// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : SA_2D
// Git hash  : cb73c1d03e6f2bcfd7eeee91a2245d4910c61e19

`timescale 1ns/1ps

module SA_2D (
  input      [7:0]    io_MatrixA_0,
  input      [7:0]    io_MatrixA_1,
  input      [7:0]    io_MatrixA_2,
  input      [7:0]    io_MatrixA_3,
  input      [7:0]    io_MatrixA_4,
  input      [7:0]    io_MatrixA_5,
  input      [7:0]    io_MatrixA_6,
  input      [7:0]    io_MatrixA_7,
  input      [7:0]    io_MatrixB_0,
  input      [7:0]    io_MatrixB_1,
  input      [7:0]    io_MatrixB_2,
  input      [7:0]    io_MatrixB_3,
  input      [7:0]    io_MatrixB_4,
  input      [7:0]    io_MatrixB_5,
  input      [7:0]    io_MatrixB_6,
  input      [7:0]    io_MatrixB_7,
  input               io_A_Valid_0,
  input               io_A_Valid_1,
  input               io_A_Valid_2,
  input               io_A_Valid_3,
  input               io_A_Valid_4,
  input               io_A_Valid_5,
  input               io_A_Valid_6,
  input               io_A_Valid_7,
  input               io_B_Valid_0,
  input               io_B_Valid_1,
  input               io_B_Valid_2,
  input               io_B_Valid_3,
  input               io_B_Valid_4,
  input               io_B_Valid_5,
  input               io_B_Valid_6,
  input               io_B_Valid_7,
  input      [15:0]   io_signCount,
  input               start,
  input               clk,
  input               reset
);

  wire                pE_64_valid;
  wire                pE_65_valid;
  wire                pE_66_valid;
  wire                pE_67_valid;
  wire                pE_68_valid;
  wire                pE_69_valid;
  wire                pE_70_valid;
  wire                pE_71_valid;
  wire                pE_72_valid;
  wire                pE_73_valid;
  wire                pE_74_valid;
  wire                pE_75_valid;
  wire                pE_76_valid;
  wire                pE_77_valid;
  wire                pE_78_valid;
  wire                pE_79_valid;
  wire                pE_80_valid;
  wire                pE_81_valid;
  wire                pE_82_valid;
  wire                pE_83_valid;
  wire                pE_84_valid;
  wire                pE_85_valid;
  wire                pE_86_valid;
  wire                pE_87_valid;
  wire                pE_88_valid;
  wire                pE_89_valid;
  wire                pE_90_valid;
  wire                pE_91_valid;
  wire                pE_92_valid;
  wire                pE_93_valid;
  wire                pE_94_valid;
  wire                pE_95_valid;
  wire                pE_96_valid;
  wire                pE_97_valid;
  wire                pE_98_valid;
  wire                pE_99_valid;
  wire                pE_100_valid;
  wire                pE_101_valid;
  wire                pE_102_valid;
  wire                pE_103_valid;
  wire                pE_104_valid;
  wire                pE_105_valid;
  wire                pE_106_valid;
  wire                pE_107_valid;
  wire                pE_108_valid;
  wire                pE_109_valid;
  wire                pE_110_valid;
  wire                pE_111_valid;
  wire                pE_112_valid;
  wire                pE_113_valid;
  wire                pE_114_valid;
  wire                pE_115_valid;
  wire                pE_116_valid;
  wire                pE_117_valid;
  wire                pE_118_valid;
  wire                pE_119_valid;
  wire                pE_120_valid;
  wire                pE_121_valid;
  wire                pE_122_valid;
  wire                pE_123_valid;
  wire                pE_124_valid;
  wire                pE_125_valid;
  wire                pE_126_valid;
  wire                pE_127_valid;
  wire       [7:0]    pE_64_acount;
  wire       [7:0]    pE_64_bcount;
  wire       [31:0]   pE_64_PE_OUT;
  wire                pE_64_finish;
  wire       [7:0]    pE_65_acount;
  wire       [7:0]    pE_65_bcount;
  wire       [31:0]   pE_65_PE_OUT;
  wire                pE_65_finish;
  wire       [7:0]    pE_66_acount;
  wire       [7:0]    pE_66_bcount;
  wire       [31:0]   pE_66_PE_OUT;
  wire                pE_66_finish;
  wire       [7:0]    pE_67_acount;
  wire       [7:0]    pE_67_bcount;
  wire       [31:0]   pE_67_PE_OUT;
  wire                pE_67_finish;
  wire       [7:0]    pE_68_acount;
  wire       [7:0]    pE_68_bcount;
  wire       [31:0]   pE_68_PE_OUT;
  wire                pE_68_finish;
  wire       [7:0]    pE_69_acount;
  wire       [7:0]    pE_69_bcount;
  wire       [31:0]   pE_69_PE_OUT;
  wire                pE_69_finish;
  wire       [7:0]    pE_70_acount;
  wire       [7:0]    pE_70_bcount;
  wire       [31:0]   pE_70_PE_OUT;
  wire                pE_70_finish;
  wire       [7:0]    pE_71_acount;
  wire       [7:0]    pE_71_bcount;
  wire       [31:0]   pE_71_PE_OUT;
  wire                pE_71_finish;
  wire       [7:0]    pE_72_acount;
  wire       [7:0]    pE_72_bcount;
  wire       [31:0]   pE_72_PE_OUT;
  wire                pE_72_finish;
  wire       [7:0]    pE_73_acount;
  wire       [7:0]    pE_73_bcount;
  wire       [31:0]   pE_73_PE_OUT;
  wire                pE_73_finish;
  wire       [7:0]    pE_74_acount;
  wire       [7:0]    pE_74_bcount;
  wire       [31:0]   pE_74_PE_OUT;
  wire                pE_74_finish;
  wire       [7:0]    pE_75_acount;
  wire       [7:0]    pE_75_bcount;
  wire       [31:0]   pE_75_PE_OUT;
  wire                pE_75_finish;
  wire       [7:0]    pE_76_acount;
  wire       [7:0]    pE_76_bcount;
  wire       [31:0]   pE_76_PE_OUT;
  wire                pE_76_finish;
  wire       [7:0]    pE_77_acount;
  wire       [7:0]    pE_77_bcount;
  wire       [31:0]   pE_77_PE_OUT;
  wire                pE_77_finish;
  wire       [7:0]    pE_78_acount;
  wire       [7:0]    pE_78_bcount;
  wire       [31:0]   pE_78_PE_OUT;
  wire                pE_78_finish;
  wire       [7:0]    pE_79_acount;
  wire       [7:0]    pE_79_bcount;
  wire       [31:0]   pE_79_PE_OUT;
  wire                pE_79_finish;
  wire       [7:0]    pE_80_acount;
  wire       [7:0]    pE_80_bcount;
  wire       [31:0]   pE_80_PE_OUT;
  wire                pE_80_finish;
  wire       [7:0]    pE_81_acount;
  wire       [7:0]    pE_81_bcount;
  wire       [31:0]   pE_81_PE_OUT;
  wire                pE_81_finish;
  wire       [7:0]    pE_82_acount;
  wire       [7:0]    pE_82_bcount;
  wire       [31:0]   pE_82_PE_OUT;
  wire                pE_82_finish;
  wire       [7:0]    pE_83_acount;
  wire       [7:0]    pE_83_bcount;
  wire       [31:0]   pE_83_PE_OUT;
  wire                pE_83_finish;
  wire       [7:0]    pE_84_acount;
  wire       [7:0]    pE_84_bcount;
  wire       [31:0]   pE_84_PE_OUT;
  wire                pE_84_finish;
  wire       [7:0]    pE_85_acount;
  wire       [7:0]    pE_85_bcount;
  wire       [31:0]   pE_85_PE_OUT;
  wire                pE_85_finish;
  wire       [7:0]    pE_86_acount;
  wire       [7:0]    pE_86_bcount;
  wire       [31:0]   pE_86_PE_OUT;
  wire                pE_86_finish;
  wire       [7:0]    pE_87_acount;
  wire       [7:0]    pE_87_bcount;
  wire       [31:0]   pE_87_PE_OUT;
  wire                pE_87_finish;
  wire       [7:0]    pE_88_acount;
  wire       [7:0]    pE_88_bcount;
  wire       [31:0]   pE_88_PE_OUT;
  wire                pE_88_finish;
  wire       [7:0]    pE_89_acount;
  wire       [7:0]    pE_89_bcount;
  wire       [31:0]   pE_89_PE_OUT;
  wire                pE_89_finish;
  wire       [7:0]    pE_90_acount;
  wire       [7:0]    pE_90_bcount;
  wire       [31:0]   pE_90_PE_OUT;
  wire                pE_90_finish;
  wire       [7:0]    pE_91_acount;
  wire       [7:0]    pE_91_bcount;
  wire       [31:0]   pE_91_PE_OUT;
  wire                pE_91_finish;
  wire       [7:0]    pE_92_acount;
  wire       [7:0]    pE_92_bcount;
  wire       [31:0]   pE_92_PE_OUT;
  wire                pE_92_finish;
  wire       [7:0]    pE_93_acount;
  wire       [7:0]    pE_93_bcount;
  wire       [31:0]   pE_93_PE_OUT;
  wire                pE_93_finish;
  wire       [7:0]    pE_94_acount;
  wire       [7:0]    pE_94_bcount;
  wire       [31:0]   pE_94_PE_OUT;
  wire                pE_94_finish;
  wire       [7:0]    pE_95_acount;
  wire       [7:0]    pE_95_bcount;
  wire       [31:0]   pE_95_PE_OUT;
  wire                pE_95_finish;
  wire       [7:0]    pE_96_acount;
  wire       [7:0]    pE_96_bcount;
  wire       [31:0]   pE_96_PE_OUT;
  wire                pE_96_finish;
  wire       [7:0]    pE_97_acount;
  wire       [7:0]    pE_97_bcount;
  wire       [31:0]   pE_97_PE_OUT;
  wire                pE_97_finish;
  wire       [7:0]    pE_98_acount;
  wire       [7:0]    pE_98_bcount;
  wire       [31:0]   pE_98_PE_OUT;
  wire                pE_98_finish;
  wire       [7:0]    pE_99_acount;
  wire       [7:0]    pE_99_bcount;
  wire       [31:0]   pE_99_PE_OUT;
  wire                pE_99_finish;
  wire       [7:0]    pE_100_acount;
  wire       [7:0]    pE_100_bcount;
  wire       [31:0]   pE_100_PE_OUT;
  wire                pE_100_finish;
  wire       [7:0]    pE_101_acount;
  wire       [7:0]    pE_101_bcount;
  wire       [31:0]   pE_101_PE_OUT;
  wire                pE_101_finish;
  wire       [7:0]    pE_102_acount;
  wire       [7:0]    pE_102_bcount;
  wire       [31:0]   pE_102_PE_OUT;
  wire                pE_102_finish;
  wire       [7:0]    pE_103_acount;
  wire       [7:0]    pE_103_bcount;
  wire       [31:0]   pE_103_PE_OUT;
  wire                pE_103_finish;
  wire       [7:0]    pE_104_acount;
  wire       [7:0]    pE_104_bcount;
  wire       [31:0]   pE_104_PE_OUT;
  wire                pE_104_finish;
  wire       [7:0]    pE_105_acount;
  wire       [7:0]    pE_105_bcount;
  wire       [31:0]   pE_105_PE_OUT;
  wire                pE_105_finish;
  wire       [7:0]    pE_106_acount;
  wire       [7:0]    pE_106_bcount;
  wire       [31:0]   pE_106_PE_OUT;
  wire                pE_106_finish;
  wire       [7:0]    pE_107_acount;
  wire       [7:0]    pE_107_bcount;
  wire       [31:0]   pE_107_PE_OUT;
  wire                pE_107_finish;
  wire       [7:0]    pE_108_acount;
  wire       [7:0]    pE_108_bcount;
  wire       [31:0]   pE_108_PE_OUT;
  wire                pE_108_finish;
  wire       [7:0]    pE_109_acount;
  wire       [7:0]    pE_109_bcount;
  wire       [31:0]   pE_109_PE_OUT;
  wire                pE_109_finish;
  wire       [7:0]    pE_110_acount;
  wire       [7:0]    pE_110_bcount;
  wire       [31:0]   pE_110_PE_OUT;
  wire                pE_110_finish;
  wire       [7:0]    pE_111_acount;
  wire       [7:0]    pE_111_bcount;
  wire       [31:0]   pE_111_PE_OUT;
  wire                pE_111_finish;
  wire       [7:0]    pE_112_acount;
  wire       [7:0]    pE_112_bcount;
  wire       [31:0]   pE_112_PE_OUT;
  wire                pE_112_finish;
  wire       [7:0]    pE_113_acount;
  wire       [7:0]    pE_113_bcount;
  wire       [31:0]   pE_113_PE_OUT;
  wire                pE_113_finish;
  wire       [7:0]    pE_114_acount;
  wire       [7:0]    pE_114_bcount;
  wire       [31:0]   pE_114_PE_OUT;
  wire                pE_114_finish;
  wire       [7:0]    pE_115_acount;
  wire       [7:0]    pE_115_bcount;
  wire       [31:0]   pE_115_PE_OUT;
  wire                pE_115_finish;
  wire       [7:0]    pE_116_acount;
  wire       [7:0]    pE_116_bcount;
  wire       [31:0]   pE_116_PE_OUT;
  wire                pE_116_finish;
  wire       [7:0]    pE_117_acount;
  wire       [7:0]    pE_117_bcount;
  wire       [31:0]   pE_117_PE_OUT;
  wire                pE_117_finish;
  wire       [7:0]    pE_118_acount;
  wire       [7:0]    pE_118_bcount;
  wire       [31:0]   pE_118_PE_OUT;
  wire                pE_118_finish;
  wire       [7:0]    pE_119_acount;
  wire       [7:0]    pE_119_bcount;
  wire       [31:0]   pE_119_PE_OUT;
  wire                pE_119_finish;
  wire       [7:0]    pE_120_acount;
  wire       [7:0]    pE_120_bcount;
  wire       [31:0]   pE_120_PE_OUT;
  wire                pE_120_finish;
  wire       [7:0]    pE_121_acount;
  wire       [7:0]    pE_121_bcount;
  wire       [31:0]   pE_121_PE_OUT;
  wire                pE_121_finish;
  wire       [7:0]    pE_122_acount;
  wire       [7:0]    pE_122_bcount;
  wire       [31:0]   pE_122_PE_OUT;
  wire                pE_122_finish;
  wire       [7:0]    pE_123_acount;
  wire       [7:0]    pE_123_bcount;
  wire       [31:0]   pE_123_PE_OUT;
  wire                pE_123_finish;
  wire       [7:0]    pE_124_acount;
  wire       [7:0]    pE_124_bcount;
  wire       [31:0]   pE_124_PE_OUT;
  wire                pE_124_finish;
  wire       [7:0]    pE_125_acount;
  wire       [7:0]    pE_125_bcount;
  wire       [31:0]   pE_125_PE_OUT;
  wire                pE_125_finish;
  wire       [7:0]    pE_126_acount;
  wire       [7:0]    pE_126_bcount;
  wire       [31:0]   pE_126_PE_OUT;
  wire                pE_126_finish;
  wire       [7:0]    pE_127_acount;
  wire       [7:0]    pE_127_bcount;
  wire       [31:0]   pE_127_PE_OUT;
  wire                pE_127_finish;
  reg        [15:0]   io_signCount_regNextWhen;
  reg                 io_A_Valid_0_delay_1;
  reg                 io_A_Valid_0_delay_1_1;
  reg                 io_A_Valid_0_delay_2;
  reg                 io_A_Valid_0_delay_1_2;
  reg                 io_A_Valid_0_delay_2_1;
  reg                 io_A_Valid_0_delay_3;
  reg                 io_A_Valid_0_delay_1_3;
  reg                 io_A_Valid_0_delay_2_2;
  reg                 io_A_Valid_0_delay_3_1;
  reg                 io_A_Valid_0_delay_4;
  reg                 io_A_Valid_0_delay_1_4;
  reg                 io_A_Valid_0_delay_2_3;
  reg                 io_A_Valid_0_delay_3_2;
  reg                 io_A_Valid_0_delay_4_1;
  reg                 io_A_Valid_0_delay_5;
  reg                 io_A_Valid_0_delay_1_5;
  reg                 io_A_Valid_0_delay_2_4;
  reg                 io_A_Valid_0_delay_3_3;
  reg                 io_A_Valid_0_delay_4_2;
  reg                 io_A_Valid_0_delay_5_1;
  reg                 io_A_Valid_0_delay_6;
  reg                 io_A_Valid_0_delay_1_6;
  reg                 io_A_Valid_0_delay_2_5;
  reg                 io_A_Valid_0_delay_3_4;
  reg                 io_A_Valid_0_delay_4_3;
  reg                 io_A_Valid_0_delay_5_2;
  reg                 io_A_Valid_0_delay_6_1;
  reg                 io_A_Valid_0_delay_7;
  reg        [15:0]   io_signCount_regNextWhen_1;
  reg                 io_B_Valid_0_delay_1;
  reg                 io_A_Valid_1_delay_1;
  reg                 io_B_Valid_1_delay_1;
  reg                 io_A_Valid_1_delay_1_1;
  reg                 io_A_Valid_1_delay_2;
  reg                 io_B_Valid_2_delay_1;
  reg                 io_A_Valid_1_delay_1_2;
  reg                 io_A_Valid_1_delay_2_1;
  reg                 io_A_Valid_1_delay_3;
  reg                 io_B_Valid_3_delay_1;
  reg                 io_A_Valid_1_delay_1_3;
  reg                 io_A_Valid_1_delay_2_2;
  reg                 io_A_Valid_1_delay_3_1;
  reg                 io_A_Valid_1_delay_4;
  reg                 io_B_Valid_4_delay_1;
  reg                 io_A_Valid_1_delay_1_4;
  reg                 io_A_Valid_1_delay_2_3;
  reg                 io_A_Valid_1_delay_3_2;
  reg                 io_A_Valid_1_delay_4_1;
  reg                 io_A_Valid_1_delay_5;
  reg                 io_B_Valid_5_delay_1;
  reg                 io_A_Valid_1_delay_1_5;
  reg                 io_A_Valid_1_delay_2_4;
  reg                 io_A_Valid_1_delay_3_3;
  reg                 io_A_Valid_1_delay_4_2;
  reg                 io_A_Valid_1_delay_5_1;
  reg                 io_A_Valid_1_delay_6;
  reg                 io_B_Valid_6_delay_1;
  reg                 io_A_Valid_1_delay_1_6;
  reg                 io_A_Valid_1_delay_2_5;
  reg                 io_A_Valid_1_delay_3_4;
  reg                 io_A_Valid_1_delay_4_3;
  reg                 io_A_Valid_1_delay_5_2;
  reg                 io_A_Valid_1_delay_6_1;
  reg                 io_A_Valid_1_delay_7;
  reg                 io_B_Valid_7_delay_1;
  reg        [15:0]   io_signCount_regNextWhen_2;
  reg                 io_B_Valid_0_delay_1_1;
  reg                 io_B_Valid_0_delay_2;
  reg                 io_A_Valid_2_delay_1;
  reg                 io_B_Valid_1_delay_1_1;
  reg                 io_B_Valid_1_delay_2;
  reg                 io_A_Valid_2_delay_1_1;
  reg                 io_A_Valid_2_delay_2;
  reg                 io_B_Valid_2_delay_1_1;
  reg                 io_B_Valid_2_delay_2;
  reg                 io_A_Valid_2_delay_1_2;
  reg                 io_A_Valid_2_delay_2_1;
  reg                 io_A_Valid_2_delay_3;
  reg                 io_B_Valid_3_delay_1_1;
  reg                 io_B_Valid_3_delay_2;
  reg                 io_A_Valid_2_delay_1_3;
  reg                 io_A_Valid_2_delay_2_2;
  reg                 io_A_Valid_2_delay_3_1;
  reg                 io_A_Valid_2_delay_4;
  reg                 io_B_Valid_4_delay_1_1;
  reg                 io_B_Valid_4_delay_2;
  reg                 io_A_Valid_2_delay_1_4;
  reg                 io_A_Valid_2_delay_2_3;
  reg                 io_A_Valid_2_delay_3_2;
  reg                 io_A_Valid_2_delay_4_1;
  reg                 io_A_Valid_2_delay_5;
  reg                 io_B_Valid_5_delay_1_1;
  reg                 io_B_Valid_5_delay_2;
  reg                 io_A_Valid_2_delay_1_5;
  reg                 io_A_Valid_2_delay_2_4;
  reg                 io_A_Valid_2_delay_3_3;
  reg                 io_A_Valid_2_delay_4_2;
  reg                 io_A_Valid_2_delay_5_1;
  reg                 io_A_Valid_2_delay_6;
  reg                 io_B_Valid_6_delay_1_1;
  reg                 io_B_Valid_6_delay_2;
  reg                 io_A_Valid_2_delay_1_6;
  reg                 io_A_Valid_2_delay_2_5;
  reg                 io_A_Valid_2_delay_3_4;
  reg                 io_A_Valid_2_delay_4_3;
  reg                 io_A_Valid_2_delay_5_2;
  reg                 io_A_Valid_2_delay_6_1;
  reg                 io_A_Valid_2_delay_7;
  reg                 io_B_Valid_7_delay_1_1;
  reg                 io_B_Valid_7_delay_2;
  reg        [15:0]   io_signCount_regNextWhen_3;
  reg                 io_B_Valid_0_delay_1_2;
  reg                 io_B_Valid_0_delay_2_1;
  reg                 io_B_Valid_0_delay_3;
  reg                 io_A_Valid_3_delay_1;
  reg                 io_B_Valid_1_delay_1_2;
  reg                 io_B_Valid_1_delay_2_1;
  reg                 io_B_Valid_1_delay_3;
  reg                 io_A_Valid_3_delay_1_1;
  reg                 io_A_Valid_3_delay_2;
  reg                 io_B_Valid_2_delay_1_2;
  reg                 io_B_Valid_2_delay_2_1;
  reg                 io_B_Valid_2_delay_3;
  reg                 io_A_Valid_3_delay_1_2;
  reg                 io_A_Valid_3_delay_2_1;
  reg                 io_A_Valid_3_delay_3;
  reg                 io_B_Valid_3_delay_1_2;
  reg                 io_B_Valid_3_delay_2_1;
  reg                 io_B_Valid_3_delay_3;
  reg                 io_A_Valid_3_delay_1_3;
  reg                 io_A_Valid_3_delay_2_2;
  reg                 io_A_Valid_3_delay_3_1;
  reg                 io_A_Valid_3_delay_4;
  reg                 io_B_Valid_4_delay_1_2;
  reg                 io_B_Valid_4_delay_2_1;
  reg                 io_B_Valid_4_delay_3;
  reg                 io_A_Valid_3_delay_1_4;
  reg                 io_A_Valid_3_delay_2_3;
  reg                 io_A_Valid_3_delay_3_2;
  reg                 io_A_Valid_3_delay_4_1;
  reg                 io_A_Valid_3_delay_5;
  reg                 io_B_Valid_5_delay_1_2;
  reg                 io_B_Valid_5_delay_2_1;
  reg                 io_B_Valid_5_delay_3;
  reg                 io_A_Valid_3_delay_1_5;
  reg                 io_A_Valid_3_delay_2_4;
  reg                 io_A_Valid_3_delay_3_3;
  reg                 io_A_Valid_3_delay_4_2;
  reg                 io_A_Valid_3_delay_5_1;
  reg                 io_A_Valid_3_delay_6;
  reg                 io_B_Valid_6_delay_1_2;
  reg                 io_B_Valid_6_delay_2_1;
  reg                 io_B_Valid_6_delay_3;
  reg                 io_A_Valid_3_delay_1_6;
  reg                 io_A_Valid_3_delay_2_5;
  reg                 io_A_Valid_3_delay_3_4;
  reg                 io_A_Valid_3_delay_4_3;
  reg                 io_A_Valid_3_delay_5_2;
  reg                 io_A_Valid_3_delay_6_1;
  reg                 io_A_Valid_3_delay_7;
  reg                 io_B_Valid_7_delay_1_2;
  reg                 io_B_Valid_7_delay_2_1;
  reg                 io_B_Valid_7_delay_3;
  reg        [15:0]   io_signCount_regNextWhen_4;
  reg                 io_B_Valid_0_delay_1_3;
  reg                 io_B_Valid_0_delay_2_2;
  reg                 io_B_Valid_0_delay_3_1;
  reg                 io_B_Valid_0_delay_4;
  reg                 io_A_Valid_4_delay_1;
  reg                 io_B_Valid_1_delay_1_3;
  reg                 io_B_Valid_1_delay_2_2;
  reg                 io_B_Valid_1_delay_3_1;
  reg                 io_B_Valid_1_delay_4;
  reg                 io_A_Valid_4_delay_1_1;
  reg                 io_A_Valid_4_delay_2;
  reg                 io_B_Valid_2_delay_1_3;
  reg                 io_B_Valid_2_delay_2_2;
  reg                 io_B_Valid_2_delay_3_1;
  reg                 io_B_Valid_2_delay_4;
  reg                 io_A_Valid_4_delay_1_2;
  reg                 io_A_Valid_4_delay_2_1;
  reg                 io_A_Valid_4_delay_3;
  reg                 io_B_Valid_3_delay_1_3;
  reg                 io_B_Valid_3_delay_2_2;
  reg                 io_B_Valid_3_delay_3_1;
  reg                 io_B_Valid_3_delay_4;
  reg                 io_A_Valid_4_delay_1_3;
  reg                 io_A_Valid_4_delay_2_2;
  reg                 io_A_Valid_4_delay_3_1;
  reg                 io_A_Valid_4_delay_4;
  reg                 io_B_Valid_4_delay_1_3;
  reg                 io_B_Valid_4_delay_2_2;
  reg                 io_B_Valid_4_delay_3_1;
  reg                 io_B_Valid_4_delay_4;
  reg                 io_A_Valid_4_delay_1_4;
  reg                 io_A_Valid_4_delay_2_3;
  reg                 io_A_Valid_4_delay_3_2;
  reg                 io_A_Valid_4_delay_4_1;
  reg                 io_A_Valid_4_delay_5;
  reg                 io_B_Valid_5_delay_1_3;
  reg                 io_B_Valid_5_delay_2_2;
  reg                 io_B_Valid_5_delay_3_1;
  reg                 io_B_Valid_5_delay_4;
  reg                 io_A_Valid_4_delay_1_5;
  reg                 io_A_Valid_4_delay_2_4;
  reg                 io_A_Valid_4_delay_3_3;
  reg                 io_A_Valid_4_delay_4_2;
  reg                 io_A_Valid_4_delay_5_1;
  reg                 io_A_Valid_4_delay_6;
  reg                 io_B_Valid_6_delay_1_3;
  reg                 io_B_Valid_6_delay_2_2;
  reg                 io_B_Valid_6_delay_3_1;
  reg                 io_B_Valid_6_delay_4;
  reg                 io_A_Valid_4_delay_1_6;
  reg                 io_A_Valid_4_delay_2_5;
  reg                 io_A_Valid_4_delay_3_4;
  reg                 io_A_Valid_4_delay_4_3;
  reg                 io_A_Valid_4_delay_5_2;
  reg                 io_A_Valid_4_delay_6_1;
  reg                 io_A_Valid_4_delay_7;
  reg                 io_B_Valid_7_delay_1_3;
  reg                 io_B_Valid_7_delay_2_2;
  reg                 io_B_Valid_7_delay_3_1;
  reg                 io_B_Valid_7_delay_4;
  reg        [15:0]   io_signCount_regNextWhen_5;
  reg                 io_B_Valid_0_delay_1_4;
  reg                 io_B_Valid_0_delay_2_3;
  reg                 io_B_Valid_0_delay_3_2;
  reg                 io_B_Valid_0_delay_4_1;
  reg                 io_B_Valid_0_delay_5;
  reg                 io_A_Valid_5_delay_1;
  reg                 io_B_Valid_1_delay_1_4;
  reg                 io_B_Valid_1_delay_2_3;
  reg                 io_B_Valid_1_delay_3_2;
  reg                 io_B_Valid_1_delay_4_1;
  reg                 io_B_Valid_1_delay_5;
  reg                 io_A_Valid_5_delay_1_1;
  reg                 io_A_Valid_5_delay_2;
  reg                 io_B_Valid_2_delay_1_4;
  reg                 io_B_Valid_2_delay_2_3;
  reg                 io_B_Valid_2_delay_3_2;
  reg                 io_B_Valid_2_delay_4_1;
  reg                 io_B_Valid_2_delay_5;
  reg                 io_A_Valid_5_delay_1_2;
  reg                 io_A_Valid_5_delay_2_1;
  reg                 io_A_Valid_5_delay_3;
  reg                 io_B_Valid_3_delay_1_4;
  reg                 io_B_Valid_3_delay_2_3;
  reg                 io_B_Valid_3_delay_3_2;
  reg                 io_B_Valid_3_delay_4_1;
  reg                 io_B_Valid_3_delay_5;
  reg                 io_A_Valid_5_delay_1_3;
  reg                 io_A_Valid_5_delay_2_2;
  reg                 io_A_Valid_5_delay_3_1;
  reg                 io_A_Valid_5_delay_4;
  reg                 io_B_Valid_4_delay_1_4;
  reg                 io_B_Valid_4_delay_2_3;
  reg                 io_B_Valid_4_delay_3_2;
  reg                 io_B_Valid_4_delay_4_1;
  reg                 io_B_Valid_4_delay_5;
  reg                 io_A_Valid_5_delay_1_4;
  reg                 io_A_Valid_5_delay_2_3;
  reg                 io_A_Valid_5_delay_3_2;
  reg                 io_A_Valid_5_delay_4_1;
  reg                 io_A_Valid_5_delay_5;
  reg                 io_B_Valid_5_delay_1_4;
  reg                 io_B_Valid_5_delay_2_3;
  reg                 io_B_Valid_5_delay_3_2;
  reg                 io_B_Valid_5_delay_4_1;
  reg                 io_B_Valid_5_delay_5;
  reg                 io_A_Valid_5_delay_1_5;
  reg                 io_A_Valid_5_delay_2_4;
  reg                 io_A_Valid_5_delay_3_3;
  reg                 io_A_Valid_5_delay_4_2;
  reg                 io_A_Valid_5_delay_5_1;
  reg                 io_A_Valid_5_delay_6;
  reg                 io_B_Valid_6_delay_1_4;
  reg                 io_B_Valid_6_delay_2_3;
  reg                 io_B_Valid_6_delay_3_2;
  reg                 io_B_Valid_6_delay_4_1;
  reg                 io_B_Valid_6_delay_5;
  reg                 io_A_Valid_5_delay_1_6;
  reg                 io_A_Valid_5_delay_2_5;
  reg                 io_A_Valid_5_delay_3_4;
  reg                 io_A_Valid_5_delay_4_3;
  reg                 io_A_Valid_5_delay_5_2;
  reg                 io_A_Valid_5_delay_6_1;
  reg                 io_A_Valid_5_delay_7;
  reg                 io_B_Valid_7_delay_1_4;
  reg                 io_B_Valid_7_delay_2_3;
  reg                 io_B_Valid_7_delay_3_2;
  reg                 io_B_Valid_7_delay_4_1;
  reg                 io_B_Valid_7_delay_5;
  reg        [15:0]   io_signCount_regNextWhen_6;
  reg                 io_B_Valid_0_delay_1_5;
  reg                 io_B_Valid_0_delay_2_4;
  reg                 io_B_Valid_0_delay_3_3;
  reg                 io_B_Valid_0_delay_4_2;
  reg                 io_B_Valid_0_delay_5_1;
  reg                 io_B_Valid_0_delay_6;
  reg                 io_A_Valid_6_delay_1;
  reg                 io_B_Valid_1_delay_1_5;
  reg                 io_B_Valid_1_delay_2_4;
  reg                 io_B_Valid_1_delay_3_3;
  reg                 io_B_Valid_1_delay_4_2;
  reg                 io_B_Valid_1_delay_5_1;
  reg                 io_B_Valid_1_delay_6;
  reg                 io_A_Valid_6_delay_1_1;
  reg                 io_A_Valid_6_delay_2;
  reg                 io_B_Valid_2_delay_1_5;
  reg                 io_B_Valid_2_delay_2_4;
  reg                 io_B_Valid_2_delay_3_3;
  reg                 io_B_Valid_2_delay_4_2;
  reg                 io_B_Valid_2_delay_5_1;
  reg                 io_B_Valid_2_delay_6;
  reg                 io_A_Valid_6_delay_1_2;
  reg                 io_A_Valid_6_delay_2_1;
  reg                 io_A_Valid_6_delay_3;
  reg                 io_B_Valid_3_delay_1_5;
  reg                 io_B_Valid_3_delay_2_4;
  reg                 io_B_Valid_3_delay_3_3;
  reg                 io_B_Valid_3_delay_4_2;
  reg                 io_B_Valid_3_delay_5_1;
  reg                 io_B_Valid_3_delay_6;
  reg                 io_A_Valid_6_delay_1_3;
  reg                 io_A_Valid_6_delay_2_2;
  reg                 io_A_Valid_6_delay_3_1;
  reg                 io_A_Valid_6_delay_4;
  reg                 io_B_Valid_4_delay_1_5;
  reg                 io_B_Valid_4_delay_2_4;
  reg                 io_B_Valid_4_delay_3_3;
  reg                 io_B_Valid_4_delay_4_2;
  reg                 io_B_Valid_4_delay_5_1;
  reg                 io_B_Valid_4_delay_6;
  reg                 io_A_Valid_6_delay_1_4;
  reg                 io_A_Valid_6_delay_2_3;
  reg                 io_A_Valid_6_delay_3_2;
  reg                 io_A_Valid_6_delay_4_1;
  reg                 io_A_Valid_6_delay_5;
  reg                 io_B_Valid_5_delay_1_5;
  reg                 io_B_Valid_5_delay_2_4;
  reg                 io_B_Valid_5_delay_3_3;
  reg                 io_B_Valid_5_delay_4_2;
  reg                 io_B_Valid_5_delay_5_1;
  reg                 io_B_Valid_5_delay_6;
  reg                 io_A_Valid_6_delay_1_5;
  reg                 io_A_Valid_6_delay_2_4;
  reg                 io_A_Valid_6_delay_3_3;
  reg                 io_A_Valid_6_delay_4_2;
  reg                 io_A_Valid_6_delay_5_1;
  reg                 io_A_Valid_6_delay_6;
  reg                 io_B_Valid_6_delay_1_5;
  reg                 io_B_Valid_6_delay_2_4;
  reg                 io_B_Valid_6_delay_3_3;
  reg                 io_B_Valid_6_delay_4_2;
  reg                 io_B_Valid_6_delay_5_1;
  reg                 io_B_Valid_6_delay_6;
  reg                 io_A_Valid_6_delay_1_6;
  reg                 io_A_Valid_6_delay_2_5;
  reg                 io_A_Valid_6_delay_3_4;
  reg                 io_A_Valid_6_delay_4_3;
  reg                 io_A_Valid_6_delay_5_2;
  reg                 io_A_Valid_6_delay_6_1;
  reg                 io_A_Valid_6_delay_7;
  reg                 io_B_Valid_7_delay_1_5;
  reg                 io_B_Valid_7_delay_2_4;
  reg                 io_B_Valid_7_delay_3_3;
  reg                 io_B_Valid_7_delay_4_2;
  reg                 io_B_Valid_7_delay_5_1;
  reg                 io_B_Valid_7_delay_6;
  reg        [15:0]   io_signCount_regNextWhen_7;
  reg                 io_B_Valid_0_delay_1_6;
  reg                 io_B_Valid_0_delay_2_5;
  reg                 io_B_Valid_0_delay_3_4;
  reg                 io_B_Valid_0_delay_4_3;
  reg                 io_B_Valid_0_delay_5_2;
  reg                 io_B_Valid_0_delay_6_1;
  reg                 io_B_Valid_0_delay_7;
  reg                 io_A_Valid_7_delay_1;
  reg                 io_B_Valid_1_delay_1_6;
  reg                 io_B_Valid_1_delay_2_5;
  reg                 io_B_Valid_1_delay_3_4;
  reg                 io_B_Valid_1_delay_4_3;
  reg                 io_B_Valid_1_delay_5_2;
  reg                 io_B_Valid_1_delay_6_1;
  reg                 io_B_Valid_1_delay_7;
  reg                 io_A_Valid_7_delay_1_1;
  reg                 io_A_Valid_7_delay_2;
  reg                 io_B_Valid_2_delay_1_6;
  reg                 io_B_Valid_2_delay_2_5;
  reg                 io_B_Valid_2_delay_3_4;
  reg                 io_B_Valid_2_delay_4_3;
  reg                 io_B_Valid_2_delay_5_2;
  reg                 io_B_Valid_2_delay_6_1;
  reg                 io_B_Valid_2_delay_7;
  reg                 io_A_Valid_7_delay_1_2;
  reg                 io_A_Valid_7_delay_2_1;
  reg                 io_A_Valid_7_delay_3;
  reg                 io_B_Valid_3_delay_1_6;
  reg                 io_B_Valid_3_delay_2_5;
  reg                 io_B_Valid_3_delay_3_4;
  reg                 io_B_Valid_3_delay_4_3;
  reg                 io_B_Valid_3_delay_5_2;
  reg                 io_B_Valid_3_delay_6_1;
  reg                 io_B_Valid_3_delay_7;
  reg                 io_A_Valid_7_delay_1_3;
  reg                 io_A_Valid_7_delay_2_2;
  reg                 io_A_Valid_7_delay_3_1;
  reg                 io_A_Valid_7_delay_4;
  reg                 io_B_Valid_4_delay_1_6;
  reg                 io_B_Valid_4_delay_2_5;
  reg                 io_B_Valid_4_delay_3_4;
  reg                 io_B_Valid_4_delay_4_3;
  reg                 io_B_Valid_4_delay_5_2;
  reg                 io_B_Valid_4_delay_6_1;
  reg                 io_B_Valid_4_delay_7;
  reg                 io_A_Valid_7_delay_1_4;
  reg                 io_A_Valid_7_delay_2_3;
  reg                 io_A_Valid_7_delay_3_2;
  reg                 io_A_Valid_7_delay_4_1;
  reg                 io_A_Valid_7_delay_5;
  reg                 io_B_Valid_5_delay_1_6;
  reg                 io_B_Valid_5_delay_2_5;
  reg                 io_B_Valid_5_delay_3_4;
  reg                 io_B_Valid_5_delay_4_3;
  reg                 io_B_Valid_5_delay_5_2;
  reg                 io_B_Valid_5_delay_6_1;
  reg                 io_B_Valid_5_delay_7;
  reg                 io_A_Valid_7_delay_1_5;
  reg                 io_A_Valid_7_delay_2_4;
  reg                 io_A_Valid_7_delay_3_3;
  reg                 io_A_Valid_7_delay_4_2;
  reg                 io_A_Valid_7_delay_5_1;
  reg                 io_A_Valid_7_delay_6;
  reg                 io_B_Valid_6_delay_1_6;
  reg                 io_B_Valid_6_delay_2_5;
  reg                 io_B_Valid_6_delay_3_4;
  reg                 io_B_Valid_6_delay_4_3;
  reg                 io_B_Valid_6_delay_5_2;
  reg                 io_B_Valid_6_delay_6_1;
  reg                 io_B_Valid_6_delay_7;
  reg                 io_A_Valid_7_delay_1_6;
  reg                 io_A_Valid_7_delay_2_5;
  reg                 io_A_Valid_7_delay_3_4;
  reg                 io_A_Valid_7_delay_4_3;
  reg                 io_A_Valid_7_delay_5_2;
  reg                 io_A_Valid_7_delay_6_1;
  reg                 io_A_Valid_7_delay_7;
  reg                 io_B_Valid_7_delay_1_6;
  reg                 io_B_Valid_7_delay_2_5;
  reg                 io_B_Valid_7_delay_3_4;
  reg                 io_B_Valid_7_delay_4_3;
  reg                 io_B_Valid_7_delay_5_2;
  reg                 io_B_Valid_7_delay_6_1;
  reg                 io_B_Valid_7_delay_7;

  PE pE_64 (
    .activate  (io_MatrixA_0[7:0]             ), //i
    .weight    (io_MatrixB_0[7:0]             ), //i
    .valid     (pE_64_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_64_acount[7:0]             ), //o
    .bcount    (pE_64_bcount[7:0]             ), //o
    .PE_OUT    (pE_64_PE_OUT[31:0]            ), //o
    .finish    (pE_64_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE pE_65 (
    .activate  (pE_64_acount[7:0]             ), //i
    .weight    (io_MatrixB_1[7:0]             ), //i
    .valid     (pE_65_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_65_acount[7:0]             ), //o
    .bcount    (pE_65_bcount[7:0]             ), //o
    .PE_OUT    (pE_65_PE_OUT[31:0]            ), //o
    .finish    (pE_65_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE pE_66 (
    .activate  (pE_65_acount[7:0]             ), //i
    .weight    (io_MatrixB_2[7:0]             ), //i
    .valid     (pE_66_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_66_acount[7:0]             ), //o
    .bcount    (pE_66_bcount[7:0]             ), //o
    .PE_OUT    (pE_66_PE_OUT[31:0]            ), //o
    .finish    (pE_66_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE pE_67 (
    .activate  (pE_66_acount[7:0]             ), //i
    .weight    (io_MatrixB_3[7:0]             ), //i
    .valid     (pE_67_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_67_acount[7:0]             ), //o
    .bcount    (pE_67_bcount[7:0]             ), //o
    .PE_OUT    (pE_67_PE_OUT[31:0]            ), //o
    .finish    (pE_67_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE pE_68 (
    .activate  (pE_67_acount[7:0]             ), //i
    .weight    (io_MatrixB_4[7:0]             ), //i
    .valid     (pE_68_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_68_acount[7:0]             ), //o
    .bcount    (pE_68_bcount[7:0]             ), //o
    .PE_OUT    (pE_68_PE_OUT[31:0]            ), //o
    .finish    (pE_68_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE pE_69 (
    .activate  (pE_68_acount[7:0]             ), //i
    .weight    (io_MatrixB_5[7:0]             ), //i
    .valid     (pE_69_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_69_acount[7:0]             ), //o
    .bcount    (pE_69_bcount[7:0]             ), //o
    .PE_OUT    (pE_69_PE_OUT[31:0]            ), //o
    .finish    (pE_69_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE pE_70 (
    .activate  (pE_69_acount[7:0]             ), //i
    .weight    (io_MatrixB_6[7:0]             ), //i
    .valid     (pE_70_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_70_acount[7:0]             ), //o
    .bcount    (pE_70_bcount[7:0]             ), //o
    .PE_OUT    (pE_70_PE_OUT[31:0]            ), //o
    .finish    (pE_70_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE pE_71 (
    .activate  (pE_70_acount[7:0]             ), //i
    .weight    (io_MatrixB_7[7:0]             ), //i
    .valid     (pE_71_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_71_acount[7:0]             ), //o
    .bcount    (pE_71_bcount[7:0]             ), //o
    .PE_OUT    (pE_71_PE_OUT[31:0]            ), //o
    .finish    (pE_71_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE pE_72 (
    .activate  (pE_72_acount[7:0]               ), //i
    .weight    (pE_64_bcount[7:0]               ), //i
    .valid     (pE_72_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_72_acount[7:0]               ), //o
    .bcount    (pE_72_bcount[7:0]               ), //o
    .PE_OUT    (pE_72_PE_OUT[31:0]              ), //o
    .finish    (pE_72_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_73 (
    .activate  (pE_64_acount[7:0]               ), //i
    .weight    (pE_64_bcount[7:0]               ), //i
    .valid     (pE_73_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_73_acount[7:0]               ), //o
    .bcount    (pE_73_bcount[7:0]               ), //o
    .PE_OUT    (pE_73_PE_OUT[31:0]              ), //o
    .finish    (pE_73_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_74 (
    .activate  (pE_65_acount[7:0]               ), //i
    .weight    (pE_65_bcount[7:0]               ), //i
    .valid     (pE_74_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_74_acount[7:0]               ), //o
    .bcount    (pE_74_bcount[7:0]               ), //o
    .PE_OUT    (pE_74_PE_OUT[31:0]              ), //o
    .finish    (pE_74_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_75 (
    .activate  (pE_66_acount[7:0]               ), //i
    .weight    (pE_66_bcount[7:0]               ), //i
    .valid     (pE_75_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_75_acount[7:0]               ), //o
    .bcount    (pE_75_bcount[7:0]               ), //o
    .PE_OUT    (pE_75_PE_OUT[31:0]              ), //o
    .finish    (pE_75_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_76 (
    .activate  (pE_67_acount[7:0]               ), //i
    .weight    (pE_67_bcount[7:0]               ), //i
    .valid     (pE_76_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_76_acount[7:0]               ), //o
    .bcount    (pE_76_bcount[7:0]               ), //o
    .PE_OUT    (pE_76_PE_OUT[31:0]              ), //o
    .finish    (pE_76_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_77 (
    .activate  (pE_68_acount[7:0]               ), //i
    .weight    (pE_68_bcount[7:0]               ), //i
    .valid     (pE_77_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_77_acount[7:0]               ), //o
    .bcount    (pE_77_bcount[7:0]               ), //o
    .PE_OUT    (pE_77_PE_OUT[31:0]              ), //o
    .finish    (pE_77_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_78 (
    .activate  (pE_69_acount[7:0]               ), //i
    .weight    (pE_69_bcount[7:0]               ), //i
    .valid     (pE_78_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_78_acount[7:0]               ), //o
    .bcount    (pE_78_bcount[7:0]               ), //o
    .PE_OUT    (pE_78_PE_OUT[31:0]              ), //o
    .finish    (pE_78_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_79 (
    .activate  (pE_70_acount[7:0]               ), //i
    .weight    (pE_70_bcount[7:0]               ), //i
    .valid     (pE_79_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_79_acount[7:0]               ), //o
    .bcount    (pE_79_bcount[7:0]               ), //o
    .PE_OUT    (pE_79_PE_OUT[31:0]              ), //o
    .finish    (pE_79_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_80 (
    .activate  (pE_80_acount[7:0]               ), //i
    .weight    (pE_72_bcount[7:0]               ), //i
    .valid     (pE_80_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_80_acount[7:0]               ), //o
    .bcount    (pE_80_bcount[7:0]               ), //o
    .PE_OUT    (pE_80_PE_OUT[31:0]              ), //o
    .finish    (pE_80_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_81 (
    .activate  (pE_72_acount[7:0]               ), //i
    .weight    (pE_72_bcount[7:0]               ), //i
    .valid     (pE_81_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_81_acount[7:0]               ), //o
    .bcount    (pE_81_bcount[7:0]               ), //o
    .PE_OUT    (pE_81_PE_OUT[31:0]              ), //o
    .finish    (pE_81_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_82 (
    .activate  (pE_73_acount[7:0]               ), //i
    .weight    (pE_73_bcount[7:0]               ), //i
    .valid     (pE_82_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_82_acount[7:0]               ), //o
    .bcount    (pE_82_bcount[7:0]               ), //o
    .PE_OUT    (pE_82_PE_OUT[31:0]              ), //o
    .finish    (pE_82_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_83 (
    .activate  (pE_74_acount[7:0]               ), //i
    .weight    (pE_74_bcount[7:0]               ), //i
    .valid     (pE_83_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_83_acount[7:0]               ), //o
    .bcount    (pE_83_bcount[7:0]               ), //o
    .PE_OUT    (pE_83_PE_OUT[31:0]              ), //o
    .finish    (pE_83_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_84 (
    .activate  (pE_75_acount[7:0]               ), //i
    .weight    (pE_75_bcount[7:0]               ), //i
    .valid     (pE_84_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_84_acount[7:0]               ), //o
    .bcount    (pE_84_bcount[7:0]               ), //o
    .PE_OUT    (pE_84_PE_OUT[31:0]              ), //o
    .finish    (pE_84_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_85 (
    .activate  (pE_76_acount[7:0]               ), //i
    .weight    (pE_76_bcount[7:0]               ), //i
    .valid     (pE_85_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_85_acount[7:0]               ), //o
    .bcount    (pE_85_bcount[7:0]               ), //o
    .PE_OUT    (pE_85_PE_OUT[31:0]              ), //o
    .finish    (pE_85_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_86 (
    .activate  (pE_77_acount[7:0]               ), //i
    .weight    (pE_77_bcount[7:0]               ), //i
    .valid     (pE_86_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_86_acount[7:0]               ), //o
    .bcount    (pE_86_bcount[7:0]               ), //o
    .PE_OUT    (pE_86_PE_OUT[31:0]              ), //o
    .finish    (pE_86_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_87 (
    .activate  (pE_78_acount[7:0]               ), //i
    .weight    (pE_78_bcount[7:0]               ), //i
    .valid     (pE_87_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_87_acount[7:0]               ), //o
    .bcount    (pE_87_bcount[7:0]               ), //o
    .PE_OUT    (pE_87_PE_OUT[31:0]              ), //o
    .finish    (pE_87_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_88 (
    .activate  (pE_88_acount[7:0]               ), //i
    .weight    (pE_80_bcount[7:0]               ), //i
    .valid     (pE_88_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_88_acount[7:0]               ), //o
    .bcount    (pE_88_bcount[7:0]               ), //o
    .PE_OUT    (pE_88_PE_OUT[31:0]              ), //o
    .finish    (pE_88_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_89 (
    .activate  (pE_80_acount[7:0]               ), //i
    .weight    (pE_80_bcount[7:0]               ), //i
    .valid     (pE_89_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_89_acount[7:0]               ), //o
    .bcount    (pE_89_bcount[7:0]               ), //o
    .PE_OUT    (pE_89_PE_OUT[31:0]              ), //o
    .finish    (pE_89_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_90 (
    .activate  (pE_81_acount[7:0]               ), //i
    .weight    (pE_81_bcount[7:0]               ), //i
    .valid     (pE_90_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_90_acount[7:0]               ), //o
    .bcount    (pE_90_bcount[7:0]               ), //o
    .PE_OUT    (pE_90_PE_OUT[31:0]              ), //o
    .finish    (pE_90_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_91 (
    .activate  (pE_82_acount[7:0]               ), //i
    .weight    (pE_82_bcount[7:0]               ), //i
    .valid     (pE_91_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_91_acount[7:0]               ), //o
    .bcount    (pE_91_bcount[7:0]               ), //o
    .PE_OUT    (pE_91_PE_OUT[31:0]              ), //o
    .finish    (pE_91_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_92 (
    .activate  (pE_83_acount[7:0]               ), //i
    .weight    (pE_83_bcount[7:0]               ), //i
    .valid     (pE_92_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_92_acount[7:0]               ), //o
    .bcount    (pE_92_bcount[7:0]               ), //o
    .PE_OUT    (pE_92_PE_OUT[31:0]              ), //o
    .finish    (pE_92_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_93 (
    .activate  (pE_84_acount[7:0]               ), //i
    .weight    (pE_84_bcount[7:0]               ), //i
    .valid     (pE_93_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_93_acount[7:0]               ), //o
    .bcount    (pE_93_bcount[7:0]               ), //o
    .PE_OUT    (pE_93_PE_OUT[31:0]              ), //o
    .finish    (pE_93_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_94 (
    .activate  (pE_85_acount[7:0]               ), //i
    .weight    (pE_85_bcount[7:0]               ), //i
    .valid     (pE_94_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_94_acount[7:0]               ), //o
    .bcount    (pE_94_bcount[7:0]               ), //o
    .PE_OUT    (pE_94_PE_OUT[31:0]              ), //o
    .finish    (pE_94_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_95 (
    .activate  (pE_86_acount[7:0]               ), //i
    .weight    (pE_86_bcount[7:0]               ), //i
    .valid     (pE_95_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_95_acount[7:0]               ), //o
    .bcount    (pE_95_bcount[7:0]               ), //o
    .PE_OUT    (pE_95_PE_OUT[31:0]              ), //o
    .finish    (pE_95_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_96 (
    .activate  (pE_96_acount[7:0]               ), //i
    .weight    (pE_88_bcount[7:0]               ), //i
    .valid     (pE_96_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_96_acount[7:0]               ), //o
    .bcount    (pE_96_bcount[7:0]               ), //o
    .PE_OUT    (pE_96_PE_OUT[31:0]              ), //o
    .finish    (pE_96_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_97 (
    .activate  (pE_88_acount[7:0]               ), //i
    .weight    (pE_88_bcount[7:0]               ), //i
    .valid     (pE_97_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_97_acount[7:0]               ), //o
    .bcount    (pE_97_bcount[7:0]               ), //o
    .PE_OUT    (pE_97_PE_OUT[31:0]              ), //o
    .finish    (pE_97_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_98 (
    .activate  (pE_89_acount[7:0]               ), //i
    .weight    (pE_89_bcount[7:0]               ), //i
    .valid     (pE_98_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_98_acount[7:0]               ), //o
    .bcount    (pE_98_bcount[7:0]               ), //o
    .PE_OUT    (pE_98_PE_OUT[31:0]              ), //o
    .finish    (pE_98_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_99 (
    .activate  (pE_90_acount[7:0]               ), //i
    .weight    (pE_90_bcount[7:0]               ), //i
    .valid     (pE_99_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_99_acount[7:0]               ), //o
    .bcount    (pE_99_bcount[7:0]               ), //o
    .PE_OUT    (pE_99_PE_OUT[31:0]              ), //o
    .finish    (pE_99_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_100 (
    .activate  (pE_91_acount[7:0]               ), //i
    .weight    (pE_91_bcount[7:0]               ), //i
    .valid     (pE_100_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_100_acount[7:0]              ), //o
    .bcount    (pE_100_bcount[7:0]              ), //o
    .PE_OUT    (pE_100_PE_OUT[31:0]             ), //o
    .finish    (pE_100_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_101 (
    .activate  (pE_92_acount[7:0]               ), //i
    .weight    (pE_92_bcount[7:0]               ), //i
    .valid     (pE_101_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_101_acount[7:0]              ), //o
    .bcount    (pE_101_bcount[7:0]              ), //o
    .PE_OUT    (pE_101_PE_OUT[31:0]             ), //o
    .finish    (pE_101_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_102 (
    .activate  (pE_93_acount[7:0]               ), //i
    .weight    (pE_93_bcount[7:0]               ), //i
    .valid     (pE_102_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_102_acount[7:0]              ), //o
    .bcount    (pE_102_bcount[7:0]              ), //o
    .PE_OUT    (pE_102_PE_OUT[31:0]             ), //o
    .finish    (pE_102_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_103 (
    .activate  (pE_94_acount[7:0]               ), //i
    .weight    (pE_94_bcount[7:0]               ), //i
    .valid     (pE_103_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_103_acount[7:0]              ), //o
    .bcount    (pE_103_bcount[7:0]              ), //o
    .PE_OUT    (pE_103_PE_OUT[31:0]             ), //o
    .finish    (pE_103_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_104 (
    .activate  (pE_104_acount[7:0]              ), //i
    .weight    (pE_96_bcount[7:0]               ), //i
    .valid     (pE_104_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_104_acount[7:0]              ), //o
    .bcount    (pE_104_bcount[7:0]              ), //o
    .PE_OUT    (pE_104_PE_OUT[31:0]             ), //o
    .finish    (pE_104_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_105 (
    .activate  (pE_96_acount[7:0]               ), //i
    .weight    (pE_96_bcount[7:0]               ), //i
    .valid     (pE_105_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_105_acount[7:0]              ), //o
    .bcount    (pE_105_bcount[7:0]              ), //o
    .PE_OUT    (pE_105_PE_OUT[31:0]             ), //o
    .finish    (pE_105_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_106 (
    .activate  (pE_97_acount[7:0]               ), //i
    .weight    (pE_97_bcount[7:0]               ), //i
    .valid     (pE_106_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_106_acount[7:0]              ), //o
    .bcount    (pE_106_bcount[7:0]              ), //o
    .PE_OUT    (pE_106_PE_OUT[31:0]             ), //o
    .finish    (pE_106_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_107 (
    .activate  (pE_98_acount[7:0]               ), //i
    .weight    (pE_98_bcount[7:0]               ), //i
    .valid     (pE_107_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_107_acount[7:0]              ), //o
    .bcount    (pE_107_bcount[7:0]              ), //o
    .PE_OUT    (pE_107_PE_OUT[31:0]             ), //o
    .finish    (pE_107_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_108 (
    .activate  (pE_99_acount[7:0]               ), //i
    .weight    (pE_99_bcount[7:0]               ), //i
    .valid     (pE_108_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_108_acount[7:0]              ), //o
    .bcount    (pE_108_bcount[7:0]              ), //o
    .PE_OUT    (pE_108_PE_OUT[31:0]             ), //o
    .finish    (pE_108_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_109 (
    .activate  (pE_100_acount[7:0]              ), //i
    .weight    (pE_100_bcount[7:0]              ), //i
    .valid     (pE_109_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_109_acount[7:0]              ), //o
    .bcount    (pE_109_bcount[7:0]              ), //o
    .PE_OUT    (pE_109_PE_OUT[31:0]             ), //o
    .finish    (pE_109_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_110 (
    .activate  (pE_101_acount[7:0]              ), //i
    .weight    (pE_101_bcount[7:0]              ), //i
    .valid     (pE_110_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_110_acount[7:0]              ), //o
    .bcount    (pE_110_bcount[7:0]              ), //o
    .PE_OUT    (pE_110_PE_OUT[31:0]             ), //o
    .finish    (pE_110_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_111 (
    .activate  (pE_102_acount[7:0]              ), //i
    .weight    (pE_102_bcount[7:0]              ), //i
    .valid     (pE_111_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_111_acount[7:0]              ), //o
    .bcount    (pE_111_bcount[7:0]              ), //o
    .PE_OUT    (pE_111_PE_OUT[31:0]             ), //o
    .finish    (pE_111_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_112 (
    .activate  (pE_112_acount[7:0]              ), //i
    .weight    (pE_104_bcount[7:0]              ), //i
    .valid     (pE_112_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_112_acount[7:0]              ), //o
    .bcount    (pE_112_bcount[7:0]              ), //o
    .PE_OUT    (pE_112_PE_OUT[31:0]             ), //o
    .finish    (pE_112_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_113 (
    .activate  (pE_104_acount[7:0]              ), //i
    .weight    (pE_104_bcount[7:0]              ), //i
    .valid     (pE_113_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_113_acount[7:0]              ), //o
    .bcount    (pE_113_bcount[7:0]              ), //o
    .PE_OUT    (pE_113_PE_OUT[31:0]             ), //o
    .finish    (pE_113_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_114 (
    .activate  (pE_105_acount[7:0]              ), //i
    .weight    (pE_105_bcount[7:0]              ), //i
    .valid     (pE_114_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_114_acount[7:0]              ), //o
    .bcount    (pE_114_bcount[7:0]              ), //o
    .PE_OUT    (pE_114_PE_OUT[31:0]             ), //o
    .finish    (pE_114_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_115 (
    .activate  (pE_106_acount[7:0]              ), //i
    .weight    (pE_106_bcount[7:0]              ), //i
    .valid     (pE_115_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_115_acount[7:0]              ), //o
    .bcount    (pE_115_bcount[7:0]              ), //o
    .PE_OUT    (pE_115_PE_OUT[31:0]             ), //o
    .finish    (pE_115_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_116 (
    .activate  (pE_107_acount[7:0]              ), //i
    .weight    (pE_107_bcount[7:0]              ), //i
    .valid     (pE_116_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_116_acount[7:0]              ), //o
    .bcount    (pE_116_bcount[7:0]              ), //o
    .PE_OUT    (pE_116_PE_OUT[31:0]             ), //o
    .finish    (pE_116_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_117 (
    .activate  (pE_108_acount[7:0]              ), //i
    .weight    (pE_108_bcount[7:0]              ), //i
    .valid     (pE_117_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_117_acount[7:0]              ), //o
    .bcount    (pE_117_bcount[7:0]              ), //o
    .PE_OUT    (pE_117_PE_OUT[31:0]             ), //o
    .finish    (pE_117_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_118 (
    .activate  (pE_109_acount[7:0]              ), //i
    .weight    (pE_109_bcount[7:0]              ), //i
    .valid     (pE_118_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_118_acount[7:0]              ), //o
    .bcount    (pE_118_bcount[7:0]              ), //o
    .PE_OUT    (pE_118_PE_OUT[31:0]             ), //o
    .finish    (pE_118_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_119 (
    .activate  (pE_110_acount[7:0]              ), //i
    .weight    (pE_110_bcount[7:0]              ), //i
    .valid     (pE_119_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_119_acount[7:0]              ), //o
    .bcount    (pE_119_bcount[7:0]              ), //o
    .PE_OUT    (pE_119_PE_OUT[31:0]             ), //o
    .finish    (pE_119_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_120 (
    .activate  (pE_120_acount[7:0]              ), //i
    .weight    (pE_112_bcount[7:0]              ), //i
    .valid     (pE_120_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_120_acount[7:0]              ), //o
    .bcount    (pE_120_bcount[7:0]              ), //o
    .PE_OUT    (pE_120_PE_OUT[31:0]             ), //o
    .finish    (pE_120_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_121 (
    .activate  (pE_112_acount[7:0]              ), //i
    .weight    (pE_112_bcount[7:0]              ), //i
    .valid     (pE_121_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_121_acount[7:0]              ), //o
    .bcount    (pE_121_bcount[7:0]              ), //o
    .PE_OUT    (pE_121_PE_OUT[31:0]             ), //o
    .finish    (pE_121_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_122 (
    .activate  (pE_113_acount[7:0]              ), //i
    .weight    (pE_113_bcount[7:0]              ), //i
    .valid     (pE_122_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_122_acount[7:0]              ), //o
    .bcount    (pE_122_bcount[7:0]              ), //o
    .PE_OUT    (pE_122_PE_OUT[31:0]             ), //o
    .finish    (pE_122_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_123 (
    .activate  (pE_114_acount[7:0]              ), //i
    .weight    (pE_114_bcount[7:0]              ), //i
    .valid     (pE_123_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_123_acount[7:0]              ), //o
    .bcount    (pE_123_bcount[7:0]              ), //o
    .PE_OUT    (pE_123_PE_OUT[31:0]             ), //o
    .finish    (pE_123_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_124 (
    .activate  (pE_115_acount[7:0]              ), //i
    .weight    (pE_115_bcount[7:0]              ), //i
    .valid     (pE_124_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_124_acount[7:0]              ), //o
    .bcount    (pE_124_bcount[7:0]              ), //o
    .PE_OUT    (pE_124_PE_OUT[31:0]             ), //o
    .finish    (pE_124_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_125 (
    .activate  (pE_116_acount[7:0]              ), //i
    .weight    (pE_116_bcount[7:0]              ), //i
    .valid     (pE_125_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_125_acount[7:0]              ), //o
    .bcount    (pE_125_bcount[7:0]              ), //o
    .PE_OUT    (pE_125_PE_OUT[31:0]             ), //o
    .finish    (pE_125_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_126 (
    .activate  (pE_117_acount[7:0]              ), //i
    .weight    (pE_117_bcount[7:0]              ), //i
    .valid     (pE_126_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_126_acount[7:0]              ), //o
    .bcount    (pE_126_bcount[7:0]              ), //o
    .PE_OUT    (pE_126_PE_OUT[31:0]             ), //o
    .finish    (pE_126_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE pE_127 (
    .activate  (pE_118_acount[7:0]              ), //i
    .weight    (pE_118_bcount[7:0]              ), //i
    .valid     (pE_127_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_127_acount[7:0]              ), //o
    .bcount    (pE_127_bcount[7:0]              ), //o
    .PE_OUT    (pE_127_PE_OUT[31:0]             ), //o
    .finish    (pE_127_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  assign pE_64_valid = (io_A_Valid_0 && io_B_Valid_0);
  assign pE_65_valid = (io_A_Valid_0_delay_1 && io_B_Valid_1);
  assign pE_66_valid = (io_A_Valid_0_delay_2 && io_B_Valid_2);
  assign pE_67_valid = (io_A_Valid_0_delay_3 && io_B_Valid_3);
  assign pE_68_valid = (io_A_Valid_0_delay_4 && io_B_Valid_4);
  assign pE_69_valid = (io_A_Valid_0_delay_5 && io_B_Valid_5);
  assign pE_70_valid = (io_A_Valid_0_delay_6 && io_B_Valid_6);
  assign pE_71_valid = (io_A_Valid_0_delay_7 && io_B_Valid_7);
  assign pE_72_valid = (io_A_Valid_1 && io_B_Valid_0_delay_1);
  assign pE_73_valid = (io_A_Valid_1_delay_1 && io_B_Valid_1_delay_1);
  assign pE_74_valid = (io_A_Valid_1_delay_2 && io_B_Valid_2_delay_1);
  assign pE_75_valid = (io_A_Valid_1_delay_3 && io_B_Valid_3_delay_1);
  assign pE_76_valid = (io_A_Valid_1_delay_4 && io_B_Valid_4_delay_1);
  assign pE_77_valid = (io_A_Valid_1_delay_5 && io_B_Valid_5_delay_1);
  assign pE_78_valid = (io_A_Valid_1_delay_6 && io_B_Valid_6_delay_1);
  assign pE_79_valid = (io_A_Valid_1_delay_7 && io_B_Valid_7_delay_1);
  assign pE_80_valid = (io_A_Valid_2 && io_B_Valid_0_delay_2);
  assign pE_81_valid = (io_A_Valid_2_delay_1 && io_B_Valid_1_delay_2);
  assign pE_82_valid = (io_A_Valid_2_delay_2 && io_B_Valid_2_delay_2);
  assign pE_83_valid = (io_A_Valid_2_delay_3 && io_B_Valid_3_delay_2);
  assign pE_84_valid = (io_A_Valid_2_delay_4 && io_B_Valid_4_delay_2);
  assign pE_85_valid = (io_A_Valid_2_delay_5 && io_B_Valid_5_delay_2);
  assign pE_86_valid = (io_A_Valid_2_delay_6 && io_B_Valid_6_delay_2);
  assign pE_87_valid = (io_A_Valid_2_delay_7 && io_B_Valid_7_delay_2);
  assign pE_88_valid = (io_A_Valid_3 && io_B_Valid_0_delay_3);
  assign pE_89_valid = (io_A_Valid_3_delay_1 && io_B_Valid_1_delay_3);
  assign pE_90_valid = (io_A_Valid_3_delay_2 && io_B_Valid_2_delay_3);
  assign pE_91_valid = (io_A_Valid_3_delay_3 && io_B_Valid_3_delay_3);
  assign pE_92_valid = (io_A_Valid_3_delay_4 && io_B_Valid_4_delay_3);
  assign pE_93_valid = (io_A_Valid_3_delay_5 && io_B_Valid_5_delay_3);
  assign pE_94_valid = (io_A_Valid_3_delay_6 && io_B_Valid_6_delay_3);
  assign pE_95_valid = (io_A_Valid_3_delay_7 && io_B_Valid_7_delay_3);
  assign pE_96_valid = (io_A_Valid_4 && io_B_Valid_0_delay_4);
  assign pE_97_valid = (io_A_Valid_4_delay_1 && io_B_Valid_1_delay_4);
  assign pE_98_valid = (io_A_Valid_4_delay_2 && io_B_Valid_2_delay_4);
  assign pE_99_valid = (io_A_Valid_4_delay_3 && io_B_Valid_3_delay_4);
  assign pE_100_valid = (io_A_Valid_4_delay_4 && io_B_Valid_4_delay_4);
  assign pE_101_valid = (io_A_Valid_4_delay_5 && io_B_Valid_5_delay_4);
  assign pE_102_valid = (io_A_Valid_4_delay_6 && io_B_Valid_6_delay_4);
  assign pE_103_valid = (io_A_Valid_4_delay_7 && io_B_Valid_7_delay_4);
  assign pE_104_valid = (io_A_Valid_5 && io_B_Valid_0_delay_5);
  assign pE_105_valid = (io_A_Valid_5_delay_1 && io_B_Valid_1_delay_5);
  assign pE_106_valid = (io_A_Valid_5_delay_2 && io_B_Valid_2_delay_5);
  assign pE_107_valid = (io_A_Valid_5_delay_3 && io_B_Valid_3_delay_5);
  assign pE_108_valid = (io_A_Valid_5_delay_4 && io_B_Valid_4_delay_5);
  assign pE_109_valid = (io_A_Valid_5_delay_5 && io_B_Valid_5_delay_5);
  assign pE_110_valid = (io_A_Valid_5_delay_6 && io_B_Valid_6_delay_5);
  assign pE_111_valid = (io_A_Valid_5_delay_7 && io_B_Valid_7_delay_5);
  assign pE_112_valid = (io_A_Valid_6 && io_B_Valid_0_delay_6);
  assign pE_113_valid = (io_A_Valid_6_delay_1 && io_B_Valid_1_delay_6);
  assign pE_114_valid = (io_A_Valid_6_delay_2 && io_B_Valid_2_delay_6);
  assign pE_115_valid = (io_A_Valid_6_delay_3 && io_B_Valid_3_delay_6);
  assign pE_116_valid = (io_A_Valid_6_delay_4 && io_B_Valid_4_delay_6);
  assign pE_117_valid = (io_A_Valid_6_delay_5 && io_B_Valid_5_delay_6);
  assign pE_118_valid = (io_A_Valid_6_delay_6 && io_B_Valid_6_delay_6);
  assign pE_119_valid = (io_A_Valid_6_delay_7 && io_B_Valid_7_delay_6);
  assign pE_120_valid = (io_A_Valid_7 && io_B_Valid_0_delay_7);
  assign pE_121_valid = (io_A_Valid_7_delay_1 && io_B_Valid_1_delay_7);
  assign pE_122_valid = (io_A_Valid_7_delay_2 && io_B_Valid_2_delay_7);
  assign pE_123_valid = (io_A_Valid_7_delay_3 && io_B_Valid_3_delay_7);
  assign pE_124_valid = (io_A_Valid_7_delay_4 && io_B_Valid_4_delay_7);
  assign pE_125_valid = (io_A_Valid_7_delay_5 && io_B_Valid_5_delay_7);
  assign pE_126_valid = (io_A_Valid_7_delay_6 && io_B_Valid_6_delay_7);
  assign pE_127_valid = (io_A_Valid_7_delay_7 && io_B_Valid_7_delay_7);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      io_signCount_regNextWhen <= 16'h0;
      io_signCount_regNextWhen_1 <= 16'h0;
      io_signCount_regNextWhen_2 <= 16'h0;
      io_signCount_regNextWhen_3 <= 16'h0;
      io_signCount_regNextWhen_4 <= 16'h0;
      io_signCount_regNextWhen_5 <= 16'h0;
      io_signCount_regNextWhen_6 <= 16'h0;
      io_signCount_regNextWhen_7 <= 16'h0;
    end else begin
      if(start) begin
        io_signCount_regNextWhen <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_1 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_2 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_3 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_4 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_5 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_6 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_7 <= io_signCount;
      end
    end
  end

  always @(posedge clk) begin
    io_A_Valid_0_delay_1 <= io_A_Valid_0;
    io_A_Valid_0_delay_1_1 <= io_A_Valid_0;
    io_A_Valid_0_delay_2 <= io_A_Valid_0_delay_1_1;
    io_A_Valid_0_delay_1_2 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_1 <= io_A_Valid_0_delay_1_2;
    io_A_Valid_0_delay_3 <= io_A_Valid_0_delay_2_1;
    io_A_Valid_0_delay_1_3 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_2 <= io_A_Valid_0_delay_1_3;
    io_A_Valid_0_delay_3_1 <= io_A_Valid_0_delay_2_2;
    io_A_Valid_0_delay_4 <= io_A_Valid_0_delay_3_1;
    io_A_Valid_0_delay_1_4 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_3 <= io_A_Valid_0_delay_1_4;
    io_A_Valid_0_delay_3_2 <= io_A_Valid_0_delay_2_3;
    io_A_Valid_0_delay_4_1 <= io_A_Valid_0_delay_3_2;
    io_A_Valid_0_delay_5 <= io_A_Valid_0_delay_4_1;
    io_A_Valid_0_delay_1_5 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_4 <= io_A_Valid_0_delay_1_5;
    io_A_Valid_0_delay_3_3 <= io_A_Valid_0_delay_2_4;
    io_A_Valid_0_delay_4_2 <= io_A_Valid_0_delay_3_3;
    io_A_Valid_0_delay_5_1 <= io_A_Valid_0_delay_4_2;
    io_A_Valid_0_delay_6 <= io_A_Valid_0_delay_5_1;
    io_A_Valid_0_delay_1_6 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_5 <= io_A_Valid_0_delay_1_6;
    io_A_Valid_0_delay_3_4 <= io_A_Valid_0_delay_2_5;
    io_A_Valid_0_delay_4_3 <= io_A_Valid_0_delay_3_4;
    io_A_Valid_0_delay_5_2 <= io_A_Valid_0_delay_4_3;
    io_A_Valid_0_delay_6_1 <= io_A_Valid_0_delay_5_2;
    io_A_Valid_0_delay_7 <= io_A_Valid_0_delay_6_1;
    io_B_Valid_0_delay_1 <= io_B_Valid_0;
    io_A_Valid_1_delay_1 <= io_A_Valid_1;
    io_B_Valid_1_delay_1 <= io_B_Valid_1;
    io_A_Valid_1_delay_1_1 <= io_A_Valid_1;
    io_A_Valid_1_delay_2 <= io_A_Valid_1_delay_1_1;
    io_B_Valid_2_delay_1 <= io_B_Valid_2;
    io_A_Valid_1_delay_1_2 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_1 <= io_A_Valid_1_delay_1_2;
    io_A_Valid_1_delay_3 <= io_A_Valid_1_delay_2_1;
    io_B_Valid_3_delay_1 <= io_B_Valid_3;
    io_A_Valid_1_delay_1_3 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_2 <= io_A_Valid_1_delay_1_3;
    io_A_Valid_1_delay_3_1 <= io_A_Valid_1_delay_2_2;
    io_A_Valid_1_delay_4 <= io_A_Valid_1_delay_3_1;
    io_B_Valid_4_delay_1 <= io_B_Valid_4;
    io_A_Valid_1_delay_1_4 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_3 <= io_A_Valid_1_delay_1_4;
    io_A_Valid_1_delay_3_2 <= io_A_Valid_1_delay_2_3;
    io_A_Valid_1_delay_4_1 <= io_A_Valid_1_delay_3_2;
    io_A_Valid_1_delay_5 <= io_A_Valid_1_delay_4_1;
    io_B_Valid_5_delay_1 <= io_B_Valid_5;
    io_A_Valid_1_delay_1_5 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_4 <= io_A_Valid_1_delay_1_5;
    io_A_Valid_1_delay_3_3 <= io_A_Valid_1_delay_2_4;
    io_A_Valid_1_delay_4_2 <= io_A_Valid_1_delay_3_3;
    io_A_Valid_1_delay_5_1 <= io_A_Valid_1_delay_4_2;
    io_A_Valid_1_delay_6 <= io_A_Valid_1_delay_5_1;
    io_B_Valid_6_delay_1 <= io_B_Valid_6;
    io_A_Valid_1_delay_1_6 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_5 <= io_A_Valid_1_delay_1_6;
    io_A_Valid_1_delay_3_4 <= io_A_Valid_1_delay_2_5;
    io_A_Valid_1_delay_4_3 <= io_A_Valid_1_delay_3_4;
    io_A_Valid_1_delay_5_2 <= io_A_Valid_1_delay_4_3;
    io_A_Valid_1_delay_6_1 <= io_A_Valid_1_delay_5_2;
    io_A_Valid_1_delay_7 <= io_A_Valid_1_delay_6_1;
    io_B_Valid_7_delay_1 <= io_B_Valid_7;
    io_B_Valid_0_delay_1_1 <= io_B_Valid_0;
    io_B_Valid_0_delay_2 <= io_B_Valid_0_delay_1_1;
    io_A_Valid_2_delay_1 <= io_A_Valid_2;
    io_B_Valid_1_delay_1_1 <= io_B_Valid_1;
    io_B_Valid_1_delay_2 <= io_B_Valid_1_delay_1_1;
    io_A_Valid_2_delay_1_1 <= io_A_Valid_2;
    io_A_Valid_2_delay_2 <= io_A_Valid_2_delay_1_1;
    io_B_Valid_2_delay_1_1 <= io_B_Valid_2;
    io_B_Valid_2_delay_2 <= io_B_Valid_2_delay_1_1;
    io_A_Valid_2_delay_1_2 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_1 <= io_A_Valid_2_delay_1_2;
    io_A_Valid_2_delay_3 <= io_A_Valid_2_delay_2_1;
    io_B_Valid_3_delay_1_1 <= io_B_Valid_3;
    io_B_Valid_3_delay_2 <= io_B_Valid_3_delay_1_1;
    io_A_Valid_2_delay_1_3 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_2 <= io_A_Valid_2_delay_1_3;
    io_A_Valid_2_delay_3_1 <= io_A_Valid_2_delay_2_2;
    io_A_Valid_2_delay_4 <= io_A_Valid_2_delay_3_1;
    io_B_Valid_4_delay_1_1 <= io_B_Valid_4;
    io_B_Valid_4_delay_2 <= io_B_Valid_4_delay_1_1;
    io_A_Valid_2_delay_1_4 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_3 <= io_A_Valid_2_delay_1_4;
    io_A_Valid_2_delay_3_2 <= io_A_Valid_2_delay_2_3;
    io_A_Valid_2_delay_4_1 <= io_A_Valid_2_delay_3_2;
    io_A_Valid_2_delay_5 <= io_A_Valid_2_delay_4_1;
    io_B_Valid_5_delay_1_1 <= io_B_Valid_5;
    io_B_Valid_5_delay_2 <= io_B_Valid_5_delay_1_1;
    io_A_Valid_2_delay_1_5 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_4 <= io_A_Valid_2_delay_1_5;
    io_A_Valid_2_delay_3_3 <= io_A_Valid_2_delay_2_4;
    io_A_Valid_2_delay_4_2 <= io_A_Valid_2_delay_3_3;
    io_A_Valid_2_delay_5_1 <= io_A_Valid_2_delay_4_2;
    io_A_Valid_2_delay_6 <= io_A_Valid_2_delay_5_1;
    io_B_Valid_6_delay_1_1 <= io_B_Valid_6;
    io_B_Valid_6_delay_2 <= io_B_Valid_6_delay_1_1;
    io_A_Valid_2_delay_1_6 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_5 <= io_A_Valid_2_delay_1_6;
    io_A_Valid_2_delay_3_4 <= io_A_Valid_2_delay_2_5;
    io_A_Valid_2_delay_4_3 <= io_A_Valid_2_delay_3_4;
    io_A_Valid_2_delay_5_2 <= io_A_Valid_2_delay_4_3;
    io_A_Valid_2_delay_6_1 <= io_A_Valid_2_delay_5_2;
    io_A_Valid_2_delay_7 <= io_A_Valid_2_delay_6_1;
    io_B_Valid_7_delay_1_1 <= io_B_Valid_7;
    io_B_Valid_7_delay_2 <= io_B_Valid_7_delay_1_1;
    io_B_Valid_0_delay_1_2 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_1 <= io_B_Valid_0_delay_1_2;
    io_B_Valid_0_delay_3 <= io_B_Valid_0_delay_2_1;
    io_A_Valid_3_delay_1 <= io_A_Valid_3;
    io_B_Valid_1_delay_1_2 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_1 <= io_B_Valid_1_delay_1_2;
    io_B_Valid_1_delay_3 <= io_B_Valid_1_delay_2_1;
    io_A_Valid_3_delay_1_1 <= io_A_Valid_3;
    io_A_Valid_3_delay_2 <= io_A_Valid_3_delay_1_1;
    io_B_Valid_2_delay_1_2 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_1 <= io_B_Valid_2_delay_1_2;
    io_B_Valid_2_delay_3 <= io_B_Valid_2_delay_2_1;
    io_A_Valid_3_delay_1_2 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_1 <= io_A_Valid_3_delay_1_2;
    io_A_Valid_3_delay_3 <= io_A_Valid_3_delay_2_1;
    io_B_Valid_3_delay_1_2 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_1 <= io_B_Valid_3_delay_1_2;
    io_B_Valid_3_delay_3 <= io_B_Valid_3_delay_2_1;
    io_A_Valid_3_delay_1_3 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_2 <= io_A_Valid_3_delay_1_3;
    io_A_Valid_3_delay_3_1 <= io_A_Valid_3_delay_2_2;
    io_A_Valid_3_delay_4 <= io_A_Valid_3_delay_3_1;
    io_B_Valid_4_delay_1_2 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_1 <= io_B_Valid_4_delay_1_2;
    io_B_Valid_4_delay_3 <= io_B_Valid_4_delay_2_1;
    io_A_Valid_3_delay_1_4 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_3 <= io_A_Valid_3_delay_1_4;
    io_A_Valid_3_delay_3_2 <= io_A_Valid_3_delay_2_3;
    io_A_Valid_3_delay_4_1 <= io_A_Valid_3_delay_3_2;
    io_A_Valid_3_delay_5 <= io_A_Valid_3_delay_4_1;
    io_B_Valid_5_delay_1_2 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_1 <= io_B_Valid_5_delay_1_2;
    io_B_Valid_5_delay_3 <= io_B_Valid_5_delay_2_1;
    io_A_Valid_3_delay_1_5 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_4 <= io_A_Valid_3_delay_1_5;
    io_A_Valid_3_delay_3_3 <= io_A_Valid_3_delay_2_4;
    io_A_Valid_3_delay_4_2 <= io_A_Valid_3_delay_3_3;
    io_A_Valid_3_delay_5_1 <= io_A_Valid_3_delay_4_2;
    io_A_Valid_3_delay_6 <= io_A_Valid_3_delay_5_1;
    io_B_Valid_6_delay_1_2 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_1 <= io_B_Valid_6_delay_1_2;
    io_B_Valid_6_delay_3 <= io_B_Valid_6_delay_2_1;
    io_A_Valid_3_delay_1_6 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_5 <= io_A_Valid_3_delay_1_6;
    io_A_Valid_3_delay_3_4 <= io_A_Valid_3_delay_2_5;
    io_A_Valid_3_delay_4_3 <= io_A_Valid_3_delay_3_4;
    io_A_Valid_3_delay_5_2 <= io_A_Valid_3_delay_4_3;
    io_A_Valid_3_delay_6_1 <= io_A_Valid_3_delay_5_2;
    io_A_Valid_3_delay_7 <= io_A_Valid_3_delay_6_1;
    io_B_Valid_7_delay_1_2 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_1 <= io_B_Valid_7_delay_1_2;
    io_B_Valid_7_delay_3 <= io_B_Valid_7_delay_2_1;
    io_B_Valid_0_delay_1_3 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_2 <= io_B_Valid_0_delay_1_3;
    io_B_Valid_0_delay_3_1 <= io_B_Valid_0_delay_2_2;
    io_B_Valid_0_delay_4 <= io_B_Valid_0_delay_3_1;
    io_A_Valid_4_delay_1 <= io_A_Valid_4;
    io_B_Valid_1_delay_1_3 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_2 <= io_B_Valid_1_delay_1_3;
    io_B_Valid_1_delay_3_1 <= io_B_Valid_1_delay_2_2;
    io_B_Valid_1_delay_4 <= io_B_Valid_1_delay_3_1;
    io_A_Valid_4_delay_1_1 <= io_A_Valid_4;
    io_A_Valid_4_delay_2 <= io_A_Valid_4_delay_1_1;
    io_B_Valid_2_delay_1_3 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_2 <= io_B_Valid_2_delay_1_3;
    io_B_Valid_2_delay_3_1 <= io_B_Valid_2_delay_2_2;
    io_B_Valid_2_delay_4 <= io_B_Valid_2_delay_3_1;
    io_A_Valid_4_delay_1_2 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_1 <= io_A_Valid_4_delay_1_2;
    io_A_Valid_4_delay_3 <= io_A_Valid_4_delay_2_1;
    io_B_Valid_3_delay_1_3 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_2 <= io_B_Valid_3_delay_1_3;
    io_B_Valid_3_delay_3_1 <= io_B_Valid_3_delay_2_2;
    io_B_Valid_3_delay_4 <= io_B_Valid_3_delay_3_1;
    io_A_Valid_4_delay_1_3 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_2 <= io_A_Valid_4_delay_1_3;
    io_A_Valid_4_delay_3_1 <= io_A_Valid_4_delay_2_2;
    io_A_Valid_4_delay_4 <= io_A_Valid_4_delay_3_1;
    io_B_Valid_4_delay_1_3 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_2 <= io_B_Valid_4_delay_1_3;
    io_B_Valid_4_delay_3_1 <= io_B_Valid_4_delay_2_2;
    io_B_Valid_4_delay_4 <= io_B_Valid_4_delay_3_1;
    io_A_Valid_4_delay_1_4 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_3 <= io_A_Valid_4_delay_1_4;
    io_A_Valid_4_delay_3_2 <= io_A_Valid_4_delay_2_3;
    io_A_Valid_4_delay_4_1 <= io_A_Valid_4_delay_3_2;
    io_A_Valid_4_delay_5 <= io_A_Valid_4_delay_4_1;
    io_B_Valid_5_delay_1_3 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_2 <= io_B_Valid_5_delay_1_3;
    io_B_Valid_5_delay_3_1 <= io_B_Valid_5_delay_2_2;
    io_B_Valid_5_delay_4 <= io_B_Valid_5_delay_3_1;
    io_A_Valid_4_delay_1_5 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_4 <= io_A_Valid_4_delay_1_5;
    io_A_Valid_4_delay_3_3 <= io_A_Valid_4_delay_2_4;
    io_A_Valid_4_delay_4_2 <= io_A_Valid_4_delay_3_3;
    io_A_Valid_4_delay_5_1 <= io_A_Valid_4_delay_4_2;
    io_A_Valid_4_delay_6 <= io_A_Valid_4_delay_5_1;
    io_B_Valid_6_delay_1_3 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_2 <= io_B_Valid_6_delay_1_3;
    io_B_Valid_6_delay_3_1 <= io_B_Valid_6_delay_2_2;
    io_B_Valid_6_delay_4 <= io_B_Valid_6_delay_3_1;
    io_A_Valid_4_delay_1_6 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_5 <= io_A_Valid_4_delay_1_6;
    io_A_Valid_4_delay_3_4 <= io_A_Valid_4_delay_2_5;
    io_A_Valid_4_delay_4_3 <= io_A_Valid_4_delay_3_4;
    io_A_Valid_4_delay_5_2 <= io_A_Valid_4_delay_4_3;
    io_A_Valid_4_delay_6_1 <= io_A_Valid_4_delay_5_2;
    io_A_Valid_4_delay_7 <= io_A_Valid_4_delay_6_1;
    io_B_Valid_7_delay_1_3 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_2 <= io_B_Valid_7_delay_1_3;
    io_B_Valid_7_delay_3_1 <= io_B_Valid_7_delay_2_2;
    io_B_Valid_7_delay_4 <= io_B_Valid_7_delay_3_1;
    io_B_Valid_0_delay_1_4 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_3 <= io_B_Valid_0_delay_1_4;
    io_B_Valid_0_delay_3_2 <= io_B_Valid_0_delay_2_3;
    io_B_Valid_0_delay_4_1 <= io_B_Valid_0_delay_3_2;
    io_B_Valid_0_delay_5 <= io_B_Valid_0_delay_4_1;
    io_A_Valid_5_delay_1 <= io_A_Valid_5;
    io_B_Valid_1_delay_1_4 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_3 <= io_B_Valid_1_delay_1_4;
    io_B_Valid_1_delay_3_2 <= io_B_Valid_1_delay_2_3;
    io_B_Valid_1_delay_4_1 <= io_B_Valid_1_delay_3_2;
    io_B_Valid_1_delay_5 <= io_B_Valid_1_delay_4_1;
    io_A_Valid_5_delay_1_1 <= io_A_Valid_5;
    io_A_Valid_5_delay_2 <= io_A_Valid_5_delay_1_1;
    io_B_Valid_2_delay_1_4 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_3 <= io_B_Valid_2_delay_1_4;
    io_B_Valid_2_delay_3_2 <= io_B_Valid_2_delay_2_3;
    io_B_Valid_2_delay_4_1 <= io_B_Valid_2_delay_3_2;
    io_B_Valid_2_delay_5 <= io_B_Valid_2_delay_4_1;
    io_A_Valid_5_delay_1_2 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_1 <= io_A_Valid_5_delay_1_2;
    io_A_Valid_5_delay_3 <= io_A_Valid_5_delay_2_1;
    io_B_Valid_3_delay_1_4 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_3 <= io_B_Valid_3_delay_1_4;
    io_B_Valid_3_delay_3_2 <= io_B_Valid_3_delay_2_3;
    io_B_Valid_3_delay_4_1 <= io_B_Valid_3_delay_3_2;
    io_B_Valid_3_delay_5 <= io_B_Valid_3_delay_4_1;
    io_A_Valid_5_delay_1_3 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_2 <= io_A_Valid_5_delay_1_3;
    io_A_Valid_5_delay_3_1 <= io_A_Valid_5_delay_2_2;
    io_A_Valid_5_delay_4 <= io_A_Valid_5_delay_3_1;
    io_B_Valid_4_delay_1_4 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_3 <= io_B_Valid_4_delay_1_4;
    io_B_Valid_4_delay_3_2 <= io_B_Valid_4_delay_2_3;
    io_B_Valid_4_delay_4_1 <= io_B_Valid_4_delay_3_2;
    io_B_Valid_4_delay_5 <= io_B_Valid_4_delay_4_1;
    io_A_Valid_5_delay_1_4 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_3 <= io_A_Valid_5_delay_1_4;
    io_A_Valid_5_delay_3_2 <= io_A_Valid_5_delay_2_3;
    io_A_Valid_5_delay_4_1 <= io_A_Valid_5_delay_3_2;
    io_A_Valid_5_delay_5 <= io_A_Valid_5_delay_4_1;
    io_B_Valid_5_delay_1_4 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_3 <= io_B_Valid_5_delay_1_4;
    io_B_Valid_5_delay_3_2 <= io_B_Valid_5_delay_2_3;
    io_B_Valid_5_delay_4_1 <= io_B_Valid_5_delay_3_2;
    io_B_Valid_5_delay_5 <= io_B_Valid_5_delay_4_1;
    io_A_Valid_5_delay_1_5 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_4 <= io_A_Valid_5_delay_1_5;
    io_A_Valid_5_delay_3_3 <= io_A_Valid_5_delay_2_4;
    io_A_Valid_5_delay_4_2 <= io_A_Valid_5_delay_3_3;
    io_A_Valid_5_delay_5_1 <= io_A_Valid_5_delay_4_2;
    io_A_Valid_5_delay_6 <= io_A_Valid_5_delay_5_1;
    io_B_Valid_6_delay_1_4 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_3 <= io_B_Valid_6_delay_1_4;
    io_B_Valid_6_delay_3_2 <= io_B_Valid_6_delay_2_3;
    io_B_Valid_6_delay_4_1 <= io_B_Valid_6_delay_3_2;
    io_B_Valid_6_delay_5 <= io_B_Valid_6_delay_4_1;
    io_A_Valid_5_delay_1_6 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_5 <= io_A_Valid_5_delay_1_6;
    io_A_Valid_5_delay_3_4 <= io_A_Valid_5_delay_2_5;
    io_A_Valid_5_delay_4_3 <= io_A_Valid_5_delay_3_4;
    io_A_Valid_5_delay_5_2 <= io_A_Valid_5_delay_4_3;
    io_A_Valid_5_delay_6_1 <= io_A_Valid_5_delay_5_2;
    io_A_Valid_5_delay_7 <= io_A_Valid_5_delay_6_1;
    io_B_Valid_7_delay_1_4 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_3 <= io_B_Valid_7_delay_1_4;
    io_B_Valid_7_delay_3_2 <= io_B_Valid_7_delay_2_3;
    io_B_Valid_7_delay_4_1 <= io_B_Valid_7_delay_3_2;
    io_B_Valid_7_delay_5 <= io_B_Valid_7_delay_4_1;
    io_B_Valid_0_delay_1_5 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_4 <= io_B_Valid_0_delay_1_5;
    io_B_Valid_0_delay_3_3 <= io_B_Valid_0_delay_2_4;
    io_B_Valid_0_delay_4_2 <= io_B_Valid_0_delay_3_3;
    io_B_Valid_0_delay_5_1 <= io_B_Valid_0_delay_4_2;
    io_B_Valid_0_delay_6 <= io_B_Valid_0_delay_5_1;
    io_A_Valid_6_delay_1 <= io_A_Valid_6;
    io_B_Valid_1_delay_1_5 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_4 <= io_B_Valid_1_delay_1_5;
    io_B_Valid_1_delay_3_3 <= io_B_Valid_1_delay_2_4;
    io_B_Valid_1_delay_4_2 <= io_B_Valid_1_delay_3_3;
    io_B_Valid_1_delay_5_1 <= io_B_Valid_1_delay_4_2;
    io_B_Valid_1_delay_6 <= io_B_Valid_1_delay_5_1;
    io_A_Valid_6_delay_1_1 <= io_A_Valid_6;
    io_A_Valid_6_delay_2 <= io_A_Valid_6_delay_1_1;
    io_B_Valid_2_delay_1_5 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_4 <= io_B_Valid_2_delay_1_5;
    io_B_Valid_2_delay_3_3 <= io_B_Valid_2_delay_2_4;
    io_B_Valid_2_delay_4_2 <= io_B_Valid_2_delay_3_3;
    io_B_Valid_2_delay_5_1 <= io_B_Valid_2_delay_4_2;
    io_B_Valid_2_delay_6 <= io_B_Valid_2_delay_5_1;
    io_A_Valid_6_delay_1_2 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_1 <= io_A_Valid_6_delay_1_2;
    io_A_Valid_6_delay_3 <= io_A_Valid_6_delay_2_1;
    io_B_Valid_3_delay_1_5 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_4 <= io_B_Valid_3_delay_1_5;
    io_B_Valid_3_delay_3_3 <= io_B_Valid_3_delay_2_4;
    io_B_Valid_3_delay_4_2 <= io_B_Valid_3_delay_3_3;
    io_B_Valid_3_delay_5_1 <= io_B_Valid_3_delay_4_2;
    io_B_Valid_3_delay_6 <= io_B_Valid_3_delay_5_1;
    io_A_Valid_6_delay_1_3 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_2 <= io_A_Valid_6_delay_1_3;
    io_A_Valid_6_delay_3_1 <= io_A_Valid_6_delay_2_2;
    io_A_Valid_6_delay_4 <= io_A_Valid_6_delay_3_1;
    io_B_Valid_4_delay_1_5 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_4 <= io_B_Valid_4_delay_1_5;
    io_B_Valid_4_delay_3_3 <= io_B_Valid_4_delay_2_4;
    io_B_Valid_4_delay_4_2 <= io_B_Valid_4_delay_3_3;
    io_B_Valid_4_delay_5_1 <= io_B_Valid_4_delay_4_2;
    io_B_Valid_4_delay_6 <= io_B_Valid_4_delay_5_1;
    io_A_Valid_6_delay_1_4 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_3 <= io_A_Valid_6_delay_1_4;
    io_A_Valid_6_delay_3_2 <= io_A_Valid_6_delay_2_3;
    io_A_Valid_6_delay_4_1 <= io_A_Valid_6_delay_3_2;
    io_A_Valid_6_delay_5 <= io_A_Valid_6_delay_4_1;
    io_B_Valid_5_delay_1_5 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_4 <= io_B_Valid_5_delay_1_5;
    io_B_Valid_5_delay_3_3 <= io_B_Valid_5_delay_2_4;
    io_B_Valid_5_delay_4_2 <= io_B_Valid_5_delay_3_3;
    io_B_Valid_5_delay_5_1 <= io_B_Valid_5_delay_4_2;
    io_B_Valid_5_delay_6 <= io_B_Valid_5_delay_5_1;
    io_A_Valid_6_delay_1_5 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_4 <= io_A_Valid_6_delay_1_5;
    io_A_Valid_6_delay_3_3 <= io_A_Valid_6_delay_2_4;
    io_A_Valid_6_delay_4_2 <= io_A_Valid_6_delay_3_3;
    io_A_Valid_6_delay_5_1 <= io_A_Valid_6_delay_4_2;
    io_A_Valid_6_delay_6 <= io_A_Valid_6_delay_5_1;
    io_B_Valid_6_delay_1_5 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_4 <= io_B_Valid_6_delay_1_5;
    io_B_Valid_6_delay_3_3 <= io_B_Valid_6_delay_2_4;
    io_B_Valid_6_delay_4_2 <= io_B_Valid_6_delay_3_3;
    io_B_Valid_6_delay_5_1 <= io_B_Valid_6_delay_4_2;
    io_B_Valid_6_delay_6 <= io_B_Valid_6_delay_5_1;
    io_A_Valid_6_delay_1_6 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_5 <= io_A_Valid_6_delay_1_6;
    io_A_Valid_6_delay_3_4 <= io_A_Valid_6_delay_2_5;
    io_A_Valid_6_delay_4_3 <= io_A_Valid_6_delay_3_4;
    io_A_Valid_6_delay_5_2 <= io_A_Valid_6_delay_4_3;
    io_A_Valid_6_delay_6_1 <= io_A_Valid_6_delay_5_2;
    io_A_Valid_6_delay_7 <= io_A_Valid_6_delay_6_1;
    io_B_Valid_7_delay_1_5 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_4 <= io_B_Valid_7_delay_1_5;
    io_B_Valid_7_delay_3_3 <= io_B_Valid_7_delay_2_4;
    io_B_Valid_7_delay_4_2 <= io_B_Valid_7_delay_3_3;
    io_B_Valid_7_delay_5_1 <= io_B_Valid_7_delay_4_2;
    io_B_Valid_7_delay_6 <= io_B_Valid_7_delay_5_1;
    io_B_Valid_0_delay_1_6 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_5 <= io_B_Valid_0_delay_1_6;
    io_B_Valid_0_delay_3_4 <= io_B_Valid_0_delay_2_5;
    io_B_Valid_0_delay_4_3 <= io_B_Valid_0_delay_3_4;
    io_B_Valid_0_delay_5_2 <= io_B_Valid_0_delay_4_3;
    io_B_Valid_0_delay_6_1 <= io_B_Valid_0_delay_5_2;
    io_B_Valid_0_delay_7 <= io_B_Valid_0_delay_6_1;
    io_A_Valid_7_delay_1 <= io_A_Valid_7;
    io_B_Valid_1_delay_1_6 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_5 <= io_B_Valid_1_delay_1_6;
    io_B_Valid_1_delay_3_4 <= io_B_Valid_1_delay_2_5;
    io_B_Valid_1_delay_4_3 <= io_B_Valid_1_delay_3_4;
    io_B_Valid_1_delay_5_2 <= io_B_Valid_1_delay_4_3;
    io_B_Valid_1_delay_6_1 <= io_B_Valid_1_delay_5_2;
    io_B_Valid_1_delay_7 <= io_B_Valid_1_delay_6_1;
    io_A_Valid_7_delay_1_1 <= io_A_Valid_7;
    io_A_Valid_7_delay_2 <= io_A_Valid_7_delay_1_1;
    io_B_Valid_2_delay_1_6 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_5 <= io_B_Valid_2_delay_1_6;
    io_B_Valid_2_delay_3_4 <= io_B_Valid_2_delay_2_5;
    io_B_Valid_2_delay_4_3 <= io_B_Valid_2_delay_3_4;
    io_B_Valid_2_delay_5_2 <= io_B_Valid_2_delay_4_3;
    io_B_Valid_2_delay_6_1 <= io_B_Valid_2_delay_5_2;
    io_B_Valid_2_delay_7 <= io_B_Valid_2_delay_6_1;
    io_A_Valid_7_delay_1_2 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_1 <= io_A_Valid_7_delay_1_2;
    io_A_Valid_7_delay_3 <= io_A_Valid_7_delay_2_1;
    io_B_Valid_3_delay_1_6 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_5 <= io_B_Valid_3_delay_1_6;
    io_B_Valid_3_delay_3_4 <= io_B_Valid_3_delay_2_5;
    io_B_Valid_3_delay_4_3 <= io_B_Valid_3_delay_3_4;
    io_B_Valid_3_delay_5_2 <= io_B_Valid_3_delay_4_3;
    io_B_Valid_3_delay_6_1 <= io_B_Valid_3_delay_5_2;
    io_B_Valid_3_delay_7 <= io_B_Valid_3_delay_6_1;
    io_A_Valid_7_delay_1_3 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_2 <= io_A_Valid_7_delay_1_3;
    io_A_Valid_7_delay_3_1 <= io_A_Valid_7_delay_2_2;
    io_A_Valid_7_delay_4 <= io_A_Valid_7_delay_3_1;
    io_B_Valid_4_delay_1_6 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_5 <= io_B_Valid_4_delay_1_6;
    io_B_Valid_4_delay_3_4 <= io_B_Valid_4_delay_2_5;
    io_B_Valid_4_delay_4_3 <= io_B_Valid_4_delay_3_4;
    io_B_Valid_4_delay_5_2 <= io_B_Valid_4_delay_4_3;
    io_B_Valid_4_delay_6_1 <= io_B_Valid_4_delay_5_2;
    io_B_Valid_4_delay_7 <= io_B_Valid_4_delay_6_1;
    io_A_Valid_7_delay_1_4 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_3 <= io_A_Valid_7_delay_1_4;
    io_A_Valid_7_delay_3_2 <= io_A_Valid_7_delay_2_3;
    io_A_Valid_7_delay_4_1 <= io_A_Valid_7_delay_3_2;
    io_A_Valid_7_delay_5 <= io_A_Valid_7_delay_4_1;
    io_B_Valid_5_delay_1_6 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_5 <= io_B_Valid_5_delay_1_6;
    io_B_Valid_5_delay_3_4 <= io_B_Valid_5_delay_2_5;
    io_B_Valid_5_delay_4_3 <= io_B_Valid_5_delay_3_4;
    io_B_Valid_5_delay_5_2 <= io_B_Valid_5_delay_4_3;
    io_B_Valid_5_delay_6_1 <= io_B_Valid_5_delay_5_2;
    io_B_Valid_5_delay_7 <= io_B_Valid_5_delay_6_1;
    io_A_Valid_7_delay_1_5 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_4 <= io_A_Valid_7_delay_1_5;
    io_A_Valid_7_delay_3_3 <= io_A_Valid_7_delay_2_4;
    io_A_Valid_7_delay_4_2 <= io_A_Valid_7_delay_3_3;
    io_A_Valid_7_delay_5_1 <= io_A_Valid_7_delay_4_2;
    io_A_Valid_7_delay_6 <= io_A_Valid_7_delay_5_1;
    io_B_Valid_6_delay_1_6 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_5 <= io_B_Valid_6_delay_1_6;
    io_B_Valid_6_delay_3_4 <= io_B_Valid_6_delay_2_5;
    io_B_Valid_6_delay_4_3 <= io_B_Valid_6_delay_3_4;
    io_B_Valid_6_delay_5_2 <= io_B_Valid_6_delay_4_3;
    io_B_Valid_6_delay_6_1 <= io_B_Valid_6_delay_5_2;
    io_B_Valid_6_delay_7 <= io_B_Valid_6_delay_6_1;
    io_A_Valid_7_delay_1_6 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_5 <= io_A_Valid_7_delay_1_6;
    io_A_Valid_7_delay_3_4 <= io_A_Valid_7_delay_2_5;
    io_A_Valid_7_delay_4_3 <= io_A_Valid_7_delay_3_4;
    io_A_Valid_7_delay_5_2 <= io_A_Valid_7_delay_4_3;
    io_A_Valid_7_delay_6_1 <= io_A_Valid_7_delay_5_2;
    io_A_Valid_7_delay_7 <= io_A_Valid_7_delay_6_1;
    io_B_Valid_7_delay_1_6 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_5 <= io_B_Valid_7_delay_1_6;
    io_B_Valid_7_delay_3_4 <= io_B_Valid_7_delay_2_5;
    io_B_Valid_7_delay_4_3 <= io_B_Valid_7_delay_3_4;
    io_B_Valid_7_delay_5_2 <= io_B_Valid_7_delay_4_3;
    io_B_Valid_7_delay_6_1 <= io_B_Valid_7_delay_5_2;
    io_B_Valid_7_delay_7 <= io_B_Valid_7_delay_6_1;
  end


endmodule

//PE_63 replaced by PE

//PE_62 replaced by PE

//PE_61 replaced by PE

//PE_60 replaced by PE

//PE_59 replaced by PE

//PE_58 replaced by PE

//PE_57 replaced by PE

//PE_56 replaced by PE

//PE_55 replaced by PE

//PE_54 replaced by PE

//PE_53 replaced by PE

//PE_52 replaced by PE

//PE_51 replaced by PE

//PE_50 replaced by PE

//PE_49 replaced by PE

//PE_48 replaced by PE

//PE_47 replaced by PE

//PE_46 replaced by PE

//PE_45 replaced by PE

//PE_44 replaced by PE

//PE_43 replaced by PE

//PE_42 replaced by PE

//PE_41 replaced by PE

//PE_40 replaced by PE

//PE_39 replaced by PE

//PE_38 replaced by PE

//PE_37 replaced by PE

//PE_36 replaced by PE

//PE_35 replaced by PE

//PE_34 replaced by PE

//PE_33 replaced by PE

//PE_32 replaced by PE

//PE_31 replaced by PE

//PE_30 replaced by PE

//PE_29 replaced by PE

//PE_28 replaced by PE

//PE_27 replaced by PE

//PE_26 replaced by PE

//PE_25 replaced by PE

//PE_24 replaced by PE

//PE_23 replaced by PE

//PE_22 replaced by PE

//PE_21 replaced by PE

//PE_20 replaced by PE

//PE_19 replaced by PE

//PE_18 replaced by PE

//PE_17 replaced by PE

//PE_16 replaced by PE

//PE_15 replaced by PE

//PE_14 replaced by PE

//PE_13 replaced by PE

//PE_12 replaced by PE

//PE_11 replaced by PE

//PE_10 replaced by PE

//PE_9 replaced by PE

//PE_8 replaced by PE

//PE_7 replaced by PE

//PE_6 replaced by PE

//PE_5 replaced by PE

//PE_4 replaced by PE

//PE_3 replaced by PE

//PE_2 replaced by PE

//PE_1 replaced by PE

module PE (
  input      [7:0]    activate,
  input      [7:0]    weight,
  input               valid,
  input      [15:0]   signCount,
  output     [7:0]    acount,
  output     [7:0]    bcount,
  output reg [31:0]   PE_OUT,
  output              finish,
  input               clk,
  input               reset
);

  wire       [15:0]   dsp_P;
  wire       [31:0]   _zz_reg1;
  wire       [31:0]   _zz_reg1_1;
  wire       [31:0]   _zz_reg1_2;
  reg        [31:0]   reg1;
  reg                 valid_regNext;
  reg                 valid_regNext_regNext;
  reg        [15:0]   finishCnt_count;
  wire                finishCnt_valid;
  reg                 valid_regNext_1;
  reg        [7:0]    activate_regNext;
  reg        [7:0]    weight_regNext;

  assign _zz_reg1 = {{16{dsp_P[15]}}, dsp_P};
  assign _zz_reg1_1 = 32'h0;
  assign _zz_reg1_2 = {{16{dsp_P[15]}}, dsp_P};
  dsp_marco dsp (
    .CLK (clk          ), //i
    .A   (activate[7:0]), //i
    .B   (weight[7:0]  ), //i
    .P   (dsp_P[15:0]  )  //o
  );
  assign finishCnt_valid = ((finishCnt_count == signCount) && valid_regNext_regNext);
  assign finish = finishCnt_valid;
  always @(*) begin
    PE_OUT = 32'h0;
    if(finishCnt_valid) begin
      PE_OUT = reg1;
    end
  end

  assign acount = activate_regNext;
  assign bcount = weight_regNext;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      reg1 <= 32'h0;
      finishCnt_count <= 16'h0;
    end else begin
      if(valid_regNext_regNext) begin
        if(finishCnt_valid) begin
          finishCnt_count <= 16'h0;
        end else begin
          finishCnt_count <= (finishCnt_count + 16'h0001);
        end
      end
      if(finishCnt_valid) begin
        reg1 <= (valid ? _zz_reg1 : _zz_reg1_1);
      end else begin
        if(valid_regNext_1) begin
          reg1 <= ($signed(_zz_reg1_2) + $signed(reg1));
        end
      end
    end
  end

  always @(posedge clk) begin
    valid_regNext <= valid;
    valid_regNext_regNext <= valid_regNext;
    valid_regNext_1 <= valid;
    activate_regNext <= activate;
    weight_regNext <= weight;
  end


endmodule
