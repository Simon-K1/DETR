// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : SA3D_Top
// Git hash  : 004d9e187bb1a9a81da41bc917389f312106aff9

`timescale 1ns/1ps

module SA3D_Top (
  input               Control_start,
  input               Control_Switch_Conv,
  input      [63:0]   s_axis_s2mm_tdata,
  input      [7:0]    s_axis_s2mm_tkeep,
  input               s_axis_s2mm_tlast,
  output              s_axis_s2mm_tready,
  input               s_axis_s2mm_tvalid,
  input      [4:0]    Img2Col_Stride,
  input      [4:0]    Img2Col_Kernel_Size,
  input      [15:0]   Img2Col_Window_Size,
  input      [15:0]   Img2Col_InFeature_Size,
  input      [15:0]   Img2Col_InFeature_Channel,
  input      [15:0]   Img2Col_OutFeature_Channel,
  input      [15:0]   Img2Col_OutFeature_Size,
  input      [12:0]   Img2Col_Sliding_Size,
  input      [15:0]   Img2Col_OutCol_Count_Times,
  input      [15:0]   Img2Col_InCol_Count_Times,
  input      [15:0]   Img2Col_OutRow_Count_Times,
  input      [15:0]   Img2Col_OutFeature_Channel_Count_Times,
  input      [15:0]   Img2Col_WeightMatrix_Row,
  input      [11:0]   Img2Col_OutMatrix_Col,
  input      [19:0]   Img2Col_OutMatrix_Row,
  input               clk,
  input               reset
);
  localparam TopCtrl_Enum_IDLE = 6'd1;
  localparam TopCtrl_Enum_INIT = 6'd2;
  localparam TopCtrl_Enum_WEIGHT_CACHE = 6'd4;
  localparam TopCtrl_Enum_RECEIVE_PICTURE = 6'd8;
  localparam TopCtrl_Enum_RECEIVE_MATRIX = 6'd16;
  localparam TopCtrl_Enum_WAIT_COMPUTE_END = 6'd32;

  reg        [1:0]    InputSwitch_Switch;
  reg                 InputSwitch_m_0_axis_mm2s_tready;
  wire                SubModule_Img2Col_start;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_0;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_0;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_7;
  wire                SubModule_SA_3D__zz_io_A_Valid_0;
  wire                SubModule_SA_3D__zz_io_A_Valid_1;
  wire                SubModule_SA_3D__zz_io_A_Valid_2;
  wire                SubModule_SA_3D__zz_io_A_Valid_3;
  wire                SubModule_SA_3D__zz_io_A_Valid_4;
  wire                SubModule_SA_3D__zz_io_A_Valid_5;
  wire                SubModule_SA_3D__zz_io_A_Valid_6;
  wire                SubModule_SA_3D__zz_io_A_Valid_7;
  wire                SubModule_SA_3D__zz_io_B_Valid_0;
  wire                SubModule_SA_3D__zz_io_B_Valid_1;
  wire                SubModule_SA_3D__zz_io_B_Valid_2;
  wire                SubModule_SA_3D__zz_io_B_Valid_3;
  wire                SubModule_SA_3D__zz_io_B_Valid_4;
  wire                SubModule_SA_3D__zz_io_B_Valid_5;
  wire                SubModule_SA_3D__zz_io_B_Valid_6;
  wire                SubModule_SA_3D__zz_io_B_Valid_7;
  wire       [15:0]   SubModule_SA_3D__zz_io_signCount;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_0_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_1_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_2_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_3_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_4_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_5_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_6_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_7_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_0_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_1_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_2_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_3_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_4_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_5_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_6_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_7_1;
  wire                SubModule_SA_3D__zz_io_A_Valid_0_1;
  wire                SubModule_SA_3D__zz_io_A_Valid_1_1;
  wire                SubModule_SA_3D__zz_io_A_Valid_2_1;
  wire                SubModule_SA_3D__zz_io_A_Valid_3_1;
  wire                SubModule_SA_3D__zz_io_A_Valid_4_1;
  wire                SubModule_SA_3D__zz_io_A_Valid_5_1;
  wire                SubModule_SA_3D__zz_io_A_Valid_6_1;
  wire                SubModule_SA_3D__zz_io_A_Valid_7_1;
  wire                SubModule_SA_3D__zz_io_B_Valid_0_1;
  wire                SubModule_SA_3D__zz_io_B_Valid_1_1;
  wire                SubModule_SA_3D__zz_io_B_Valid_2_1;
  wire                SubModule_SA_3D__zz_io_B_Valid_3_1;
  wire                SubModule_SA_3D__zz_io_B_Valid_4_1;
  wire                SubModule_SA_3D__zz_io_B_Valid_5_1;
  wire                SubModule_SA_3D__zz_io_B_Valid_6_1;
  wire                SubModule_SA_3D__zz_io_B_Valid_7_1;
  wire       [15:0]   SubModule_SA_3D__zz_io_signCount_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_0_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_1_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_2_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_3_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_4_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_5_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_6_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_7_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_0_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_1_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_2_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_3_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_4_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_5_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_6_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_7_2;
  wire                SubModule_SA_3D__zz_io_A_Valid_0_2;
  wire                SubModule_SA_3D__zz_io_A_Valid_1_2;
  wire                SubModule_SA_3D__zz_io_A_Valid_2_2;
  wire                SubModule_SA_3D__zz_io_A_Valid_3_2;
  wire                SubModule_SA_3D__zz_io_A_Valid_4_2;
  wire                SubModule_SA_3D__zz_io_A_Valid_5_2;
  wire                SubModule_SA_3D__zz_io_A_Valid_6_2;
  wire                SubModule_SA_3D__zz_io_A_Valid_7_2;
  wire                SubModule_SA_3D__zz_io_B_Valid_0_2;
  wire                SubModule_SA_3D__zz_io_B_Valid_1_2;
  wire                SubModule_SA_3D__zz_io_B_Valid_2_2;
  wire                SubModule_SA_3D__zz_io_B_Valid_3_2;
  wire                SubModule_SA_3D__zz_io_B_Valid_4_2;
  wire                SubModule_SA_3D__zz_io_B_Valid_5_2;
  wire                SubModule_SA_3D__zz_io_B_Valid_6_2;
  wire                SubModule_SA_3D__zz_io_B_Valid_7_2;
  wire       [15:0]   SubModule_SA_3D__zz_io_signCount_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_0_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_1_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_2_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_3_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_4_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_5_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_6_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_7_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_0_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_1_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_2_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_3_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_4_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_5_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_6_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_7_3;
  wire                SubModule_SA_3D__zz_io_A_Valid_0_3;
  wire                SubModule_SA_3D__zz_io_A_Valid_1_3;
  wire                SubModule_SA_3D__zz_io_A_Valid_2_3;
  wire                SubModule_SA_3D__zz_io_A_Valid_3_3;
  wire                SubModule_SA_3D__zz_io_A_Valid_4_3;
  wire                SubModule_SA_3D__zz_io_A_Valid_5_3;
  wire                SubModule_SA_3D__zz_io_A_Valid_6_3;
  wire                SubModule_SA_3D__zz_io_A_Valid_7_3;
  wire                SubModule_SA_3D__zz_io_B_Valid_0_3;
  wire                SubModule_SA_3D__zz_io_B_Valid_1_3;
  wire                SubModule_SA_3D__zz_io_B_Valid_2_3;
  wire                SubModule_SA_3D__zz_io_B_Valid_3_3;
  wire                SubModule_SA_3D__zz_io_B_Valid_4_3;
  wire                SubModule_SA_3D__zz_io_B_Valid_5_3;
  wire                SubModule_SA_3D__zz_io_B_Valid_6_3;
  wire                SubModule_SA_3D__zz_io_B_Valid_7_3;
  wire       [15:0]   SubModule_SA_3D__zz_io_signCount_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_0_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_1_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_2_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_3_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_4_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_5_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_6_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_7_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_0_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_1_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_2_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_3_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_4_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_5_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_6_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_7_4;
  wire                SubModule_SA_3D__zz_io_A_Valid_0_4;
  wire                SubModule_SA_3D__zz_io_A_Valid_1_4;
  wire                SubModule_SA_3D__zz_io_A_Valid_2_4;
  wire                SubModule_SA_3D__zz_io_A_Valid_3_4;
  wire                SubModule_SA_3D__zz_io_A_Valid_4_4;
  wire                SubModule_SA_3D__zz_io_A_Valid_5_4;
  wire                SubModule_SA_3D__zz_io_A_Valid_6_4;
  wire                SubModule_SA_3D__zz_io_A_Valid_7_4;
  wire                SubModule_SA_3D__zz_io_B_Valid_0_4;
  wire                SubModule_SA_3D__zz_io_B_Valid_1_4;
  wire                SubModule_SA_3D__zz_io_B_Valid_2_4;
  wire                SubModule_SA_3D__zz_io_B_Valid_3_4;
  wire                SubModule_SA_3D__zz_io_B_Valid_4_4;
  wire                SubModule_SA_3D__zz_io_B_Valid_5_4;
  wire                SubModule_SA_3D__zz_io_B_Valid_6_4;
  wire                SubModule_SA_3D__zz_io_B_Valid_7_4;
  wire       [15:0]   SubModule_SA_3D__zz_io_signCount_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_0_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_1_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_2_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_3_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_4_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_5_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_6_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_7_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_0_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_1_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_2_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_3_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_4_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_5_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_6_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_7_5;
  wire                SubModule_SA_3D__zz_io_A_Valid_0_5;
  wire                SubModule_SA_3D__zz_io_A_Valid_1_5;
  wire                SubModule_SA_3D__zz_io_A_Valid_2_5;
  wire                SubModule_SA_3D__zz_io_A_Valid_3_5;
  wire                SubModule_SA_3D__zz_io_A_Valid_4_5;
  wire                SubModule_SA_3D__zz_io_A_Valid_5_5;
  wire                SubModule_SA_3D__zz_io_A_Valid_6_5;
  wire                SubModule_SA_3D__zz_io_A_Valid_7_5;
  wire                SubModule_SA_3D__zz_io_B_Valid_0_5;
  wire                SubModule_SA_3D__zz_io_B_Valid_1_5;
  wire                SubModule_SA_3D__zz_io_B_Valid_2_5;
  wire                SubModule_SA_3D__zz_io_B_Valid_3_5;
  wire                SubModule_SA_3D__zz_io_B_Valid_4_5;
  wire                SubModule_SA_3D__zz_io_B_Valid_5_5;
  wire                SubModule_SA_3D__zz_io_B_Valid_6_5;
  wire                SubModule_SA_3D__zz_io_B_Valid_7_5;
  wire       [15:0]   SubModule_SA_3D__zz_io_signCount_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_0_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_1_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_2_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_3_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_4_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_5_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_6_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_7_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_0_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_1_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_2_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_3_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_4_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_5_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_6_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_7_6;
  wire                SubModule_SA_3D__zz_io_A_Valid_0_6;
  wire                SubModule_SA_3D__zz_io_A_Valid_1_6;
  wire                SubModule_SA_3D__zz_io_A_Valid_2_6;
  wire                SubModule_SA_3D__zz_io_A_Valid_3_6;
  wire                SubModule_SA_3D__zz_io_A_Valid_4_6;
  wire                SubModule_SA_3D__zz_io_A_Valid_5_6;
  wire                SubModule_SA_3D__zz_io_A_Valid_6_6;
  wire                SubModule_SA_3D__zz_io_A_Valid_7_6;
  wire                SubModule_SA_3D__zz_io_B_Valid_0_6;
  wire                SubModule_SA_3D__zz_io_B_Valid_1_6;
  wire                SubModule_SA_3D__zz_io_B_Valid_2_6;
  wire                SubModule_SA_3D__zz_io_B_Valid_3_6;
  wire                SubModule_SA_3D__zz_io_B_Valid_4_6;
  wire                SubModule_SA_3D__zz_io_B_Valid_5_6;
  wire                SubModule_SA_3D__zz_io_B_Valid_6_6;
  wire                SubModule_SA_3D__zz_io_B_Valid_7_6;
  wire       [15:0]   SubModule_SA_3D__zz_io_signCount_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_0_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_1_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_2_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_3_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_4_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_5_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_6_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_7_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_0_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_1_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_2_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_3_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_4_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_5_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_6_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_7_7;
  wire                SubModule_SA_3D__zz_io_A_Valid_0_7;
  wire                SubModule_SA_3D__zz_io_A_Valid_1_7;
  wire                SubModule_SA_3D__zz_io_A_Valid_2_7;
  wire                SubModule_SA_3D__zz_io_A_Valid_3_7;
  wire                SubModule_SA_3D__zz_io_A_Valid_4_7;
  wire                SubModule_SA_3D__zz_io_A_Valid_5_7;
  wire                SubModule_SA_3D__zz_io_A_Valid_6_7;
  wire                SubModule_SA_3D__zz_io_A_Valid_7_7;
  wire                SubModule_SA_3D__zz_io_B_Valid_0_7;
  wire                SubModule_SA_3D__zz_io_B_Valid_1_7;
  wire                SubModule_SA_3D__zz_io_B_Valid_2_7;
  wire                SubModule_SA_3D__zz_io_B_Valid_3_7;
  wire                SubModule_SA_3D__zz_io_B_Valid_4_7;
  wire                SubModule_SA_3D__zz_io_B_Valid_5_7;
  wire                SubModule_SA_3D__zz_io_B_Valid_6_7;
  wire                SubModule_SA_3D__zz_io_B_Valid_7_7;
  wire       [15:0]   SubModule_SA_3D__zz_io_signCount_7;
  wire                InputSwitch_s0_axis_s2mm_tready;
  wire       [63:0]   InputSwitch_m_0_axis_mm2s_tdata;
  wire       [7:0]    InputSwitch_m_0_axis_mm2s_tkeep;
  wire                InputSwitch_m_0_axis_mm2s_tlast;
  wire                InputSwitch_m_0_axis_mm2s_tvalid;
  wire       [63:0]   InputSwitch_m_1_axis_mm2s_tdata;
  wire       [7:0]    InputSwitch_m_1_axis_mm2s_tkeep;
  wire                InputSwitch_m_1_axis_mm2s_tlast;
  wire                InputSwitch_m_1_axis_mm2s_tvalid;
  wire       [63:0]   SubModule_Img2Col_mData;
  wire       [7:0]    SubModule_Img2Col_mValid;
  wire                SubModule_Img2Col_s_axis_s2mm_tready;
  wire                SubModule_Img2Col_Raddr_Valid;
  wire                SubModule_Img2Col_LayerEnd;
  wire                SubModule_WeightCache_s_axis_s2mm_tready;
  wire       [7:0]    SubModule_WeightCache_mData_0;
  wire       [7:0]    SubModule_WeightCache_mData_1;
  wire       [7:0]    SubModule_WeightCache_mData_2;
  wire       [7:0]    SubModule_WeightCache_mData_3;
  wire       [7:0]    SubModule_WeightCache_mData_4;
  wire       [7:0]    SubModule_WeightCache_mData_5;
  wire       [7:0]    SubModule_WeightCache_mData_6;
  wire       [7:0]    SubModule_WeightCache_mData_7;
  wire       [7:0]    SubModule_WeightCache_mData_8;
  wire       [7:0]    SubModule_WeightCache_mData_9;
  wire       [7:0]    SubModule_WeightCache_mData_10;
  wire       [7:0]    SubModule_WeightCache_mData_11;
  wire       [7:0]    SubModule_WeightCache_mData_12;
  wire       [7:0]    SubModule_WeightCache_mData_13;
  wire       [7:0]    SubModule_WeightCache_mData_14;
  wire       [7:0]    SubModule_WeightCache_mData_15;
  wire       [7:0]    SubModule_WeightCache_mData_16;
  wire       [7:0]    SubModule_WeightCache_mData_17;
  wire       [7:0]    SubModule_WeightCache_mData_18;
  wire       [7:0]    SubModule_WeightCache_mData_19;
  wire       [7:0]    SubModule_WeightCache_mData_20;
  wire       [7:0]    SubModule_WeightCache_mData_21;
  wire       [7:0]    SubModule_WeightCache_mData_22;
  wire       [7:0]    SubModule_WeightCache_mData_23;
  wire       [7:0]    SubModule_WeightCache_mData_24;
  wire       [7:0]    SubModule_WeightCache_mData_25;
  wire       [7:0]    SubModule_WeightCache_mData_26;
  wire       [7:0]    SubModule_WeightCache_mData_27;
  wire       [7:0]    SubModule_WeightCache_mData_28;
  wire       [7:0]    SubModule_WeightCache_mData_29;
  wire       [7:0]    SubModule_WeightCache_mData_30;
  wire       [7:0]    SubModule_WeightCache_mData_31;
  wire       [7:0]    SubModule_WeightCache_mData_32;
  wire       [7:0]    SubModule_WeightCache_mData_33;
  wire       [7:0]    SubModule_WeightCache_mData_34;
  wire       [7:0]    SubModule_WeightCache_mData_35;
  wire       [7:0]    SubModule_WeightCache_mData_36;
  wire       [7:0]    SubModule_WeightCache_mData_37;
  wire       [7:0]    SubModule_WeightCache_mData_38;
  wire       [7:0]    SubModule_WeightCache_mData_39;
  wire       [7:0]    SubModule_WeightCache_mData_40;
  wire       [7:0]    SubModule_WeightCache_mData_41;
  wire       [7:0]    SubModule_WeightCache_mData_42;
  wire       [7:0]    SubModule_WeightCache_mData_43;
  wire       [7:0]    SubModule_WeightCache_mData_44;
  wire       [7:0]    SubModule_WeightCache_mData_45;
  wire       [7:0]    SubModule_WeightCache_mData_46;
  wire       [7:0]    SubModule_WeightCache_mData_47;
  wire       [7:0]    SubModule_WeightCache_mData_48;
  wire       [7:0]    SubModule_WeightCache_mData_49;
  wire       [7:0]    SubModule_WeightCache_mData_50;
  wire       [7:0]    SubModule_WeightCache_mData_51;
  wire       [7:0]    SubModule_WeightCache_mData_52;
  wire       [7:0]    SubModule_WeightCache_mData_53;
  wire       [7:0]    SubModule_WeightCache_mData_54;
  wire       [7:0]    SubModule_WeightCache_mData_55;
  wire       [7:0]    SubModule_WeightCache_mData_56;
  wire       [7:0]    SubModule_WeightCache_mData_57;
  wire       [7:0]    SubModule_WeightCache_mData_58;
  wire       [7:0]    SubModule_WeightCache_mData_59;
  wire       [7:0]    SubModule_WeightCache_mData_60;
  wire       [7:0]    SubModule_WeightCache_mData_61;
  wire       [7:0]    SubModule_WeightCache_mData_62;
  wire       [7:0]    SubModule_WeightCache_mData_63;
  wire                SubModule_WeightCache_Weight_Cached;
  wire       [63:0]   SubModule_WeightCache_MatrixCol_Switch;
  reg        [5:0]    Fsm_currentState;
  reg        [5:0]    Fsm_nextState;
  wire                Fsm_Inited;
  wire                Fsm_WeightCached;
  wire                Fsm_Picture_Received;
  wire                Fsm_Matrix_Received;
  wire                Fsm_Compute_End;
  wire                Fsm_Switch_Conv;
  wire                when_SA3D_Top_l46;
  wire                when_SA3D_Top_l48;
  wire                LayerEnd;
  wire                when_WaCounter_l19;
  reg        [2:0]    InitCnt_count;
  reg                 InitCnt_valid;
  wire                when_WaCounter_l14;
  wire                when_SA3D_Top_l131;
  reg                 toplevel_SubModule_WeightCache_Weight_Cached_delay_1;
  reg                 toplevel_SubModule_WeightCache_Weight_Cached_delay_2;
  reg                 toplevel_SubModule_WeightCache_Weight_Cached_delay_3;
  reg                 _zz_start;
  reg                 _zz_start_1;
  reg                 _zz_start_2;
  `ifndef SYNTHESIS
  reg [127:0] Fsm_currentState_string;
  reg [127:0] Fsm_nextState_string;
  `endif


  Compute_DataIn_Switch InputSwitch (
    .Switch               (InputSwitch_Switch[1:0]              ), //i
    .s0_axis_s2mm_tdata   (s_axis_s2mm_tdata[63:0]              ), //i
    .s0_axis_s2mm_tkeep   (s_axis_s2mm_tkeep[7:0]               ), //i
    .s0_axis_s2mm_tlast   (s_axis_s2mm_tlast                    ), //i
    .s0_axis_s2mm_tready  (InputSwitch_s0_axis_s2mm_tready      ), //o
    .s0_axis_s2mm_tvalid  (s_axis_s2mm_tvalid                   ), //i
    .m_0_axis_mm2s_tdata  (InputSwitch_m_0_axis_mm2s_tdata[63:0]), //o
    .m_0_axis_mm2s_tkeep  (InputSwitch_m_0_axis_mm2s_tkeep[7:0] ), //o
    .m_0_axis_mm2s_tlast  (InputSwitch_m_0_axis_mm2s_tlast      ), //o
    .m_0_axis_mm2s_tready (InputSwitch_m_0_axis_mm2s_tready     ), //i
    .m_0_axis_mm2s_tvalid (InputSwitch_m_0_axis_mm2s_tvalid     ), //o
    .m_1_axis_mm2s_tdata  (InputSwitch_m_1_axis_mm2s_tdata[63:0]), //o
    .m_1_axis_mm2s_tkeep  (InputSwitch_m_1_axis_mm2s_tkeep[7:0] ), //o
    .m_1_axis_mm2s_tlast  (InputSwitch_m_1_axis_mm2s_tlast      ), //o
    .m_1_axis_mm2s_tready (SubModule_Img2Col_s_axis_s2mm_tready ), //i
    .m_1_axis_mm2s_tvalid (InputSwitch_m_1_axis_mm2s_tvalid     )  //o
  );
  Img2ColStreamV2 SubModule_Img2Col (
    .mData                          (SubModule_Img2Col_mData[63:0]               ), //o
    .mValid                         (SubModule_Img2Col_mValid[7:0]               ), //o
    .s_axis_s2mm_tdata              (InputSwitch_m_1_axis_mm2s_tdata[63:0]       ), //i
    .s_axis_s2mm_tkeep              (InputSwitch_m_1_axis_mm2s_tkeep[7:0]        ), //i
    .s_axis_s2mm_tlast              (InputSwitch_m_1_axis_mm2s_tlast             ), //i
    .s_axis_s2mm_tready             (SubModule_Img2Col_s_axis_s2mm_tready        ), //o
    .s_axis_s2mm_tvalid             (InputSwitch_m_1_axis_mm2s_tvalid            ), //i
    .start                          (SubModule_Img2Col_start                     ), //i
    .Raddr_Valid                    (SubModule_Img2Col_Raddr_Valid               ), //o
    .LayerEnd                       (SubModule_Img2Col_LayerEnd                  ), //o
    .Stride                         (Img2Col_Stride[4:0]                         ), //i
    .Kernel_Size                    (Img2Col_Kernel_Size[4:0]                    ), //i
    .Window_Size                    (Img2Col_Window_Size[15:0]                   ), //i
    .InFeature_Size                 (Img2Col_InFeature_Size[15:0]                ), //i
    .InFeature_Channel              (Img2Col_InFeature_Channel[15:0]             ), //i
    .OutFeature_Channel             (Img2Col_OutFeature_Channel[15:0]            ), //i
    .OutFeature_Size                (Img2Col_OutFeature_Size[15:0]               ), //i
    .OutCol_Count_Times             (Img2Col_OutCol_Count_Times[15:0]            ), //i
    .InCol_Count_Times              (Img2Col_InCol_Count_Times[15:0]             ), //i
    .OutRow_Count_Times             (Img2Col_OutRow_Count_Times[15:0]            ), //i
    .OutFeature_Channel_Count_Times (Img2Col_OutFeature_Channel_Count_Times[15:0]), //i
    .Sliding_Size                   (Img2Col_Sliding_Size[12:0]                  ), //i
    .clk                            (clk                                         ), //i
    .reset                          (reset                                       )  //i
  );
  SA_3D SubModule_SA_3D (
    ._zz_io_MatrixA_0   (SubModule_SA_3D__zz_io_MatrixA_0[7:0]   ), //i
    ._zz_io_MatrixA_1   (SubModule_SA_3D__zz_io_MatrixA_1[7:0]   ), //i
    ._zz_io_MatrixA_2   (SubModule_SA_3D__zz_io_MatrixA_2[7:0]   ), //i
    ._zz_io_MatrixA_3   (SubModule_SA_3D__zz_io_MatrixA_3[7:0]   ), //i
    ._zz_io_MatrixA_4   (SubModule_SA_3D__zz_io_MatrixA_4[7:0]   ), //i
    ._zz_io_MatrixA_5   (SubModule_SA_3D__zz_io_MatrixA_5[7:0]   ), //i
    ._zz_io_MatrixA_6   (SubModule_SA_3D__zz_io_MatrixA_6[7:0]   ), //i
    ._zz_io_MatrixA_7   (SubModule_SA_3D__zz_io_MatrixA_7[7:0]   ), //i
    ._zz_io_MatrixB_0   (SubModule_SA_3D__zz_io_MatrixB_0[7:0]   ), //i
    ._zz_io_MatrixB_1   (SubModule_SA_3D__zz_io_MatrixB_1[7:0]   ), //i
    ._zz_io_MatrixB_2   (SubModule_SA_3D__zz_io_MatrixB_2[7:0]   ), //i
    ._zz_io_MatrixB_3   (SubModule_SA_3D__zz_io_MatrixB_3[7:0]   ), //i
    ._zz_io_MatrixB_4   (SubModule_SA_3D__zz_io_MatrixB_4[7:0]   ), //i
    ._zz_io_MatrixB_5   (SubModule_SA_3D__zz_io_MatrixB_5[7:0]   ), //i
    ._zz_io_MatrixB_6   (SubModule_SA_3D__zz_io_MatrixB_6[7:0]   ), //i
    ._zz_io_MatrixB_7   (SubModule_SA_3D__zz_io_MatrixB_7[7:0]   ), //i
    ._zz_io_A_Valid_0   (SubModule_SA_3D__zz_io_A_Valid_0        ), //i
    ._zz_io_A_Valid_1   (SubModule_SA_3D__zz_io_A_Valid_1        ), //i
    ._zz_io_A_Valid_2   (SubModule_SA_3D__zz_io_A_Valid_2        ), //i
    ._zz_io_A_Valid_3   (SubModule_SA_3D__zz_io_A_Valid_3        ), //i
    ._zz_io_A_Valid_4   (SubModule_SA_3D__zz_io_A_Valid_4        ), //i
    ._zz_io_A_Valid_5   (SubModule_SA_3D__zz_io_A_Valid_5        ), //i
    ._zz_io_A_Valid_6   (SubModule_SA_3D__zz_io_A_Valid_6        ), //i
    ._zz_io_A_Valid_7   (SubModule_SA_3D__zz_io_A_Valid_7        ), //i
    ._zz_io_B_Valid_0   (SubModule_SA_3D__zz_io_B_Valid_0        ), //i
    ._zz_io_B_Valid_1   (SubModule_SA_3D__zz_io_B_Valid_1        ), //i
    ._zz_io_B_Valid_2   (SubModule_SA_3D__zz_io_B_Valid_2        ), //i
    ._zz_io_B_Valid_3   (SubModule_SA_3D__zz_io_B_Valid_3        ), //i
    ._zz_io_B_Valid_4   (SubModule_SA_3D__zz_io_B_Valid_4        ), //i
    ._zz_io_B_Valid_5   (SubModule_SA_3D__zz_io_B_Valid_5        ), //i
    ._zz_io_B_Valid_6   (SubModule_SA_3D__zz_io_B_Valid_6        ), //i
    ._zz_io_B_Valid_7   (SubModule_SA_3D__zz_io_B_Valid_7        ), //i
    ._zz_io_signCount   (SubModule_SA_3D__zz_io_signCount[15:0]  ), //i
    .clk                (clk                                     ), //i
    ._zz_io_MatrixA_0_1 (SubModule_SA_3D__zz_io_MatrixA_0_1[7:0] ), //i
    ._zz_io_MatrixA_1_1 (SubModule_SA_3D__zz_io_MatrixA_1_1[7:0] ), //i
    ._zz_io_MatrixA_2_1 (SubModule_SA_3D__zz_io_MatrixA_2_1[7:0] ), //i
    ._zz_io_MatrixA_3_1 (SubModule_SA_3D__zz_io_MatrixA_3_1[7:0] ), //i
    ._zz_io_MatrixA_4_1 (SubModule_SA_3D__zz_io_MatrixA_4_1[7:0] ), //i
    ._zz_io_MatrixA_5_1 (SubModule_SA_3D__zz_io_MatrixA_5_1[7:0] ), //i
    ._zz_io_MatrixA_6_1 (SubModule_SA_3D__zz_io_MatrixA_6_1[7:0] ), //i
    ._zz_io_MatrixA_7_1 (SubModule_SA_3D__zz_io_MatrixA_7_1[7:0] ), //i
    ._zz_io_MatrixB_0_1 (SubModule_SA_3D__zz_io_MatrixB_0_1[7:0] ), //i
    ._zz_io_MatrixB_1_1 (SubModule_SA_3D__zz_io_MatrixB_1_1[7:0] ), //i
    ._zz_io_MatrixB_2_1 (SubModule_SA_3D__zz_io_MatrixB_2_1[7:0] ), //i
    ._zz_io_MatrixB_3_1 (SubModule_SA_3D__zz_io_MatrixB_3_1[7:0] ), //i
    ._zz_io_MatrixB_4_1 (SubModule_SA_3D__zz_io_MatrixB_4_1[7:0] ), //i
    ._zz_io_MatrixB_5_1 (SubModule_SA_3D__zz_io_MatrixB_5_1[7:0] ), //i
    ._zz_io_MatrixB_6_1 (SubModule_SA_3D__zz_io_MatrixB_6_1[7:0] ), //i
    ._zz_io_MatrixB_7_1 (SubModule_SA_3D__zz_io_MatrixB_7_1[7:0] ), //i
    ._zz_io_A_Valid_0_1 (SubModule_SA_3D__zz_io_A_Valid_0_1      ), //i
    ._zz_io_A_Valid_1_1 (SubModule_SA_3D__zz_io_A_Valid_1_1      ), //i
    ._zz_io_A_Valid_2_1 (SubModule_SA_3D__zz_io_A_Valid_2_1      ), //i
    ._zz_io_A_Valid_3_1 (SubModule_SA_3D__zz_io_A_Valid_3_1      ), //i
    ._zz_io_A_Valid_4_1 (SubModule_SA_3D__zz_io_A_Valid_4_1      ), //i
    ._zz_io_A_Valid_5_1 (SubModule_SA_3D__zz_io_A_Valid_5_1      ), //i
    ._zz_io_A_Valid_6_1 (SubModule_SA_3D__zz_io_A_Valid_6_1      ), //i
    ._zz_io_A_Valid_7_1 (SubModule_SA_3D__zz_io_A_Valid_7_1      ), //i
    ._zz_io_B_Valid_0_1 (SubModule_SA_3D__zz_io_B_Valid_0_1      ), //i
    ._zz_io_B_Valid_1_1 (SubModule_SA_3D__zz_io_B_Valid_1_1      ), //i
    ._zz_io_B_Valid_2_1 (SubModule_SA_3D__zz_io_B_Valid_2_1      ), //i
    ._zz_io_B_Valid_3_1 (SubModule_SA_3D__zz_io_B_Valid_3_1      ), //i
    ._zz_io_B_Valid_4_1 (SubModule_SA_3D__zz_io_B_Valid_4_1      ), //i
    ._zz_io_B_Valid_5_1 (SubModule_SA_3D__zz_io_B_Valid_5_1      ), //i
    ._zz_io_B_Valid_6_1 (SubModule_SA_3D__zz_io_B_Valid_6_1      ), //i
    ._zz_io_B_Valid_7_1 (SubModule_SA_3D__zz_io_B_Valid_7_1      ), //i
    ._zz_io_signCount_1 (SubModule_SA_3D__zz_io_signCount_1[15:0]), //i
    ._zz_io_MatrixA_0_2 (SubModule_SA_3D__zz_io_MatrixA_0_2[7:0] ), //i
    ._zz_io_MatrixA_1_2 (SubModule_SA_3D__zz_io_MatrixA_1_2[7:0] ), //i
    ._zz_io_MatrixA_2_2 (SubModule_SA_3D__zz_io_MatrixA_2_2[7:0] ), //i
    ._zz_io_MatrixA_3_2 (SubModule_SA_3D__zz_io_MatrixA_3_2[7:0] ), //i
    ._zz_io_MatrixA_4_2 (SubModule_SA_3D__zz_io_MatrixA_4_2[7:0] ), //i
    ._zz_io_MatrixA_5_2 (SubModule_SA_3D__zz_io_MatrixA_5_2[7:0] ), //i
    ._zz_io_MatrixA_6_2 (SubModule_SA_3D__zz_io_MatrixA_6_2[7:0] ), //i
    ._zz_io_MatrixA_7_2 (SubModule_SA_3D__zz_io_MatrixA_7_2[7:0] ), //i
    ._zz_io_MatrixB_0_2 (SubModule_SA_3D__zz_io_MatrixB_0_2[7:0] ), //i
    ._zz_io_MatrixB_1_2 (SubModule_SA_3D__zz_io_MatrixB_1_2[7:0] ), //i
    ._zz_io_MatrixB_2_2 (SubModule_SA_3D__zz_io_MatrixB_2_2[7:0] ), //i
    ._zz_io_MatrixB_3_2 (SubModule_SA_3D__zz_io_MatrixB_3_2[7:0] ), //i
    ._zz_io_MatrixB_4_2 (SubModule_SA_3D__zz_io_MatrixB_4_2[7:0] ), //i
    ._zz_io_MatrixB_5_2 (SubModule_SA_3D__zz_io_MatrixB_5_2[7:0] ), //i
    ._zz_io_MatrixB_6_2 (SubModule_SA_3D__zz_io_MatrixB_6_2[7:0] ), //i
    ._zz_io_MatrixB_7_2 (SubModule_SA_3D__zz_io_MatrixB_7_2[7:0] ), //i
    ._zz_io_A_Valid_0_2 (SubModule_SA_3D__zz_io_A_Valid_0_2      ), //i
    ._zz_io_A_Valid_1_2 (SubModule_SA_3D__zz_io_A_Valid_1_2      ), //i
    ._zz_io_A_Valid_2_2 (SubModule_SA_3D__zz_io_A_Valid_2_2      ), //i
    ._zz_io_A_Valid_3_2 (SubModule_SA_3D__zz_io_A_Valid_3_2      ), //i
    ._zz_io_A_Valid_4_2 (SubModule_SA_3D__zz_io_A_Valid_4_2      ), //i
    ._zz_io_A_Valid_5_2 (SubModule_SA_3D__zz_io_A_Valid_5_2      ), //i
    ._zz_io_A_Valid_6_2 (SubModule_SA_3D__zz_io_A_Valid_6_2      ), //i
    ._zz_io_A_Valid_7_2 (SubModule_SA_3D__zz_io_A_Valid_7_2      ), //i
    ._zz_io_B_Valid_0_2 (SubModule_SA_3D__zz_io_B_Valid_0_2      ), //i
    ._zz_io_B_Valid_1_2 (SubModule_SA_3D__zz_io_B_Valid_1_2      ), //i
    ._zz_io_B_Valid_2_2 (SubModule_SA_3D__zz_io_B_Valid_2_2      ), //i
    ._zz_io_B_Valid_3_2 (SubModule_SA_3D__zz_io_B_Valid_3_2      ), //i
    ._zz_io_B_Valid_4_2 (SubModule_SA_3D__zz_io_B_Valid_4_2      ), //i
    ._zz_io_B_Valid_5_2 (SubModule_SA_3D__zz_io_B_Valid_5_2      ), //i
    ._zz_io_B_Valid_6_2 (SubModule_SA_3D__zz_io_B_Valid_6_2      ), //i
    ._zz_io_B_Valid_7_2 (SubModule_SA_3D__zz_io_B_Valid_7_2      ), //i
    ._zz_io_signCount_2 (SubModule_SA_3D__zz_io_signCount_2[15:0]), //i
    ._zz_io_MatrixA_0_3 (SubModule_SA_3D__zz_io_MatrixA_0_3[7:0] ), //i
    ._zz_io_MatrixA_1_3 (SubModule_SA_3D__zz_io_MatrixA_1_3[7:0] ), //i
    ._zz_io_MatrixA_2_3 (SubModule_SA_3D__zz_io_MatrixA_2_3[7:0] ), //i
    ._zz_io_MatrixA_3_3 (SubModule_SA_3D__zz_io_MatrixA_3_3[7:0] ), //i
    ._zz_io_MatrixA_4_3 (SubModule_SA_3D__zz_io_MatrixA_4_3[7:0] ), //i
    ._zz_io_MatrixA_5_3 (SubModule_SA_3D__zz_io_MatrixA_5_3[7:0] ), //i
    ._zz_io_MatrixA_6_3 (SubModule_SA_3D__zz_io_MatrixA_6_3[7:0] ), //i
    ._zz_io_MatrixA_7_3 (SubModule_SA_3D__zz_io_MatrixA_7_3[7:0] ), //i
    ._zz_io_MatrixB_0_3 (SubModule_SA_3D__zz_io_MatrixB_0_3[7:0] ), //i
    ._zz_io_MatrixB_1_3 (SubModule_SA_3D__zz_io_MatrixB_1_3[7:0] ), //i
    ._zz_io_MatrixB_2_3 (SubModule_SA_3D__zz_io_MatrixB_2_3[7:0] ), //i
    ._zz_io_MatrixB_3_3 (SubModule_SA_3D__zz_io_MatrixB_3_3[7:0] ), //i
    ._zz_io_MatrixB_4_3 (SubModule_SA_3D__zz_io_MatrixB_4_3[7:0] ), //i
    ._zz_io_MatrixB_5_3 (SubModule_SA_3D__zz_io_MatrixB_5_3[7:0] ), //i
    ._zz_io_MatrixB_6_3 (SubModule_SA_3D__zz_io_MatrixB_6_3[7:0] ), //i
    ._zz_io_MatrixB_7_3 (SubModule_SA_3D__zz_io_MatrixB_7_3[7:0] ), //i
    ._zz_io_A_Valid_0_3 (SubModule_SA_3D__zz_io_A_Valid_0_3      ), //i
    ._zz_io_A_Valid_1_3 (SubModule_SA_3D__zz_io_A_Valid_1_3      ), //i
    ._zz_io_A_Valid_2_3 (SubModule_SA_3D__zz_io_A_Valid_2_3      ), //i
    ._zz_io_A_Valid_3_3 (SubModule_SA_3D__zz_io_A_Valid_3_3      ), //i
    ._zz_io_A_Valid_4_3 (SubModule_SA_3D__zz_io_A_Valid_4_3      ), //i
    ._zz_io_A_Valid_5_3 (SubModule_SA_3D__zz_io_A_Valid_5_3      ), //i
    ._zz_io_A_Valid_6_3 (SubModule_SA_3D__zz_io_A_Valid_6_3      ), //i
    ._zz_io_A_Valid_7_3 (SubModule_SA_3D__zz_io_A_Valid_7_3      ), //i
    ._zz_io_B_Valid_0_3 (SubModule_SA_3D__zz_io_B_Valid_0_3      ), //i
    ._zz_io_B_Valid_1_3 (SubModule_SA_3D__zz_io_B_Valid_1_3      ), //i
    ._zz_io_B_Valid_2_3 (SubModule_SA_3D__zz_io_B_Valid_2_3      ), //i
    ._zz_io_B_Valid_3_3 (SubModule_SA_3D__zz_io_B_Valid_3_3      ), //i
    ._zz_io_B_Valid_4_3 (SubModule_SA_3D__zz_io_B_Valid_4_3      ), //i
    ._zz_io_B_Valid_5_3 (SubModule_SA_3D__zz_io_B_Valid_5_3      ), //i
    ._zz_io_B_Valid_6_3 (SubModule_SA_3D__zz_io_B_Valid_6_3      ), //i
    ._zz_io_B_Valid_7_3 (SubModule_SA_3D__zz_io_B_Valid_7_3      ), //i
    ._zz_io_signCount_3 (SubModule_SA_3D__zz_io_signCount_3[15:0]), //i
    ._zz_io_MatrixA_0_4 (SubModule_SA_3D__zz_io_MatrixA_0_4[7:0] ), //i
    ._zz_io_MatrixA_1_4 (SubModule_SA_3D__zz_io_MatrixA_1_4[7:0] ), //i
    ._zz_io_MatrixA_2_4 (SubModule_SA_3D__zz_io_MatrixA_2_4[7:0] ), //i
    ._zz_io_MatrixA_3_4 (SubModule_SA_3D__zz_io_MatrixA_3_4[7:0] ), //i
    ._zz_io_MatrixA_4_4 (SubModule_SA_3D__zz_io_MatrixA_4_4[7:0] ), //i
    ._zz_io_MatrixA_5_4 (SubModule_SA_3D__zz_io_MatrixA_5_4[7:0] ), //i
    ._zz_io_MatrixA_6_4 (SubModule_SA_3D__zz_io_MatrixA_6_4[7:0] ), //i
    ._zz_io_MatrixA_7_4 (SubModule_SA_3D__zz_io_MatrixA_7_4[7:0] ), //i
    ._zz_io_MatrixB_0_4 (SubModule_SA_3D__zz_io_MatrixB_0_4[7:0] ), //i
    ._zz_io_MatrixB_1_4 (SubModule_SA_3D__zz_io_MatrixB_1_4[7:0] ), //i
    ._zz_io_MatrixB_2_4 (SubModule_SA_3D__zz_io_MatrixB_2_4[7:0] ), //i
    ._zz_io_MatrixB_3_4 (SubModule_SA_3D__zz_io_MatrixB_3_4[7:0] ), //i
    ._zz_io_MatrixB_4_4 (SubModule_SA_3D__zz_io_MatrixB_4_4[7:0] ), //i
    ._zz_io_MatrixB_5_4 (SubModule_SA_3D__zz_io_MatrixB_5_4[7:0] ), //i
    ._zz_io_MatrixB_6_4 (SubModule_SA_3D__zz_io_MatrixB_6_4[7:0] ), //i
    ._zz_io_MatrixB_7_4 (SubModule_SA_3D__zz_io_MatrixB_7_4[7:0] ), //i
    ._zz_io_A_Valid_0_4 (SubModule_SA_3D__zz_io_A_Valid_0_4      ), //i
    ._zz_io_A_Valid_1_4 (SubModule_SA_3D__zz_io_A_Valid_1_4      ), //i
    ._zz_io_A_Valid_2_4 (SubModule_SA_3D__zz_io_A_Valid_2_4      ), //i
    ._zz_io_A_Valid_3_4 (SubModule_SA_3D__zz_io_A_Valid_3_4      ), //i
    ._zz_io_A_Valid_4_4 (SubModule_SA_3D__zz_io_A_Valid_4_4      ), //i
    ._zz_io_A_Valid_5_4 (SubModule_SA_3D__zz_io_A_Valid_5_4      ), //i
    ._zz_io_A_Valid_6_4 (SubModule_SA_3D__zz_io_A_Valid_6_4      ), //i
    ._zz_io_A_Valid_7_4 (SubModule_SA_3D__zz_io_A_Valid_7_4      ), //i
    ._zz_io_B_Valid_0_4 (SubModule_SA_3D__zz_io_B_Valid_0_4      ), //i
    ._zz_io_B_Valid_1_4 (SubModule_SA_3D__zz_io_B_Valid_1_4      ), //i
    ._zz_io_B_Valid_2_4 (SubModule_SA_3D__zz_io_B_Valid_2_4      ), //i
    ._zz_io_B_Valid_3_4 (SubModule_SA_3D__zz_io_B_Valid_3_4      ), //i
    ._zz_io_B_Valid_4_4 (SubModule_SA_3D__zz_io_B_Valid_4_4      ), //i
    ._zz_io_B_Valid_5_4 (SubModule_SA_3D__zz_io_B_Valid_5_4      ), //i
    ._zz_io_B_Valid_6_4 (SubModule_SA_3D__zz_io_B_Valid_6_4      ), //i
    ._zz_io_B_Valid_7_4 (SubModule_SA_3D__zz_io_B_Valid_7_4      ), //i
    ._zz_io_signCount_4 (SubModule_SA_3D__zz_io_signCount_4[15:0]), //i
    ._zz_io_MatrixA_0_5 (SubModule_SA_3D__zz_io_MatrixA_0_5[7:0] ), //i
    ._zz_io_MatrixA_1_5 (SubModule_SA_3D__zz_io_MatrixA_1_5[7:0] ), //i
    ._zz_io_MatrixA_2_5 (SubModule_SA_3D__zz_io_MatrixA_2_5[7:0] ), //i
    ._zz_io_MatrixA_3_5 (SubModule_SA_3D__zz_io_MatrixA_3_5[7:0] ), //i
    ._zz_io_MatrixA_4_5 (SubModule_SA_3D__zz_io_MatrixA_4_5[7:0] ), //i
    ._zz_io_MatrixA_5_5 (SubModule_SA_3D__zz_io_MatrixA_5_5[7:0] ), //i
    ._zz_io_MatrixA_6_5 (SubModule_SA_3D__zz_io_MatrixA_6_5[7:0] ), //i
    ._zz_io_MatrixA_7_5 (SubModule_SA_3D__zz_io_MatrixA_7_5[7:0] ), //i
    ._zz_io_MatrixB_0_5 (SubModule_SA_3D__zz_io_MatrixB_0_5[7:0] ), //i
    ._zz_io_MatrixB_1_5 (SubModule_SA_3D__zz_io_MatrixB_1_5[7:0] ), //i
    ._zz_io_MatrixB_2_5 (SubModule_SA_3D__zz_io_MatrixB_2_5[7:0] ), //i
    ._zz_io_MatrixB_3_5 (SubModule_SA_3D__zz_io_MatrixB_3_5[7:0] ), //i
    ._zz_io_MatrixB_4_5 (SubModule_SA_3D__zz_io_MatrixB_4_5[7:0] ), //i
    ._zz_io_MatrixB_5_5 (SubModule_SA_3D__zz_io_MatrixB_5_5[7:0] ), //i
    ._zz_io_MatrixB_6_5 (SubModule_SA_3D__zz_io_MatrixB_6_5[7:0] ), //i
    ._zz_io_MatrixB_7_5 (SubModule_SA_3D__zz_io_MatrixB_7_5[7:0] ), //i
    ._zz_io_A_Valid_0_5 (SubModule_SA_3D__zz_io_A_Valid_0_5      ), //i
    ._zz_io_A_Valid_1_5 (SubModule_SA_3D__zz_io_A_Valid_1_5      ), //i
    ._zz_io_A_Valid_2_5 (SubModule_SA_3D__zz_io_A_Valid_2_5      ), //i
    ._zz_io_A_Valid_3_5 (SubModule_SA_3D__zz_io_A_Valid_3_5      ), //i
    ._zz_io_A_Valid_4_5 (SubModule_SA_3D__zz_io_A_Valid_4_5      ), //i
    ._zz_io_A_Valid_5_5 (SubModule_SA_3D__zz_io_A_Valid_5_5      ), //i
    ._zz_io_A_Valid_6_5 (SubModule_SA_3D__zz_io_A_Valid_6_5      ), //i
    ._zz_io_A_Valid_7_5 (SubModule_SA_3D__zz_io_A_Valid_7_5      ), //i
    ._zz_io_B_Valid_0_5 (SubModule_SA_3D__zz_io_B_Valid_0_5      ), //i
    ._zz_io_B_Valid_1_5 (SubModule_SA_3D__zz_io_B_Valid_1_5      ), //i
    ._zz_io_B_Valid_2_5 (SubModule_SA_3D__zz_io_B_Valid_2_5      ), //i
    ._zz_io_B_Valid_3_5 (SubModule_SA_3D__zz_io_B_Valid_3_5      ), //i
    ._zz_io_B_Valid_4_5 (SubModule_SA_3D__zz_io_B_Valid_4_5      ), //i
    ._zz_io_B_Valid_5_5 (SubModule_SA_3D__zz_io_B_Valid_5_5      ), //i
    ._zz_io_B_Valid_6_5 (SubModule_SA_3D__zz_io_B_Valid_6_5      ), //i
    ._zz_io_B_Valid_7_5 (SubModule_SA_3D__zz_io_B_Valid_7_5      ), //i
    ._zz_io_signCount_5 (SubModule_SA_3D__zz_io_signCount_5[15:0]), //i
    ._zz_io_MatrixA_0_6 (SubModule_SA_3D__zz_io_MatrixA_0_6[7:0] ), //i
    ._zz_io_MatrixA_1_6 (SubModule_SA_3D__zz_io_MatrixA_1_6[7:0] ), //i
    ._zz_io_MatrixA_2_6 (SubModule_SA_3D__zz_io_MatrixA_2_6[7:0] ), //i
    ._zz_io_MatrixA_3_6 (SubModule_SA_3D__zz_io_MatrixA_3_6[7:0] ), //i
    ._zz_io_MatrixA_4_6 (SubModule_SA_3D__zz_io_MatrixA_4_6[7:0] ), //i
    ._zz_io_MatrixA_5_6 (SubModule_SA_3D__zz_io_MatrixA_5_6[7:0] ), //i
    ._zz_io_MatrixA_6_6 (SubModule_SA_3D__zz_io_MatrixA_6_6[7:0] ), //i
    ._zz_io_MatrixA_7_6 (SubModule_SA_3D__zz_io_MatrixA_7_6[7:0] ), //i
    ._zz_io_MatrixB_0_6 (SubModule_SA_3D__zz_io_MatrixB_0_6[7:0] ), //i
    ._zz_io_MatrixB_1_6 (SubModule_SA_3D__zz_io_MatrixB_1_6[7:0] ), //i
    ._zz_io_MatrixB_2_6 (SubModule_SA_3D__zz_io_MatrixB_2_6[7:0] ), //i
    ._zz_io_MatrixB_3_6 (SubModule_SA_3D__zz_io_MatrixB_3_6[7:0] ), //i
    ._zz_io_MatrixB_4_6 (SubModule_SA_3D__zz_io_MatrixB_4_6[7:0] ), //i
    ._zz_io_MatrixB_5_6 (SubModule_SA_3D__zz_io_MatrixB_5_6[7:0] ), //i
    ._zz_io_MatrixB_6_6 (SubModule_SA_3D__zz_io_MatrixB_6_6[7:0] ), //i
    ._zz_io_MatrixB_7_6 (SubModule_SA_3D__zz_io_MatrixB_7_6[7:0] ), //i
    ._zz_io_A_Valid_0_6 (SubModule_SA_3D__zz_io_A_Valid_0_6      ), //i
    ._zz_io_A_Valid_1_6 (SubModule_SA_3D__zz_io_A_Valid_1_6      ), //i
    ._zz_io_A_Valid_2_6 (SubModule_SA_3D__zz_io_A_Valid_2_6      ), //i
    ._zz_io_A_Valid_3_6 (SubModule_SA_3D__zz_io_A_Valid_3_6      ), //i
    ._zz_io_A_Valid_4_6 (SubModule_SA_3D__zz_io_A_Valid_4_6      ), //i
    ._zz_io_A_Valid_5_6 (SubModule_SA_3D__zz_io_A_Valid_5_6      ), //i
    ._zz_io_A_Valid_6_6 (SubModule_SA_3D__zz_io_A_Valid_6_6      ), //i
    ._zz_io_A_Valid_7_6 (SubModule_SA_3D__zz_io_A_Valid_7_6      ), //i
    ._zz_io_B_Valid_0_6 (SubModule_SA_3D__zz_io_B_Valid_0_6      ), //i
    ._zz_io_B_Valid_1_6 (SubModule_SA_3D__zz_io_B_Valid_1_6      ), //i
    ._zz_io_B_Valid_2_6 (SubModule_SA_3D__zz_io_B_Valid_2_6      ), //i
    ._zz_io_B_Valid_3_6 (SubModule_SA_3D__zz_io_B_Valid_3_6      ), //i
    ._zz_io_B_Valid_4_6 (SubModule_SA_3D__zz_io_B_Valid_4_6      ), //i
    ._zz_io_B_Valid_5_6 (SubModule_SA_3D__zz_io_B_Valid_5_6      ), //i
    ._zz_io_B_Valid_6_6 (SubModule_SA_3D__zz_io_B_Valid_6_6      ), //i
    ._zz_io_B_Valid_7_6 (SubModule_SA_3D__zz_io_B_Valid_7_6      ), //i
    ._zz_io_signCount_6 (SubModule_SA_3D__zz_io_signCount_6[15:0]), //i
    ._zz_io_MatrixA_0_7 (SubModule_SA_3D__zz_io_MatrixA_0_7[7:0] ), //i
    ._zz_io_MatrixA_1_7 (SubModule_SA_3D__zz_io_MatrixA_1_7[7:0] ), //i
    ._zz_io_MatrixA_2_7 (SubModule_SA_3D__zz_io_MatrixA_2_7[7:0] ), //i
    ._zz_io_MatrixA_3_7 (SubModule_SA_3D__zz_io_MatrixA_3_7[7:0] ), //i
    ._zz_io_MatrixA_4_7 (SubModule_SA_3D__zz_io_MatrixA_4_7[7:0] ), //i
    ._zz_io_MatrixA_5_7 (SubModule_SA_3D__zz_io_MatrixA_5_7[7:0] ), //i
    ._zz_io_MatrixA_6_7 (SubModule_SA_3D__zz_io_MatrixA_6_7[7:0] ), //i
    ._zz_io_MatrixA_7_7 (SubModule_SA_3D__zz_io_MatrixA_7_7[7:0] ), //i
    ._zz_io_MatrixB_0_7 (SubModule_SA_3D__zz_io_MatrixB_0_7[7:0] ), //i
    ._zz_io_MatrixB_1_7 (SubModule_SA_3D__zz_io_MatrixB_1_7[7:0] ), //i
    ._zz_io_MatrixB_2_7 (SubModule_SA_3D__zz_io_MatrixB_2_7[7:0] ), //i
    ._zz_io_MatrixB_3_7 (SubModule_SA_3D__zz_io_MatrixB_3_7[7:0] ), //i
    ._zz_io_MatrixB_4_7 (SubModule_SA_3D__zz_io_MatrixB_4_7[7:0] ), //i
    ._zz_io_MatrixB_5_7 (SubModule_SA_3D__zz_io_MatrixB_5_7[7:0] ), //i
    ._zz_io_MatrixB_6_7 (SubModule_SA_3D__zz_io_MatrixB_6_7[7:0] ), //i
    ._zz_io_MatrixB_7_7 (SubModule_SA_3D__zz_io_MatrixB_7_7[7:0] ), //i
    ._zz_io_A_Valid_0_7 (SubModule_SA_3D__zz_io_A_Valid_0_7      ), //i
    ._zz_io_A_Valid_1_7 (SubModule_SA_3D__zz_io_A_Valid_1_7      ), //i
    ._zz_io_A_Valid_2_7 (SubModule_SA_3D__zz_io_A_Valid_2_7      ), //i
    ._zz_io_A_Valid_3_7 (SubModule_SA_3D__zz_io_A_Valid_3_7      ), //i
    ._zz_io_A_Valid_4_7 (SubModule_SA_3D__zz_io_A_Valid_4_7      ), //i
    ._zz_io_A_Valid_5_7 (SubModule_SA_3D__zz_io_A_Valid_5_7      ), //i
    ._zz_io_A_Valid_6_7 (SubModule_SA_3D__zz_io_A_Valid_6_7      ), //i
    ._zz_io_A_Valid_7_7 (SubModule_SA_3D__zz_io_A_Valid_7_7      ), //i
    ._zz_io_B_Valid_0_7 (SubModule_SA_3D__zz_io_B_Valid_0_7      ), //i
    ._zz_io_B_Valid_1_7 (SubModule_SA_3D__zz_io_B_Valid_1_7      ), //i
    ._zz_io_B_Valid_2_7 (SubModule_SA_3D__zz_io_B_Valid_2_7      ), //i
    ._zz_io_B_Valid_3_7 (SubModule_SA_3D__zz_io_B_Valid_3_7      ), //i
    ._zz_io_B_Valid_4_7 (SubModule_SA_3D__zz_io_B_Valid_4_7      ), //i
    ._zz_io_B_Valid_5_7 (SubModule_SA_3D__zz_io_B_Valid_5_7      ), //i
    ._zz_io_B_Valid_6_7 (SubModule_SA_3D__zz_io_B_Valid_6_7      ), //i
    ._zz_io_B_Valid_7_7 (SubModule_SA_3D__zz_io_B_Valid_7_7      ), //i
    ._zz_io_signCount_7 (SubModule_SA_3D__zz_io_signCount_7[15:0]), //i
    .reset              (reset                                   )  //i
  );
  WeightCache_Stream SubModule_WeightCache (
    .s_axis_s2mm_tdata  (InputSwitch_m_0_axis_mm2s_tdata[63:0]       ), //i
    .s_axis_s2mm_tkeep  (InputSwitch_m_0_axis_mm2s_tkeep[7:0]        ), //i
    .s_axis_s2mm_tlast  (InputSwitch_m_0_axis_mm2s_tlast             ), //i
    .s_axis_s2mm_tready (SubModule_WeightCache_s_axis_s2mm_tready    ), //o
    .s_axis_s2mm_tvalid (InputSwitch_m_0_axis_mm2s_tvalid            ), //i
    .start              (_zz_start_2                                 ), //i
    .Matrix_Row         (Img2Col_WeightMatrix_Row[15:0]              ), //i
    .Matrix_Col         (Img2Col_OutFeature_Channel[15:0]            ), //i
    .mData_0            (SubModule_WeightCache_mData_0[7:0]          ), //o
    .mData_1            (SubModule_WeightCache_mData_1[7:0]          ), //o
    .mData_2            (SubModule_WeightCache_mData_2[7:0]          ), //o
    .mData_3            (SubModule_WeightCache_mData_3[7:0]          ), //o
    .mData_4            (SubModule_WeightCache_mData_4[7:0]          ), //o
    .mData_5            (SubModule_WeightCache_mData_5[7:0]          ), //o
    .mData_6            (SubModule_WeightCache_mData_6[7:0]          ), //o
    .mData_7            (SubModule_WeightCache_mData_7[7:0]          ), //o
    .mData_8            (SubModule_WeightCache_mData_8[7:0]          ), //o
    .mData_9            (SubModule_WeightCache_mData_9[7:0]          ), //o
    .mData_10           (SubModule_WeightCache_mData_10[7:0]         ), //o
    .mData_11           (SubModule_WeightCache_mData_11[7:0]         ), //o
    .mData_12           (SubModule_WeightCache_mData_12[7:0]         ), //o
    .mData_13           (SubModule_WeightCache_mData_13[7:0]         ), //o
    .mData_14           (SubModule_WeightCache_mData_14[7:0]         ), //o
    .mData_15           (SubModule_WeightCache_mData_15[7:0]         ), //o
    .mData_16           (SubModule_WeightCache_mData_16[7:0]         ), //o
    .mData_17           (SubModule_WeightCache_mData_17[7:0]         ), //o
    .mData_18           (SubModule_WeightCache_mData_18[7:0]         ), //o
    .mData_19           (SubModule_WeightCache_mData_19[7:0]         ), //o
    .mData_20           (SubModule_WeightCache_mData_20[7:0]         ), //o
    .mData_21           (SubModule_WeightCache_mData_21[7:0]         ), //o
    .mData_22           (SubModule_WeightCache_mData_22[7:0]         ), //o
    .mData_23           (SubModule_WeightCache_mData_23[7:0]         ), //o
    .mData_24           (SubModule_WeightCache_mData_24[7:0]         ), //o
    .mData_25           (SubModule_WeightCache_mData_25[7:0]         ), //o
    .mData_26           (SubModule_WeightCache_mData_26[7:0]         ), //o
    .mData_27           (SubModule_WeightCache_mData_27[7:0]         ), //o
    .mData_28           (SubModule_WeightCache_mData_28[7:0]         ), //o
    .mData_29           (SubModule_WeightCache_mData_29[7:0]         ), //o
    .mData_30           (SubModule_WeightCache_mData_30[7:0]         ), //o
    .mData_31           (SubModule_WeightCache_mData_31[7:0]         ), //o
    .mData_32           (SubModule_WeightCache_mData_32[7:0]         ), //o
    .mData_33           (SubModule_WeightCache_mData_33[7:0]         ), //o
    .mData_34           (SubModule_WeightCache_mData_34[7:0]         ), //o
    .mData_35           (SubModule_WeightCache_mData_35[7:0]         ), //o
    .mData_36           (SubModule_WeightCache_mData_36[7:0]         ), //o
    .mData_37           (SubModule_WeightCache_mData_37[7:0]         ), //o
    .mData_38           (SubModule_WeightCache_mData_38[7:0]         ), //o
    .mData_39           (SubModule_WeightCache_mData_39[7:0]         ), //o
    .mData_40           (SubModule_WeightCache_mData_40[7:0]         ), //o
    .mData_41           (SubModule_WeightCache_mData_41[7:0]         ), //o
    .mData_42           (SubModule_WeightCache_mData_42[7:0]         ), //o
    .mData_43           (SubModule_WeightCache_mData_43[7:0]         ), //o
    .mData_44           (SubModule_WeightCache_mData_44[7:0]         ), //o
    .mData_45           (SubModule_WeightCache_mData_45[7:0]         ), //o
    .mData_46           (SubModule_WeightCache_mData_46[7:0]         ), //o
    .mData_47           (SubModule_WeightCache_mData_47[7:0]         ), //o
    .mData_48           (SubModule_WeightCache_mData_48[7:0]         ), //o
    .mData_49           (SubModule_WeightCache_mData_49[7:0]         ), //o
    .mData_50           (SubModule_WeightCache_mData_50[7:0]         ), //o
    .mData_51           (SubModule_WeightCache_mData_51[7:0]         ), //o
    .mData_52           (SubModule_WeightCache_mData_52[7:0]         ), //o
    .mData_53           (SubModule_WeightCache_mData_53[7:0]         ), //o
    .mData_54           (SubModule_WeightCache_mData_54[7:0]         ), //o
    .mData_55           (SubModule_WeightCache_mData_55[7:0]         ), //o
    .mData_56           (SubModule_WeightCache_mData_56[7:0]         ), //o
    .mData_57           (SubModule_WeightCache_mData_57[7:0]         ), //o
    .mData_58           (SubModule_WeightCache_mData_58[7:0]         ), //o
    .mData_59           (SubModule_WeightCache_mData_59[7:0]         ), //o
    .mData_60           (SubModule_WeightCache_mData_60[7:0]         ), //o
    .mData_61           (SubModule_WeightCache_mData_61[7:0]         ), //o
    .mData_62           (SubModule_WeightCache_mData_62[7:0]         ), //o
    .mData_63           (SubModule_WeightCache_mData_63[7:0]         ), //o
    .Raddr_Valid        (SubModule_Img2Col_Raddr_Valid               ), //i
    .Weight_Cached      (SubModule_WeightCache_Weight_Cached         ), //o
    .LayerEnd           (LayerEnd                                    ), //i
    .MatrixCol_Switch   (SubModule_WeightCache_MatrixCol_Switch[63:0]), //o
    .clk                (clk                                         ), //i
    .reset              (reset                                       )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      TopCtrl_Enum_IDLE : Fsm_currentState_string = "IDLE            ";
      TopCtrl_Enum_INIT : Fsm_currentState_string = "INIT            ";
      TopCtrl_Enum_WEIGHT_CACHE : Fsm_currentState_string = "WEIGHT_CACHE    ";
      TopCtrl_Enum_RECEIVE_PICTURE : Fsm_currentState_string = "RECEIVE_PICTURE ";
      TopCtrl_Enum_RECEIVE_MATRIX : Fsm_currentState_string = "RECEIVE_MATRIX  ";
      TopCtrl_Enum_WAIT_COMPUTE_END : Fsm_currentState_string = "WAIT_COMPUTE_END";
      default : Fsm_currentState_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      TopCtrl_Enum_IDLE : Fsm_nextState_string = "IDLE            ";
      TopCtrl_Enum_INIT : Fsm_nextState_string = "INIT            ";
      TopCtrl_Enum_WEIGHT_CACHE : Fsm_nextState_string = "WEIGHT_CACHE    ";
      TopCtrl_Enum_RECEIVE_PICTURE : Fsm_nextState_string = "RECEIVE_PICTURE ";
      TopCtrl_Enum_RECEIVE_MATRIX : Fsm_nextState_string = "RECEIVE_MATRIX  ";
      TopCtrl_Enum_WAIT_COMPUTE_END : Fsm_nextState_string = "WAIT_COMPUTE_END";
      default : Fsm_nextState_string = "????????????????";
    endcase
  end
  `endif

  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & TopCtrl_Enum_IDLE) == TopCtrl_Enum_IDLE) : begin
        if(Control_start) begin
          Fsm_nextState = TopCtrl_Enum_INIT;
        end else begin
          Fsm_nextState = TopCtrl_Enum_IDLE;
        end
      end
      (((Fsm_currentState) & TopCtrl_Enum_INIT) == TopCtrl_Enum_INIT) : begin
        if(Fsm_Inited) begin
          Fsm_nextState = TopCtrl_Enum_WEIGHT_CACHE;
        end else begin
          Fsm_nextState = TopCtrl_Enum_INIT;
        end
      end
      (((Fsm_currentState) & TopCtrl_Enum_WEIGHT_CACHE) == TopCtrl_Enum_WEIGHT_CACHE) : begin
        if(when_SA3D_Top_l46) begin
          Fsm_nextState = TopCtrl_Enum_RECEIVE_PICTURE;
        end else begin
          if(when_SA3D_Top_l48) begin
            Fsm_nextState = TopCtrl_Enum_RECEIVE_MATRIX;
          end else begin
            Fsm_nextState = TopCtrl_Enum_WEIGHT_CACHE;
          end
        end
      end
      (((Fsm_currentState) & TopCtrl_Enum_RECEIVE_PICTURE) == TopCtrl_Enum_RECEIVE_PICTURE) : begin
        if(Fsm_Picture_Received) begin
          Fsm_nextState = TopCtrl_Enum_WAIT_COMPUTE_END;
        end else begin
          Fsm_nextState = TopCtrl_Enum_RECEIVE_PICTURE;
        end
      end
      (((Fsm_currentState) & TopCtrl_Enum_RECEIVE_MATRIX) == TopCtrl_Enum_RECEIVE_MATRIX) : begin
        if(Fsm_Matrix_Received) begin
          Fsm_nextState = TopCtrl_Enum_WAIT_COMPUTE_END;
        end else begin
          Fsm_nextState = TopCtrl_Enum_RECEIVE_MATRIX;
        end
      end
      default : begin
        if(Fsm_Compute_End) begin
          Fsm_nextState = TopCtrl_Enum_IDLE;
        end else begin
          Fsm_nextState = TopCtrl_Enum_WAIT_COMPUTE_END;
        end
      end
    endcase
  end

  assign when_SA3D_Top_l46 = (Fsm_WeightCached && Fsm_Switch_Conv);
  assign when_SA3D_Top_l48 = (Fsm_WeightCached && (! Fsm_Switch_Conv));
  assign Fsm_Compute_End = LayerEnd;
  assign when_WaCounter_l19 = ((Fsm_currentState & TopCtrl_Enum_INIT) != 6'b000000);
  assign when_WaCounter_l14 = (InitCnt_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l14) begin
      InitCnt_valid = 1'b1;
    end else begin
      InitCnt_valid = 1'b0;
    end
  end

  assign Fsm_Inited = InitCnt_valid;
  assign s_axis_s2mm_tready = InputSwitch_s0_axis_s2mm_tready;
  assign when_SA3D_Top_l131 = ((Fsm_currentState & TopCtrl_Enum_WEIGHT_CACHE) != 6'b000000);
  always @(*) begin
    if(when_SA3D_Top_l131) begin
      InputSwitch_Switch = 2'b00;
    end else begin
      if(Control_Switch_Conv) begin
        InputSwitch_Switch = 2'b01;
      end else begin
        InputSwitch_Switch = 2'b10;
      end
    end
  end

  assign SubModule_SA_3D__zz_io_signCount = (Img2Col_WeightMatrix_Row - 16'h0001);
  assign SubModule_SA_3D__zz_io_MatrixA_0 = SubModule_Img2Col_mData[7 : 0];
  assign SubModule_SA_3D__zz_io_A_Valid_0 = SubModule_Img2Col_mValid[0];
  assign SubModule_SA_3D__zz_io_MatrixA_1 = SubModule_Img2Col_mData[7 : 0];
  assign SubModule_SA_3D__zz_io_A_Valid_1 = SubModule_Img2Col_mValid[0];
  assign SubModule_SA_3D__zz_io_MatrixA_2 = SubModule_Img2Col_mData[7 : 0];
  assign SubModule_SA_3D__zz_io_A_Valid_2 = SubModule_Img2Col_mValid[0];
  assign SubModule_SA_3D__zz_io_MatrixA_3 = SubModule_Img2Col_mData[7 : 0];
  assign SubModule_SA_3D__zz_io_A_Valid_3 = SubModule_Img2Col_mValid[0];
  assign SubModule_SA_3D__zz_io_MatrixA_4 = SubModule_Img2Col_mData[7 : 0];
  assign SubModule_SA_3D__zz_io_A_Valid_4 = SubModule_Img2Col_mValid[0];
  assign SubModule_SA_3D__zz_io_MatrixA_5 = SubModule_Img2Col_mData[7 : 0];
  assign SubModule_SA_3D__zz_io_A_Valid_5 = SubModule_Img2Col_mValid[0];
  assign SubModule_SA_3D__zz_io_MatrixA_6 = SubModule_Img2Col_mData[7 : 0];
  assign SubModule_SA_3D__zz_io_A_Valid_6 = SubModule_Img2Col_mValid[0];
  assign SubModule_SA_3D__zz_io_MatrixA_7 = SubModule_Img2Col_mData[7 : 0];
  assign SubModule_SA_3D__zz_io_A_Valid_7 = SubModule_Img2Col_mValid[0];
  assign SubModule_SA_3D__zz_io_signCount_1 = (Img2Col_WeightMatrix_Row - 16'h0001);
  assign SubModule_SA_3D__zz_io_MatrixA_0_1 = SubModule_Img2Col_mData[15 : 8];
  assign SubModule_SA_3D__zz_io_A_Valid_0_1 = SubModule_Img2Col_mValid[1];
  assign SubModule_SA_3D__zz_io_MatrixA_1_1 = SubModule_Img2Col_mData[15 : 8];
  assign SubModule_SA_3D__zz_io_A_Valid_1_1 = SubModule_Img2Col_mValid[1];
  assign SubModule_SA_3D__zz_io_MatrixA_2_1 = SubModule_Img2Col_mData[15 : 8];
  assign SubModule_SA_3D__zz_io_A_Valid_2_1 = SubModule_Img2Col_mValid[1];
  assign SubModule_SA_3D__zz_io_MatrixA_3_1 = SubModule_Img2Col_mData[15 : 8];
  assign SubModule_SA_3D__zz_io_A_Valid_3_1 = SubModule_Img2Col_mValid[1];
  assign SubModule_SA_3D__zz_io_MatrixA_4_1 = SubModule_Img2Col_mData[15 : 8];
  assign SubModule_SA_3D__zz_io_A_Valid_4_1 = SubModule_Img2Col_mValid[1];
  assign SubModule_SA_3D__zz_io_MatrixA_5_1 = SubModule_Img2Col_mData[15 : 8];
  assign SubModule_SA_3D__zz_io_A_Valid_5_1 = SubModule_Img2Col_mValid[1];
  assign SubModule_SA_3D__zz_io_MatrixA_6_1 = SubModule_Img2Col_mData[15 : 8];
  assign SubModule_SA_3D__zz_io_A_Valid_6_1 = SubModule_Img2Col_mValid[1];
  assign SubModule_SA_3D__zz_io_MatrixA_7_1 = SubModule_Img2Col_mData[15 : 8];
  assign SubModule_SA_3D__zz_io_A_Valid_7_1 = SubModule_Img2Col_mValid[1];
  assign SubModule_SA_3D__zz_io_signCount_2 = (Img2Col_WeightMatrix_Row - 16'h0001);
  assign SubModule_SA_3D__zz_io_MatrixA_0_2 = SubModule_Img2Col_mData[23 : 16];
  assign SubModule_SA_3D__zz_io_A_Valid_0_2 = SubModule_Img2Col_mValid[2];
  assign SubModule_SA_3D__zz_io_MatrixA_1_2 = SubModule_Img2Col_mData[23 : 16];
  assign SubModule_SA_3D__zz_io_A_Valid_1_2 = SubModule_Img2Col_mValid[2];
  assign SubModule_SA_3D__zz_io_MatrixA_2_2 = SubModule_Img2Col_mData[23 : 16];
  assign SubModule_SA_3D__zz_io_A_Valid_2_2 = SubModule_Img2Col_mValid[2];
  assign SubModule_SA_3D__zz_io_MatrixA_3_2 = SubModule_Img2Col_mData[23 : 16];
  assign SubModule_SA_3D__zz_io_A_Valid_3_2 = SubModule_Img2Col_mValid[2];
  assign SubModule_SA_3D__zz_io_MatrixA_4_2 = SubModule_Img2Col_mData[23 : 16];
  assign SubModule_SA_3D__zz_io_A_Valid_4_2 = SubModule_Img2Col_mValid[2];
  assign SubModule_SA_3D__zz_io_MatrixA_5_2 = SubModule_Img2Col_mData[23 : 16];
  assign SubModule_SA_3D__zz_io_A_Valid_5_2 = SubModule_Img2Col_mValid[2];
  assign SubModule_SA_3D__zz_io_MatrixA_6_2 = SubModule_Img2Col_mData[23 : 16];
  assign SubModule_SA_3D__zz_io_A_Valid_6_2 = SubModule_Img2Col_mValid[2];
  assign SubModule_SA_3D__zz_io_MatrixA_7_2 = SubModule_Img2Col_mData[23 : 16];
  assign SubModule_SA_3D__zz_io_A_Valid_7_2 = SubModule_Img2Col_mValid[2];
  assign SubModule_SA_3D__zz_io_signCount_3 = (Img2Col_WeightMatrix_Row - 16'h0001);
  assign SubModule_SA_3D__zz_io_MatrixA_0_3 = SubModule_Img2Col_mData[31 : 24];
  assign SubModule_SA_3D__zz_io_A_Valid_0_3 = SubModule_Img2Col_mValid[3];
  assign SubModule_SA_3D__zz_io_MatrixA_1_3 = SubModule_Img2Col_mData[31 : 24];
  assign SubModule_SA_3D__zz_io_A_Valid_1_3 = SubModule_Img2Col_mValid[3];
  assign SubModule_SA_3D__zz_io_MatrixA_2_3 = SubModule_Img2Col_mData[31 : 24];
  assign SubModule_SA_3D__zz_io_A_Valid_2_3 = SubModule_Img2Col_mValid[3];
  assign SubModule_SA_3D__zz_io_MatrixA_3_3 = SubModule_Img2Col_mData[31 : 24];
  assign SubModule_SA_3D__zz_io_A_Valid_3_3 = SubModule_Img2Col_mValid[3];
  assign SubModule_SA_3D__zz_io_MatrixA_4_3 = SubModule_Img2Col_mData[31 : 24];
  assign SubModule_SA_3D__zz_io_A_Valid_4_3 = SubModule_Img2Col_mValid[3];
  assign SubModule_SA_3D__zz_io_MatrixA_5_3 = SubModule_Img2Col_mData[31 : 24];
  assign SubModule_SA_3D__zz_io_A_Valid_5_3 = SubModule_Img2Col_mValid[3];
  assign SubModule_SA_3D__zz_io_MatrixA_6_3 = SubModule_Img2Col_mData[31 : 24];
  assign SubModule_SA_3D__zz_io_A_Valid_6_3 = SubModule_Img2Col_mValid[3];
  assign SubModule_SA_3D__zz_io_MatrixA_7_3 = SubModule_Img2Col_mData[31 : 24];
  assign SubModule_SA_3D__zz_io_A_Valid_7_3 = SubModule_Img2Col_mValid[3];
  assign SubModule_SA_3D__zz_io_signCount_4 = (Img2Col_WeightMatrix_Row - 16'h0001);
  assign SubModule_SA_3D__zz_io_MatrixA_0_4 = SubModule_Img2Col_mData[39 : 32];
  assign SubModule_SA_3D__zz_io_A_Valid_0_4 = SubModule_Img2Col_mValid[4];
  assign SubModule_SA_3D__zz_io_MatrixA_1_4 = SubModule_Img2Col_mData[39 : 32];
  assign SubModule_SA_3D__zz_io_A_Valid_1_4 = SubModule_Img2Col_mValid[4];
  assign SubModule_SA_3D__zz_io_MatrixA_2_4 = SubModule_Img2Col_mData[39 : 32];
  assign SubModule_SA_3D__zz_io_A_Valid_2_4 = SubModule_Img2Col_mValid[4];
  assign SubModule_SA_3D__zz_io_MatrixA_3_4 = SubModule_Img2Col_mData[39 : 32];
  assign SubModule_SA_3D__zz_io_A_Valid_3_4 = SubModule_Img2Col_mValid[4];
  assign SubModule_SA_3D__zz_io_MatrixA_4_4 = SubModule_Img2Col_mData[39 : 32];
  assign SubModule_SA_3D__zz_io_A_Valid_4_4 = SubModule_Img2Col_mValid[4];
  assign SubModule_SA_3D__zz_io_MatrixA_5_4 = SubModule_Img2Col_mData[39 : 32];
  assign SubModule_SA_3D__zz_io_A_Valid_5_4 = SubModule_Img2Col_mValid[4];
  assign SubModule_SA_3D__zz_io_MatrixA_6_4 = SubModule_Img2Col_mData[39 : 32];
  assign SubModule_SA_3D__zz_io_A_Valid_6_4 = SubModule_Img2Col_mValid[4];
  assign SubModule_SA_3D__zz_io_MatrixA_7_4 = SubModule_Img2Col_mData[39 : 32];
  assign SubModule_SA_3D__zz_io_A_Valid_7_4 = SubModule_Img2Col_mValid[4];
  assign SubModule_SA_3D__zz_io_signCount_5 = (Img2Col_WeightMatrix_Row - 16'h0001);
  assign SubModule_SA_3D__zz_io_MatrixA_0_5 = SubModule_Img2Col_mData[47 : 40];
  assign SubModule_SA_3D__zz_io_A_Valid_0_5 = SubModule_Img2Col_mValid[5];
  assign SubModule_SA_3D__zz_io_MatrixA_1_5 = SubModule_Img2Col_mData[47 : 40];
  assign SubModule_SA_3D__zz_io_A_Valid_1_5 = SubModule_Img2Col_mValid[5];
  assign SubModule_SA_3D__zz_io_MatrixA_2_5 = SubModule_Img2Col_mData[47 : 40];
  assign SubModule_SA_3D__zz_io_A_Valid_2_5 = SubModule_Img2Col_mValid[5];
  assign SubModule_SA_3D__zz_io_MatrixA_3_5 = SubModule_Img2Col_mData[47 : 40];
  assign SubModule_SA_3D__zz_io_A_Valid_3_5 = SubModule_Img2Col_mValid[5];
  assign SubModule_SA_3D__zz_io_MatrixA_4_5 = SubModule_Img2Col_mData[47 : 40];
  assign SubModule_SA_3D__zz_io_A_Valid_4_5 = SubModule_Img2Col_mValid[5];
  assign SubModule_SA_3D__zz_io_MatrixA_5_5 = SubModule_Img2Col_mData[47 : 40];
  assign SubModule_SA_3D__zz_io_A_Valid_5_5 = SubModule_Img2Col_mValid[5];
  assign SubModule_SA_3D__zz_io_MatrixA_6_5 = SubModule_Img2Col_mData[47 : 40];
  assign SubModule_SA_3D__zz_io_A_Valid_6_5 = SubModule_Img2Col_mValid[5];
  assign SubModule_SA_3D__zz_io_MatrixA_7_5 = SubModule_Img2Col_mData[47 : 40];
  assign SubModule_SA_3D__zz_io_A_Valid_7_5 = SubModule_Img2Col_mValid[5];
  assign SubModule_SA_3D__zz_io_signCount_6 = (Img2Col_WeightMatrix_Row - 16'h0001);
  assign SubModule_SA_3D__zz_io_MatrixA_0_6 = SubModule_Img2Col_mData[55 : 48];
  assign SubModule_SA_3D__zz_io_A_Valid_0_6 = SubModule_Img2Col_mValid[6];
  assign SubModule_SA_3D__zz_io_MatrixA_1_6 = SubModule_Img2Col_mData[55 : 48];
  assign SubModule_SA_3D__zz_io_A_Valid_1_6 = SubModule_Img2Col_mValid[6];
  assign SubModule_SA_3D__zz_io_MatrixA_2_6 = SubModule_Img2Col_mData[55 : 48];
  assign SubModule_SA_3D__zz_io_A_Valid_2_6 = SubModule_Img2Col_mValid[6];
  assign SubModule_SA_3D__zz_io_MatrixA_3_6 = SubModule_Img2Col_mData[55 : 48];
  assign SubModule_SA_3D__zz_io_A_Valid_3_6 = SubModule_Img2Col_mValid[6];
  assign SubModule_SA_3D__zz_io_MatrixA_4_6 = SubModule_Img2Col_mData[55 : 48];
  assign SubModule_SA_3D__zz_io_A_Valid_4_6 = SubModule_Img2Col_mValid[6];
  assign SubModule_SA_3D__zz_io_MatrixA_5_6 = SubModule_Img2Col_mData[55 : 48];
  assign SubModule_SA_3D__zz_io_A_Valid_5_6 = SubModule_Img2Col_mValid[6];
  assign SubModule_SA_3D__zz_io_MatrixA_6_6 = SubModule_Img2Col_mData[55 : 48];
  assign SubModule_SA_3D__zz_io_A_Valid_6_6 = SubModule_Img2Col_mValid[6];
  assign SubModule_SA_3D__zz_io_MatrixA_7_6 = SubModule_Img2Col_mData[55 : 48];
  assign SubModule_SA_3D__zz_io_A_Valid_7_6 = SubModule_Img2Col_mValid[6];
  assign SubModule_SA_3D__zz_io_signCount_7 = (Img2Col_WeightMatrix_Row - 16'h0001);
  assign SubModule_SA_3D__zz_io_MatrixA_0_7 = SubModule_Img2Col_mData[63 : 56];
  assign SubModule_SA_3D__zz_io_A_Valid_0_7 = SubModule_Img2Col_mValid[7];
  assign SubModule_SA_3D__zz_io_MatrixA_1_7 = SubModule_Img2Col_mData[63 : 56];
  assign SubModule_SA_3D__zz_io_A_Valid_1_7 = SubModule_Img2Col_mValid[7];
  assign SubModule_SA_3D__zz_io_MatrixA_2_7 = SubModule_Img2Col_mData[63 : 56];
  assign SubModule_SA_3D__zz_io_A_Valid_2_7 = SubModule_Img2Col_mValid[7];
  assign SubModule_SA_3D__zz_io_MatrixA_3_7 = SubModule_Img2Col_mData[63 : 56];
  assign SubModule_SA_3D__zz_io_A_Valid_3_7 = SubModule_Img2Col_mValid[7];
  assign SubModule_SA_3D__zz_io_MatrixA_4_7 = SubModule_Img2Col_mData[63 : 56];
  assign SubModule_SA_3D__zz_io_A_Valid_4_7 = SubModule_Img2Col_mValid[7];
  assign SubModule_SA_3D__zz_io_MatrixA_5_7 = SubModule_Img2Col_mData[63 : 56];
  assign SubModule_SA_3D__zz_io_A_Valid_5_7 = SubModule_Img2Col_mValid[7];
  assign SubModule_SA_3D__zz_io_MatrixA_6_7 = SubModule_Img2Col_mData[63 : 56];
  assign SubModule_SA_3D__zz_io_A_Valid_6_7 = SubModule_Img2Col_mValid[7];
  assign SubModule_SA_3D__zz_io_MatrixA_7_7 = SubModule_Img2Col_mData[63 : 56];
  assign SubModule_SA_3D__zz_io_A_Valid_7_7 = SubModule_Img2Col_mValid[7];
  assign SubModule_SA_3D__zz_io_MatrixB_0 = SubModule_WeightCache_mData_0;
  assign SubModule_SA_3D__zz_io_B_Valid_0 = SubModule_WeightCache_MatrixCol_Switch[0];
  assign SubModule_SA_3D__zz_io_MatrixB_0_1 = SubModule_WeightCache_mData_1;
  assign SubModule_SA_3D__zz_io_B_Valid_0_1 = SubModule_WeightCache_MatrixCol_Switch[1];
  assign SubModule_SA_3D__zz_io_MatrixB_0_2 = SubModule_WeightCache_mData_2;
  assign SubModule_SA_3D__zz_io_B_Valid_0_2 = SubModule_WeightCache_MatrixCol_Switch[2];
  assign SubModule_SA_3D__zz_io_MatrixB_0_3 = SubModule_WeightCache_mData_3;
  assign SubModule_SA_3D__zz_io_B_Valid_0_3 = SubModule_WeightCache_MatrixCol_Switch[3];
  assign SubModule_SA_3D__zz_io_MatrixB_0_4 = SubModule_WeightCache_mData_4;
  assign SubModule_SA_3D__zz_io_B_Valid_0_4 = SubModule_WeightCache_MatrixCol_Switch[4];
  assign SubModule_SA_3D__zz_io_MatrixB_0_5 = SubModule_WeightCache_mData_5;
  assign SubModule_SA_3D__zz_io_B_Valid_0_5 = SubModule_WeightCache_MatrixCol_Switch[5];
  assign SubModule_SA_3D__zz_io_MatrixB_0_6 = SubModule_WeightCache_mData_6;
  assign SubModule_SA_3D__zz_io_B_Valid_0_6 = SubModule_WeightCache_MatrixCol_Switch[6];
  assign SubModule_SA_3D__zz_io_MatrixB_0_7 = SubModule_WeightCache_mData_7;
  assign SubModule_SA_3D__zz_io_B_Valid_0_7 = SubModule_WeightCache_MatrixCol_Switch[7];
  assign SubModule_SA_3D__zz_io_MatrixB_1 = SubModule_WeightCache_mData_8;
  assign SubModule_SA_3D__zz_io_B_Valid_1 = SubModule_WeightCache_MatrixCol_Switch[8];
  assign SubModule_SA_3D__zz_io_MatrixB_1_1 = SubModule_WeightCache_mData_9;
  assign SubModule_SA_3D__zz_io_B_Valid_1_1 = SubModule_WeightCache_MatrixCol_Switch[9];
  assign SubModule_SA_3D__zz_io_MatrixB_1_2 = SubModule_WeightCache_mData_10;
  assign SubModule_SA_3D__zz_io_B_Valid_1_2 = SubModule_WeightCache_MatrixCol_Switch[10];
  assign SubModule_SA_3D__zz_io_MatrixB_1_3 = SubModule_WeightCache_mData_11;
  assign SubModule_SA_3D__zz_io_B_Valid_1_3 = SubModule_WeightCache_MatrixCol_Switch[11];
  assign SubModule_SA_3D__zz_io_MatrixB_1_4 = SubModule_WeightCache_mData_12;
  assign SubModule_SA_3D__zz_io_B_Valid_1_4 = SubModule_WeightCache_MatrixCol_Switch[12];
  assign SubModule_SA_3D__zz_io_MatrixB_1_5 = SubModule_WeightCache_mData_13;
  assign SubModule_SA_3D__zz_io_B_Valid_1_5 = SubModule_WeightCache_MatrixCol_Switch[13];
  assign SubModule_SA_3D__zz_io_MatrixB_1_6 = SubModule_WeightCache_mData_14;
  assign SubModule_SA_3D__zz_io_B_Valid_1_6 = SubModule_WeightCache_MatrixCol_Switch[14];
  assign SubModule_SA_3D__zz_io_MatrixB_1_7 = SubModule_WeightCache_mData_15;
  assign SubModule_SA_3D__zz_io_B_Valid_1_7 = SubModule_WeightCache_MatrixCol_Switch[15];
  assign SubModule_SA_3D__zz_io_MatrixB_2 = SubModule_WeightCache_mData_16;
  assign SubModule_SA_3D__zz_io_B_Valid_2 = SubModule_WeightCache_MatrixCol_Switch[16];
  assign SubModule_SA_3D__zz_io_MatrixB_2_1 = SubModule_WeightCache_mData_17;
  assign SubModule_SA_3D__zz_io_B_Valid_2_1 = SubModule_WeightCache_MatrixCol_Switch[17];
  assign SubModule_SA_3D__zz_io_MatrixB_2_2 = SubModule_WeightCache_mData_18;
  assign SubModule_SA_3D__zz_io_B_Valid_2_2 = SubModule_WeightCache_MatrixCol_Switch[18];
  assign SubModule_SA_3D__zz_io_MatrixB_2_3 = SubModule_WeightCache_mData_19;
  assign SubModule_SA_3D__zz_io_B_Valid_2_3 = SubModule_WeightCache_MatrixCol_Switch[19];
  assign SubModule_SA_3D__zz_io_MatrixB_2_4 = SubModule_WeightCache_mData_20;
  assign SubModule_SA_3D__zz_io_B_Valid_2_4 = SubModule_WeightCache_MatrixCol_Switch[20];
  assign SubModule_SA_3D__zz_io_MatrixB_2_5 = SubModule_WeightCache_mData_21;
  assign SubModule_SA_3D__zz_io_B_Valid_2_5 = SubModule_WeightCache_MatrixCol_Switch[21];
  assign SubModule_SA_3D__zz_io_MatrixB_2_6 = SubModule_WeightCache_mData_22;
  assign SubModule_SA_3D__zz_io_B_Valid_2_6 = SubModule_WeightCache_MatrixCol_Switch[22];
  assign SubModule_SA_3D__zz_io_MatrixB_2_7 = SubModule_WeightCache_mData_23;
  assign SubModule_SA_3D__zz_io_B_Valid_2_7 = SubModule_WeightCache_MatrixCol_Switch[23];
  assign SubModule_SA_3D__zz_io_MatrixB_3 = SubModule_WeightCache_mData_24;
  assign SubModule_SA_3D__zz_io_B_Valid_3 = SubModule_WeightCache_MatrixCol_Switch[24];
  assign SubModule_SA_3D__zz_io_MatrixB_3_1 = SubModule_WeightCache_mData_25;
  assign SubModule_SA_3D__zz_io_B_Valid_3_1 = SubModule_WeightCache_MatrixCol_Switch[25];
  assign SubModule_SA_3D__zz_io_MatrixB_3_2 = SubModule_WeightCache_mData_26;
  assign SubModule_SA_3D__zz_io_B_Valid_3_2 = SubModule_WeightCache_MatrixCol_Switch[26];
  assign SubModule_SA_3D__zz_io_MatrixB_3_3 = SubModule_WeightCache_mData_27;
  assign SubModule_SA_3D__zz_io_B_Valid_3_3 = SubModule_WeightCache_MatrixCol_Switch[27];
  assign SubModule_SA_3D__zz_io_MatrixB_3_4 = SubModule_WeightCache_mData_28;
  assign SubModule_SA_3D__zz_io_B_Valid_3_4 = SubModule_WeightCache_MatrixCol_Switch[28];
  assign SubModule_SA_3D__zz_io_MatrixB_3_5 = SubModule_WeightCache_mData_29;
  assign SubModule_SA_3D__zz_io_B_Valid_3_5 = SubModule_WeightCache_MatrixCol_Switch[29];
  assign SubModule_SA_3D__zz_io_MatrixB_3_6 = SubModule_WeightCache_mData_30;
  assign SubModule_SA_3D__zz_io_B_Valid_3_6 = SubModule_WeightCache_MatrixCol_Switch[30];
  assign SubModule_SA_3D__zz_io_MatrixB_3_7 = SubModule_WeightCache_mData_31;
  assign SubModule_SA_3D__zz_io_B_Valid_3_7 = SubModule_WeightCache_MatrixCol_Switch[31];
  assign SubModule_SA_3D__zz_io_MatrixB_4 = SubModule_WeightCache_mData_32;
  assign SubModule_SA_3D__zz_io_B_Valid_4 = SubModule_WeightCache_MatrixCol_Switch[32];
  assign SubModule_SA_3D__zz_io_MatrixB_4_1 = SubModule_WeightCache_mData_33;
  assign SubModule_SA_3D__zz_io_B_Valid_4_1 = SubModule_WeightCache_MatrixCol_Switch[33];
  assign SubModule_SA_3D__zz_io_MatrixB_4_2 = SubModule_WeightCache_mData_34;
  assign SubModule_SA_3D__zz_io_B_Valid_4_2 = SubModule_WeightCache_MatrixCol_Switch[34];
  assign SubModule_SA_3D__zz_io_MatrixB_4_3 = SubModule_WeightCache_mData_35;
  assign SubModule_SA_3D__zz_io_B_Valid_4_3 = SubModule_WeightCache_MatrixCol_Switch[35];
  assign SubModule_SA_3D__zz_io_MatrixB_4_4 = SubModule_WeightCache_mData_36;
  assign SubModule_SA_3D__zz_io_B_Valid_4_4 = SubModule_WeightCache_MatrixCol_Switch[36];
  assign SubModule_SA_3D__zz_io_MatrixB_4_5 = SubModule_WeightCache_mData_37;
  assign SubModule_SA_3D__zz_io_B_Valid_4_5 = SubModule_WeightCache_MatrixCol_Switch[37];
  assign SubModule_SA_3D__zz_io_MatrixB_4_6 = SubModule_WeightCache_mData_38;
  assign SubModule_SA_3D__zz_io_B_Valid_4_6 = SubModule_WeightCache_MatrixCol_Switch[38];
  assign SubModule_SA_3D__zz_io_MatrixB_4_7 = SubModule_WeightCache_mData_39;
  assign SubModule_SA_3D__zz_io_B_Valid_4_7 = SubModule_WeightCache_MatrixCol_Switch[39];
  assign SubModule_SA_3D__zz_io_MatrixB_5 = SubModule_WeightCache_mData_40;
  assign SubModule_SA_3D__zz_io_B_Valid_5 = SubModule_WeightCache_MatrixCol_Switch[40];
  assign SubModule_SA_3D__zz_io_MatrixB_5_1 = SubModule_WeightCache_mData_41;
  assign SubModule_SA_3D__zz_io_B_Valid_5_1 = SubModule_WeightCache_MatrixCol_Switch[41];
  assign SubModule_SA_3D__zz_io_MatrixB_5_2 = SubModule_WeightCache_mData_42;
  assign SubModule_SA_3D__zz_io_B_Valid_5_2 = SubModule_WeightCache_MatrixCol_Switch[42];
  assign SubModule_SA_3D__zz_io_MatrixB_5_3 = SubModule_WeightCache_mData_43;
  assign SubModule_SA_3D__zz_io_B_Valid_5_3 = SubModule_WeightCache_MatrixCol_Switch[43];
  assign SubModule_SA_3D__zz_io_MatrixB_5_4 = SubModule_WeightCache_mData_44;
  assign SubModule_SA_3D__zz_io_B_Valid_5_4 = SubModule_WeightCache_MatrixCol_Switch[44];
  assign SubModule_SA_3D__zz_io_MatrixB_5_5 = SubModule_WeightCache_mData_45;
  assign SubModule_SA_3D__zz_io_B_Valid_5_5 = SubModule_WeightCache_MatrixCol_Switch[45];
  assign SubModule_SA_3D__zz_io_MatrixB_5_6 = SubModule_WeightCache_mData_46;
  assign SubModule_SA_3D__zz_io_B_Valid_5_6 = SubModule_WeightCache_MatrixCol_Switch[46];
  assign SubModule_SA_3D__zz_io_MatrixB_5_7 = SubModule_WeightCache_mData_47;
  assign SubModule_SA_3D__zz_io_B_Valid_5_7 = SubModule_WeightCache_MatrixCol_Switch[47];
  assign SubModule_SA_3D__zz_io_MatrixB_6 = SubModule_WeightCache_mData_48;
  assign SubModule_SA_3D__zz_io_B_Valid_6 = SubModule_WeightCache_MatrixCol_Switch[48];
  assign SubModule_SA_3D__zz_io_MatrixB_6_1 = SubModule_WeightCache_mData_49;
  assign SubModule_SA_3D__zz_io_B_Valid_6_1 = SubModule_WeightCache_MatrixCol_Switch[49];
  assign SubModule_SA_3D__zz_io_MatrixB_6_2 = SubModule_WeightCache_mData_50;
  assign SubModule_SA_3D__zz_io_B_Valid_6_2 = SubModule_WeightCache_MatrixCol_Switch[50];
  assign SubModule_SA_3D__zz_io_MatrixB_6_3 = SubModule_WeightCache_mData_51;
  assign SubModule_SA_3D__zz_io_B_Valid_6_3 = SubModule_WeightCache_MatrixCol_Switch[51];
  assign SubModule_SA_3D__zz_io_MatrixB_6_4 = SubModule_WeightCache_mData_52;
  assign SubModule_SA_3D__zz_io_B_Valid_6_4 = SubModule_WeightCache_MatrixCol_Switch[52];
  assign SubModule_SA_3D__zz_io_MatrixB_6_5 = SubModule_WeightCache_mData_53;
  assign SubModule_SA_3D__zz_io_B_Valid_6_5 = SubModule_WeightCache_MatrixCol_Switch[53];
  assign SubModule_SA_3D__zz_io_MatrixB_6_6 = SubModule_WeightCache_mData_54;
  assign SubModule_SA_3D__zz_io_B_Valid_6_6 = SubModule_WeightCache_MatrixCol_Switch[54];
  assign SubModule_SA_3D__zz_io_MatrixB_6_7 = SubModule_WeightCache_mData_55;
  assign SubModule_SA_3D__zz_io_B_Valid_6_7 = SubModule_WeightCache_MatrixCol_Switch[55];
  assign SubModule_SA_3D__zz_io_MatrixB_7 = SubModule_WeightCache_mData_56;
  assign SubModule_SA_3D__zz_io_B_Valid_7 = SubModule_WeightCache_MatrixCol_Switch[56];
  assign SubModule_SA_3D__zz_io_MatrixB_7_1 = SubModule_WeightCache_mData_57;
  assign SubModule_SA_3D__zz_io_B_Valid_7_1 = SubModule_WeightCache_MatrixCol_Switch[57];
  assign SubModule_SA_3D__zz_io_MatrixB_7_2 = SubModule_WeightCache_mData_58;
  assign SubModule_SA_3D__zz_io_B_Valid_7_2 = SubModule_WeightCache_MatrixCol_Switch[58];
  assign SubModule_SA_3D__zz_io_MatrixB_7_3 = SubModule_WeightCache_mData_59;
  assign SubModule_SA_3D__zz_io_B_Valid_7_3 = SubModule_WeightCache_MatrixCol_Switch[59];
  assign SubModule_SA_3D__zz_io_MatrixB_7_4 = SubModule_WeightCache_mData_60;
  assign SubModule_SA_3D__zz_io_B_Valid_7_4 = SubModule_WeightCache_MatrixCol_Switch[60];
  assign SubModule_SA_3D__zz_io_MatrixB_7_5 = SubModule_WeightCache_mData_61;
  assign SubModule_SA_3D__zz_io_B_Valid_7_5 = SubModule_WeightCache_MatrixCol_Switch[61];
  assign SubModule_SA_3D__zz_io_MatrixB_7_6 = SubModule_WeightCache_mData_62;
  assign SubModule_SA_3D__zz_io_B_Valid_7_6 = SubModule_WeightCache_MatrixCol_Switch[62];
  assign SubModule_SA_3D__zz_io_MatrixB_7_7 = SubModule_WeightCache_mData_63;
  assign SubModule_SA_3D__zz_io_B_Valid_7_7 = SubModule_WeightCache_MatrixCol_Switch[63];
  assign SubModule_Img2Col_start = (toplevel_SubModule_WeightCache_Weight_Cached_delay_3 && Control_Switch_Conv);
  assign Fsm_Picture_Received = SubModule_Img2Col_LayerEnd;
  assign Fsm_Switch_Conv = Control_Switch_Conv;
  assign Fsm_WeightCached = SubModule_WeightCache_Weight_Cached;
  always @(*) begin
    InputSwitch_m_0_axis_mm2s_tready = SubModule_WeightCache_s_axis_s2mm_tready;
    if(SubModule_WeightCache_s_axis_s2mm_tready) begin
      InputSwitch_m_0_axis_mm2s_tready = SubModule_WeightCache_s_axis_s2mm_tready;
    end else begin
      InputSwitch_m_0_axis_mm2s_tready = 1'b0;
    end
  end

  assign Fsm_Matrix_Received = 1'b0;
  assign LayerEnd = SubModule_Img2Col_LayerEnd;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= TopCtrl_Enum_IDLE;
      InitCnt_count <= 3'b000;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l19) begin
        InitCnt_count <= (InitCnt_count + 3'b001);
        if(InitCnt_valid) begin
          InitCnt_count <= 3'b000;
        end
      end
    end
  end

  always @(posedge clk) begin
    toplevel_SubModule_WeightCache_Weight_Cached_delay_1 <= SubModule_WeightCache_Weight_Cached;
    toplevel_SubModule_WeightCache_Weight_Cached_delay_2 <= toplevel_SubModule_WeightCache_Weight_Cached_delay_1;
    toplevel_SubModule_WeightCache_Weight_Cached_delay_3 <= toplevel_SubModule_WeightCache_Weight_Cached_delay_2;
    _zz_start <= ((Fsm_nextState & TopCtrl_Enum_WEIGHT_CACHE) != 6'b000000);
    _zz_start_1 <= _zz_start;
    _zz_start_2 <= _zz_start_1;
  end


endmodule

module WeightCache_Stream (
  input      [63:0]   s_axis_s2mm_tdata,
  input      [7:0]    s_axis_s2mm_tkeep,
  input               s_axis_s2mm_tlast,
  output              s_axis_s2mm_tready,
  input               s_axis_s2mm_tvalid,
  input               start,
  input      [15:0]   Matrix_Row,
  input      [15:0]   Matrix_Col,
  output     [7:0]    mData_0,
  output     [7:0]    mData_1,
  output     [7:0]    mData_2,
  output     [7:0]    mData_3,
  output     [7:0]    mData_4,
  output     [7:0]    mData_5,
  output     [7:0]    mData_6,
  output     [7:0]    mData_7,
  output     [7:0]    mData_8,
  output     [7:0]    mData_9,
  output     [7:0]    mData_10,
  output     [7:0]    mData_11,
  output     [7:0]    mData_12,
  output     [7:0]    mData_13,
  output     [7:0]    mData_14,
  output     [7:0]    mData_15,
  output     [7:0]    mData_16,
  output     [7:0]    mData_17,
  output     [7:0]    mData_18,
  output     [7:0]    mData_19,
  output     [7:0]    mData_20,
  output     [7:0]    mData_21,
  output     [7:0]    mData_22,
  output     [7:0]    mData_23,
  output     [7:0]    mData_24,
  output     [7:0]    mData_25,
  output     [7:0]    mData_26,
  output     [7:0]    mData_27,
  output     [7:0]    mData_28,
  output     [7:0]    mData_29,
  output     [7:0]    mData_30,
  output     [7:0]    mData_31,
  output     [7:0]    mData_32,
  output     [7:0]    mData_33,
  output     [7:0]    mData_34,
  output     [7:0]    mData_35,
  output     [7:0]    mData_36,
  output     [7:0]    mData_37,
  output     [7:0]    mData_38,
  output     [7:0]    mData_39,
  output     [7:0]    mData_40,
  output     [7:0]    mData_41,
  output     [7:0]    mData_42,
  output     [7:0]    mData_43,
  output     [7:0]    mData_44,
  output     [7:0]    mData_45,
  output     [7:0]    mData_46,
  output     [7:0]    mData_47,
  output     [7:0]    mData_48,
  output     [7:0]    mData_49,
  output     [7:0]    mData_50,
  output     [7:0]    mData_51,
  output     [7:0]    mData_52,
  output     [7:0]    mData_53,
  output     [7:0]    mData_54,
  output     [7:0]    mData_55,
  output     [7:0]    mData_56,
  output     [7:0]    mData_57,
  output     [7:0]    mData_58,
  output     [7:0]    mData_59,
  output     [7:0]    mData_60,
  output     [7:0]    mData_61,
  output     [7:0]    mData_62,
  output     [7:0]    mData_63,
  input               Raddr_Valid,
  output              Weight_Cached,
  input               LayerEnd,
  output     [63:0]   MatrixCol_Switch,
  input               clk,
  input               reset
);

  wire                WeightCache_sData_ready;
  wire       [7:0]    WeightCache_mData_0;
  wire       [7:0]    WeightCache_mData_1;
  wire       [7:0]    WeightCache_mData_2;
  wire       [7:0]    WeightCache_mData_3;
  wire       [7:0]    WeightCache_mData_4;
  wire       [7:0]    WeightCache_mData_5;
  wire       [7:0]    WeightCache_mData_6;
  wire       [7:0]    WeightCache_mData_7;
  wire       [7:0]    WeightCache_mData_8;
  wire       [7:0]    WeightCache_mData_9;
  wire       [7:0]    WeightCache_mData_10;
  wire       [7:0]    WeightCache_mData_11;
  wire       [7:0]    WeightCache_mData_12;
  wire       [7:0]    WeightCache_mData_13;
  wire       [7:0]    WeightCache_mData_14;
  wire       [7:0]    WeightCache_mData_15;
  wire       [7:0]    WeightCache_mData_16;
  wire       [7:0]    WeightCache_mData_17;
  wire       [7:0]    WeightCache_mData_18;
  wire       [7:0]    WeightCache_mData_19;
  wire       [7:0]    WeightCache_mData_20;
  wire       [7:0]    WeightCache_mData_21;
  wire       [7:0]    WeightCache_mData_22;
  wire       [7:0]    WeightCache_mData_23;
  wire       [7:0]    WeightCache_mData_24;
  wire       [7:0]    WeightCache_mData_25;
  wire       [7:0]    WeightCache_mData_26;
  wire       [7:0]    WeightCache_mData_27;
  wire       [7:0]    WeightCache_mData_28;
  wire       [7:0]    WeightCache_mData_29;
  wire       [7:0]    WeightCache_mData_30;
  wire       [7:0]    WeightCache_mData_31;
  wire       [7:0]    WeightCache_mData_32;
  wire       [7:0]    WeightCache_mData_33;
  wire       [7:0]    WeightCache_mData_34;
  wire       [7:0]    WeightCache_mData_35;
  wire       [7:0]    WeightCache_mData_36;
  wire       [7:0]    WeightCache_mData_37;
  wire       [7:0]    WeightCache_mData_38;
  wire       [7:0]    WeightCache_mData_39;
  wire       [7:0]    WeightCache_mData_40;
  wire       [7:0]    WeightCache_mData_41;
  wire       [7:0]    WeightCache_mData_42;
  wire       [7:0]    WeightCache_mData_43;
  wire       [7:0]    WeightCache_mData_44;
  wire       [7:0]    WeightCache_mData_45;
  wire       [7:0]    WeightCache_mData_46;
  wire       [7:0]    WeightCache_mData_47;
  wire       [7:0]    WeightCache_mData_48;
  wire       [7:0]    WeightCache_mData_49;
  wire       [7:0]    WeightCache_mData_50;
  wire       [7:0]    WeightCache_mData_51;
  wire       [7:0]    WeightCache_mData_52;
  wire       [7:0]    WeightCache_mData_53;
  wire       [7:0]    WeightCache_mData_54;
  wire       [7:0]    WeightCache_mData_55;
  wire       [7:0]    WeightCache_mData_56;
  wire       [7:0]    WeightCache_mData_57;
  wire       [7:0]    WeightCache_mData_58;
  wire       [7:0]    WeightCache_mData_59;
  wire       [7:0]    WeightCache_mData_60;
  wire       [7:0]    WeightCache_mData_61;
  wire       [7:0]    WeightCache_mData_62;
  wire       [7:0]    WeightCache_mData_63;
  wire                WeightCache_Weight_Cached;
  wire       [63:0]   WeightCache_MatrixCol_Switch;

  Weight_Cache WeightCache (
    .start            (start                             ), //i
    .sData_valid      (s_axis_s2mm_tvalid                ), //i
    .sData_ready      (WeightCache_sData_ready           ), //o
    .sData_payload    (s_axis_s2mm_tdata[63:0]           ), //i
    .Matrix_Row       (Matrix_Row[15:0]                  ), //i
    .Matrix_Col       (Matrix_Col[15:0]                  ), //i
    .mData_0          (WeightCache_mData_0[7:0]          ), //o
    .mData_1          (WeightCache_mData_1[7:0]          ), //o
    .mData_2          (WeightCache_mData_2[7:0]          ), //o
    .mData_3          (WeightCache_mData_3[7:0]          ), //o
    .mData_4          (WeightCache_mData_4[7:0]          ), //o
    .mData_5          (WeightCache_mData_5[7:0]          ), //o
    .mData_6          (WeightCache_mData_6[7:0]          ), //o
    .mData_7          (WeightCache_mData_7[7:0]          ), //o
    .mData_8          (WeightCache_mData_8[7:0]          ), //o
    .mData_9          (WeightCache_mData_9[7:0]          ), //o
    .mData_10         (WeightCache_mData_10[7:0]         ), //o
    .mData_11         (WeightCache_mData_11[7:0]         ), //o
    .mData_12         (WeightCache_mData_12[7:0]         ), //o
    .mData_13         (WeightCache_mData_13[7:0]         ), //o
    .mData_14         (WeightCache_mData_14[7:0]         ), //o
    .mData_15         (WeightCache_mData_15[7:0]         ), //o
    .mData_16         (WeightCache_mData_16[7:0]         ), //o
    .mData_17         (WeightCache_mData_17[7:0]         ), //o
    .mData_18         (WeightCache_mData_18[7:0]         ), //o
    .mData_19         (WeightCache_mData_19[7:0]         ), //o
    .mData_20         (WeightCache_mData_20[7:0]         ), //o
    .mData_21         (WeightCache_mData_21[7:0]         ), //o
    .mData_22         (WeightCache_mData_22[7:0]         ), //o
    .mData_23         (WeightCache_mData_23[7:0]         ), //o
    .mData_24         (WeightCache_mData_24[7:0]         ), //o
    .mData_25         (WeightCache_mData_25[7:0]         ), //o
    .mData_26         (WeightCache_mData_26[7:0]         ), //o
    .mData_27         (WeightCache_mData_27[7:0]         ), //o
    .mData_28         (WeightCache_mData_28[7:0]         ), //o
    .mData_29         (WeightCache_mData_29[7:0]         ), //o
    .mData_30         (WeightCache_mData_30[7:0]         ), //o
    .mData_31         (WeightCache_mData_31[7:0]         ), //o
    .mData_32         (WeightCache_mData_32[7:0]         ), //o
    .mData_33         (WeightCache_mData_33[7:0]         ), //o
    .mData_34         (WeightCache_mData_34[7:0]         ), //o
    .mData_35         (WeightCache_mData_35[7:0]         ), //o
    .mData_36         (WeightCache_mData_36[7:0]         ), //o
    .mData_37         (WeightCache_mData_37[7:0]         ), //o
    .mData_38         (WeightCache_mData_38[7:0]         ), //o
    .mData_39         (WeightCache_mData_39[7:0]         ), //o
    .mData_40         (WeightCache_mData_40[7:0]         ), //o
    .mData_41         (WeightCache_mData_41[7:0]         ), //o
    .mData_42         (WeightCache_mData_42[7:0]         ), //o
    .mData_43         (WeightCache_mData_43[7:0]         ), //o
    .mData_44         (WeightCache_mData_44[7:0]         ), //o
    .mData_45         (WeightCache_mData_45[7:0]         ), //o
    .mData_46         (WeightCache_mData_46[7:0]         ), //o
    .mData_47         (WeightCache_mData_47[7:0]         ), //o
    .mData_48         (WeightCache_mData_48[7:0]         ), //o
    .mData_49         (WeightCache_mData_49[7:0]         ), //o
    .mData_50         (WeightCache_mData_50[7:0]         ), //o
    .mData_51         (WeightCache_mData_51[7:0]         ), //o
    .mData_52         (WeightCache_mData_52[7:0]         ), //o
    .mData_53         (WeightCache_mData_53[7:0]         ), //o
    .mData_54         (WeightCache_mData_54[7:0]         ), //o
    .mData_55         (WeightCache_mData_55[7:0]         ), //o
    .mData_56         (WeightCache_mData_56[7:0]         ), //o
    .mData_57         (WeightCache_mData_57[7:0]         ), //o
    .mData_58         (WeightCache_mData_58[7:0]         ), //o
    .mData_59         (WeightCache_mData_59[7:0]         ), //o
    .mData_60         (WeightCache_mData_60[7:0]         ), //o
    .mData_61         (WeightCache_mData_61[7:0]         ), //o
    .mData_62         (WeightCache_mData_62[7:0]         ), //o
    .mData_63         (WeightCache_mData_63[7:0]         ), //o
    .Raddr_Valid      (Raddr_Valid                       ), //i
    .Weight_Cached    (WeightCache_Weight_Cached         ), //o
    .LayerEnd         (LayerEnd                          ), //i
    .MatrixCol_Switch (WeightCache_MatrixCol_Switch[63:0]), //o
    .clk              (clk                               ), //i
    .reset            (reset                             )  //i
  );
  assign mData_0 = WeightCache_mData_0;
  assign mData_1 = WeightCache_mData_1;
  assign mData_2 = WeightCache_mData_2;
  assign mData_3 = WeightCache_mData_3;
  assign mData_4 = WeightCache_mData_4;
  assign mData_5 = WeightCache_mData_5;
  assign mData_6 = WeightCache_mData_6;
  assign mData_7 = WeightCache_mData_7;
  assign mData_8 = WeightCache_mData_8;
  assign mData_9 = WeightCache_mData_9;
  assign mData_10 = WeightCache_mData_10;
  assign mData_11 = WeightCache_mData_11;
  assign mData_12 = WeightCache_mData_12;
  assign mData_13 = WeightCache_mData_13;
  assign mData_14 = WeightCache_mData_14;
  assign mData_15 = WeightCache_mData_15;
  assign mData_16 = WeightCache_mData_16;
  assign mData_17 = WeightCache_mData_17;
  assign mData_18 = WeightCache_mData_18;
  assign mData_19 = WeightCache_mData_19;
  assign mData_20 = WeightCache_mData_20;
  assign mData_21 = WeightCache_mData_21;
  assign mData_22 = WeightCache_mData_22;
  assign mData_23 = WeightCache_mData_23;
  assign mData_24 = WeightCache_mData_24;
  assign mData_25 = WeightCache_mData_25;
  assign mData_26 = WeightCache_mData_26;
  assign mData_27 = WeightCache_mData_27;
  assign mData_28 = WeightCache_mData_28;
  assign mData_29 = WeightCache_mData_29;
  assign mData_30 = WeightCache_mData_30;
  assign mData_31 = WeightCache_mData_31;
  assign mData_32 = WeightCache_mData_32;
  assign mData_33 = WeightCache_mData_33;
  assign mData_34 = WeightCache_mData_34;
  assign mData_35 = WeightCache_mData_35;
  assign mData_36 = WeightCache_mData_36;
  assign mData_37 = WeightCache_mData_37;
  assign mData_38 = WeightCache_mData_38;
  assign mData_39 = WeightCache_mData_39;
  assign mData_40 = WeightCache_mData_40;
  assign mData_41 = WeightCache_mData_41;
  assign mData_42 = WeightCache_mData_42;
  assign mData_43 = WeightCache_mData_43;
  assign mData_44 = WeightCache_mData_44;
  assign mData_45 = WeightCache_mData_45;
  assign mData_46 = WeightCache_mData_46;
  assign mData_47 = WeightCache_mData_47;
  assign mData_48 = WeightCache_mData_48;
  assign mData_49 = WeightCache_mData_49;
  assign mData_50 = WeightCache_mData_50;
  assign mData_51 = WeightCache_mData_51;
  assign mData_52 = WeightCache_mData_52;
  assign mData_53 = WeightCache_mData_53;
  assign mData_54 = WeightCache_mData_54;
  assign mData_55 = WeightCache_mData_55;
  assign mData_56 = WeightCache_mData_56;
  assign mData_57 = WeightCache_mData_57;
  assign mData_58 = WeightCache_mData_58;
  assign mData_59 = WeightCache_mData_59;
  assign mData_60 = WeightCache_mData_60;
  assign mData_61 = WeightCache_mData_61;
  assign mData_62 = WeightCache_mData_62;
  assign mData_63 = WeightCache_mData_63;
  assign Weight_Cached = WeightCache_Weight_Cached;
  assign MatrixCol_Switch = WeightCache_MatrixCol_Switch;
  assign s_axis_s2mm_tready = WeightCache_sData_ready;

endmodule

module SA_3D (
  input      [7:0]    _zz_io_MatrixA_0,
  input      [7:0]    _zz_io_MatrixA_1,
  input      [7:0]    _zz_io_MatrixA_2,
  input      [7:0]    _zz_io_MatrixA_3,
  input      [7:0]    _zz_io_MatrixA_4,
  input      [7:0]    _zz_io_MatrixA_5,
  input      [7:0]    _zz_io_MatrixA_6,
  input      [7:0]    _zz_io_MatrixA_7,
  input      [7:0]    _zz_io_MatrixB_0,
  input      [7:0]    _zz_io_MatrixB_1,
  input      [7:0]    _zz_io_MatrixB_2,
  input      [7:0]    _zz_io_MatrixB_3,
  input      [7:0]    _zz_io_MatrixB_4,
  input      [7:0]    _zz_io_MatrixB_5,
  input      [7:0]    _zz_io_MatrixB_6,
  input      [7:0]    _zz_io_MatrixB_7,
  input               _zz_io_A_Valid_0,
  input               _zz_io_A_Valid_1,
  input               _zz_io_A_Valid_2,
  input               _zz_io_A_Valid_3,
  input               _zz_io_A_Valid_4,
  input               _zz_io_A_Valid_5,
  input               _zz_io_A_Valid_6,
  input               _zz_io_A_Valid_7,
  input               _zz_io_B_Valid_0,
  input               _zz_io_B_Valid_1,
  input               _zz_io_B_Valid_2,
  input               _zz_io_B_Valid_3,
  input               _zz_io_B_Valid_4,
  input               _zz_io_B_Valid_5,
  input               _zz_io_B_Valid_6,
  input               _zz_io_B_Valid_7,
  input      [15:0]   _zz_io_signCount,
  input               clk,
  input      [7:0]    _zz_io_MatrixA_0_1,
  input      [7:0]    _zz_io_MatrixA_1_1,
  input      [7:0]    _zz_io_MatrixA_2_1,
  input      [7:0]    _zz_io_MatrixA_3_1,
  input      [7:0]    _zz_io_MatrixA_4_1,
  input      [7:0]    _zz_io_MatrixA_5_1,
  input      [7:0]    _zz_io_MatrixA_6_1,
  input      [7:0]    _zz_io_MatrixA_7_1,
  input      [7:0]    _zz_io_MatrixB_0_1,
  input      [7:0]    _zz_io_MatrixB_1_1,
  input      [7:0]    _zz_io_MatrixB_2_1,
  input      [7:0]    _zz_io_MatrixB_3_1,
  input      [7:0]    _zz_io_MatrixB_4_1,
  input      [7:0]    _zz_io_MatrixB_5_1,
  input      [7:0]    _zz_io_MatrixB_6_1,
  input      [7:0]    _zz_io_MatrixB_7_1,
  input               _zz_io_A_Valid_0_1,
  input               _zz_io_A_Valid_1_1,
  input               _zz_io_A_Valid_2_1,
  input               _zz_io_A_Valid_3_1,
  input               _zz_io_A_Valid_4_1,
  input               _zz_io_A_Valid_5_1,
  input               _zz_io_A_Valid_6_1,
  input               _zz_io_A_Valid_7_1,
  input               _zz_io_B_Valid_0_1,
  input               _zz_io_B_Valid_1_1,
  input               _zz_io_B_Valid_2_1,
  input               _zz_io_B_Valid_3_1,
  input               _zz_io_B_Valid_4_1,
  input               _zz_io_B_Valid_5_1,
  input               _zz_io_B_Valid_6_1,
  input               _zz_io_B_Valid_7_1,
  input      [15:0]   _zz_io_signCount_1,
  input      [7:0]    _zz_io_MatrixA_0_2,
  input      [7:0]    _zz_io_MatrixA_1_2,
  input      [7:0]    _zz_io_MatrixA_2_2,
  input      [7:0]    _zz_io_MatrixA_3_2,
  input      [7:0]    _zz_io_MatrixA_4_2,
  input      [7:0]    _zz_io_MatrixA_5_2,
  input      [7:0]    _zz_io_MatrixA_6_2,
  input      [7:0]    _zz_io_MatrixA_7_2,
  input      [7:0]    _zz_io_MatrixB_0_2,
  input      [7:0]    _zz_io_MatrixB_1_2,
  input      [7:0]    _zz_io_MatrixB_2_2,
  input      [7:0]    _zz_io_MatrixB_3_2,
  input      [7:0]    _zz_io_MatrixB_4_2,
  input      [7:0]    _zz_io_MatrixB_5_2,
  input      [7:0]    _zz_io_MatrixB_6_2,
  input      [7:0]    _zz_io_MatrixB_7_2,
  input               _zz_io_A_Valid_0_2,
  input               _zz_io_A_Valid_1_2,
  input               _zz_io_A_Valid_2_2,
  input               _zz_io_A_Valid_3_2,
  input               _zz_io_A_Valid_4_2,
  input               _zz_io_A_Valid_5_2,
  input               _zz_io_A_Valid_6_2,
  input               _zz_io_A_Valid_7_2,
  input               _zz_io_B_Valid_0_2,
  input               _zz_io_B_Valid_1_2,
  input               _zz_io_B_Valid_2_2,
  input               _zz_io_B_Valid_3_2,
  input               _zz_io_B_Valid_4_2,
  input               _zz_io_B_Valid_5_2,
  input               _zz_io_B_Valid_6_2,
  input               _zz_io_B_Valid_7_2,
  input      [15:0]   _zz_io_signCount_2,
  input      [7:0]    _zz_io_MatrixA_0_3,
  input      [7:0]    _zz_io_MatrixA_1_3,
  input      [7:0]    _zz_io_MatrixA_2_3,
  input      [7:0]    _zz_io_MatrixA_3_3,
  input      [7:0]    _zz_io_MatrixA_4_3,
  input      [7:0]    _zz_io_MatrixA_5_3,
  input      [7:0]    _zz_io_MatrixA_6_3,
  input      [7:0]    _zz_io_MatrixA_7_3,
  input      [7:0]    _zz_io_MatrixB_0_3,
  input      [7:0]    _zz_io_MatrixB_1_3,
  input      [7:0]    _zz_io_MatrixB_2_3,
  input      [7:0]    _zz_io_MatrixB_3_3,
  input      [7:0]    _zz_io_MatrixB_4_3,
  input      [7:0]    _zz_io_MatrixB_5_3,
  input      [7:0]    _zz_io_MatrixB_6_3,
  input      [7:0]    _zz_io_MatrixB_7_3,
  input               _zz_io_A_Valid_0_3,
  input               _zz_io_A_Valid_1_3,
  input               _zz_io_A_Valid_2_3,
  input               _zz_io_A_Valid_3_3,
  input               _zz_io_A_Valid_4_3,
  input               _zz_io_A_Valid_5_3,
  input               _zz_io_A_Valid_6_3,
  input               _zz_io_A_Valid_7_3,
  input               _zz_io_B_Valid_0_3,
  input               _zz_io_B_Valid_1_3,
  input               _zz_io_B_Valid_2_3,
  input               _zz_io_B_Valid_3_3,
  input               _zz_io_B_Valid_4_3,
  input               _zz_io_B_Valid_5_3,
  input               _zz_io_B_Valid_6_3,
  input               _zz_io_B_Valid_7_3,
  input      [15:0]   _zz_io_signCount_3,
  input      [7:0]    _zz_io_MatrixA_0_4,
  input      [7:0]    _zz_io_MatrixA_1_4,
  input      [7:0]    _zz_io_MatrixA_2_4,
  input      [7:0]    _zz_io_MatrixA_3_4,
  input      [7:0]    _zz_io_MatrixA_4_4,
  input      [7:0]    _zz_io_MatrixA_5_4,
  input      [7:0]    _zz_io_MatrixA_6_4,
  input      [7:0]    _zz_io_MatrixA_7_4,
  input      [7:0]    _zz_io_MatrixB_0_4,
  input      [7:0]    _zz_io_MatrixB_1_4,
  input      [7:0]    _zz_io_MatrixB_2_4,
  input      [7:0]    _zz_io_MatrixB_3_4,
  input      [7:0]    _zz_io_MatrixB_4_4,
  input      [7:0]    _zz_io_MatrixB_5_4,
  input      [7:0]    _zz_io_MatrixB_6_4,
  input      [7:0]    _zz_io_MatrixB_7_4,
  input               _zz_io_A_Valid_0_4,
  input               _zz_io_A_Valid_1_4,
  input               _zz_io_A_Valid_2_4,
  input               _zz_io_A_Valid_3_4,
  input               _zz_io_A_Valid_4_4,
  input               _zz_io_A_Valid_5_4,
  input               _zz_io_A_Valid_6_4,
  input               _zz_io_A_Valid_7_4,
  input               _zz_io_B_Valid_0_4,
  input               _zz_io_B_Valid_1_4,
  input               _zz_io_B_Valid_2_4,
  input               _zz_io_B_Valid_3_4,
  input               _zz_io_B_Valid_4_4,
  input               _zz_io_B_Valid_5_4,
  input               _zz_io_B_Valid_6_4,
  input               _zz_io_B_Valid_7_4,
  input      [15:0]   _zz_io_signCount_4,
  input      [7:0]    _zz_io_MatrixA_0_5,
  input      [7:0]    _zz_io_MatrixA_1_5,
  input      [7:0]    _zz_io_MatrixA_2_5,
  input      [7:0]    _zz_io_MatrixA_3_5,
  input      [7:0]    _zz_io_MatrixA_4_5,
  input      [7:0]    _zz_io_MatrixA_5_5,
  input      [7:0]    _zz_io_MatrixA_6_5,
  input      [7:0]    _zz_io_MatrixA_7_5,
  input      [7:0]    _zz_io_MatrixB_0_5,
  input      [7:0]    _zz_io_MatrixB_1_5,
  input      [7:0]    _zz_io_MatrixB_2_5,
  input      [7:0]    _zz_io_MatrixB_3_5,
  input      [7:0]    _zz_io_MatrixB_4_5,
  input      [7:0]    _zz_io_MatrixB_5_5,
  input      [7:0]    _zz_io_MatrixB_6_5,
  input      [7:0]    _zz_io_MatrixB_7_5,
  input               _zz_io_A_Valid_0_5,
  input               _zz_io_A_Valid_1_5,
  input               _zz_io_A_Valid_2_5,
  input               _zz_io_A_Valid_3_5,
  input               _zz_io_A_Valid_4_5,
  input               _zz_io_A_Valid_5_5,
  input               _zz_io_A_Valid_6_5,
  input               _zz_io_A_Valid_7_5,
  input               _zz_io_B_Valid_0_5,
  input               _zz_io_B_Valid_1_5,
  input               _zz_io_B_Valid_2_5,
  input               _zz_io_B_Valid_3_5,
  input               _zz_io_B_Valid_4_5,
  input               _zz_io_B_Valid_5_5,
  input               _zz_io_B_Valid_6_5,
  input               _zz_io_B_Valid_7_5,
  input      [15:0]   _zz_io_signCount_5,
  input      [7:0]    _zz_io_MatrixA_0_6,
  input      [7:0]    _zz_io_MatrixA_1_6,
  input      [7:0]    _zz_io_MatrixA_2_6,
  input      [7:0]    _zz_io_MatrixA_3_6,
  input      [7:0]    _zz_io_MatrixA_4_6,
  input      [7:0]    _zz_io_MatrixA_5_6,
  input      [7:0]    _zz_io_MatrixA_6_6,
  input      [7:0]    _zz_io_MatrixA_7_6,
  input      [7:0]    _zz_io_MatrixB_0_6,
  input      [7:0]    _zz_io_MatrixB_1_6,
  input      [7:0]    _zz_io_MatrixB_2_6,
  input      [7:0]    _zz_io_MatrixB_3_6,
  input      [7:0]    _zz_io_MatrixB_4_6,
  input      [7:0]    _zz_io_MatrixB_5_6,
  input      [7:0]    _zz_io_MatrixB_6_6,
  input      [7:0]    _zz_io_MatrixB_7_6,
  input               _zz_io_A_Valid_0_6,
  input               _zz_io_A_Valid_1_6,
  input               _zz_io_A_Valid_2_6,
  input               _zz_io_A_Valid_3_6,
  input               _zz_io_A_Valid_4_6,
  input               _zz_io_A_Valid_5_6,
  input               _zz_io_A_Valid_6_6,
  input               _zz_io_A_Valid_7_6,
  input               _zz_io_B_Valid_0_6,
  input               _zz_io_B_Valid_1_6,
  input               _zz_io_B_Valid_2_6,
  input               _zz_io_B_Valid_3_6,
  input               _zz_io_B_Valid_4_6,
  input               _zz_io_B_Valid_5_6,
  input               _zz_io_B_Valid_6_6,
  input               _zz_io_B_Valid_7_6,
  input      [15:0]   _zz_io_signCount_6,
  input      [7:0]    _zz_io_MatrixA_0_7,
  input      [7:0]    _zz_io_MatrixA_1_7,
  input      [7:0]    _zz_io_MatrixA_2_7,
  input      [7:0]    _zz_io_MatrixA_3_7,
  input      [7:0]    _zz_io_MatrixA_4_7,
  input      [7:0]    _zz_io_MatrixA_5_7,
  input      [7:0]    _zz_io_MatrixA_6_7,
  input      [7:0]    _zz_io_MatrixA_7_7,
  input      [7:0]    _zz_io_MatrixB_0_7,
  input      [7:0]    _zz_io_MatrixB_1_7,
  input      [7:0]    _zz_io_MatrixB_2_7,
  input      [7:0]    _zz_io_MatrixB_3_7,
  input      [7:0]    _zz_io_MatrixB_4_7,
  input      [7:0]    _zz_io_MatrixB_5_7,
  input      [7:0]    _zz_io_MatrixB_6_7,
  input      [7:0]    _zz_io_MatrixB_7_7,
  input               _zz_io_A_Valid_0_7,
  input               _zz_io_A_Valid_1_7,
  input               _zz_io_A_Valid_2_7,
  input               _zz_io_A_Valid_3_7,
  input               _zz_io_A_Valid_4_7,
  input               _zz_io_A_Valid_5_7,
  input               _zz_io_A_Valid_6_7,
  input               _zz_io_A_Valid_7_7,
  input               _zz_io_B_Valid_0_7,
  input               _zz_io_B_Valid_1_7,
  input               _zz_io_B_Valid_2_7,
  input               _zz_io_B_Valid_3_7,
  input               _zz_io_B_Valid_4_7,
  input               _zz_io_B_Valid_5_7,
  input               _zz_io_B_Valid_6_7,
  input               _zz_io_B_Valid_7_7,
  input      [15:0]   _zz_io_signCount_7,
  input               reset
);

  wire                sA_2D_8_start;
  wire                sA_2D_9_start;
  wire                sA_2D_10_start;
  wire                sA_2D_11_start;
  wire                sA_2D_12_start;
  wire                sA_2D_13_start;
  wire                sA_2D_14_start;
  wire                sA_2D_15_start;
  wire       [31:0]   sA_2D_8_MatrixC_0;
  wire       [31:0]   sA_2D_8_MatrixC_1;
  wire       [31:0]   sA_2D_8_MatrixC_2;
  wire       [31:0]   sA_2D_8_MatrixC_3;
  wire       [31:0]   sA_2D_8_MatrixC_4;
  wire       [31:0]   sA_2D_8_MatrixC_5;
  wire       [31:0]   sA_2D_8_MatrixC_6;
  wire       [31:0]   sA_2D_8_MatrixC_7;
  wire                sA_2D_8_C_Valid_0;
  wire                sA_2D_8_C_Valid_1;
  wire                sA_2D_8_C_Valid_2;
  wire                sA_2D_8_C_Valid_3;
  wire                sA_2D_8_C_Valid_4;
  wire                sA_2D_8_C_Valid_5;
  wire                sA_2D_8_C_Valid_6;
  wire                sA_2D_8_C_Valid_7;
  wire       [31:0]   sA_2D_9_MatrixC_0;
  wire       [31:0]   sA_2D_9_MatrixC_1;
  wire       [31:0]   sA_2D_9_MatrixC_2;
  wire       [31:0]   sA_2D_9_MatrixC_3;
  wire       [31:0]   sA_2D_9_MatrixC_4;
  wire       [31:0]   sA_2D_9_MatrixC_5;
  wire       [31:0]   sA_2D_9_MatrixC_6;
  wire       [31:0]   sA_2D_9_MatrixC_7;
  wire                sA_2D_9_C_Valid_0;
  wire                sA_2D_9_C_Valid_1;
  wire                sA_2D_9_C_Valid_2;
  wire                sA_2D_9_C_Valid_3;
  wire                sA_2D_9_C_Valid_4;
  wire                sA_2D_9_C_Valid_5;
  wire                sA_2D_9_C_Valid_6;
  wire                sA_2D_9_C_Valid_7;
  wire       [31:0]   sA_2D_10_MatrixC_0;
  wire       [31:0]   sA_2D_10_MatrixC_1;
  wire       [31:0]   sA_2D_10_MatrixC_2;
  wire       [31:0]   sA_2D_10_MatrixC_3;
  wire       [31:0]   sA_2D_10_MatrixC_4;
  wire       [31:0]   sA_2D_10_MatrixC_5;
  wire       [31:0]   sA_2D_10_MatrixC_6;
  wire       [31:0]   sA_2D_10_MatrixC_7;
  wire                sA_2D_10_C_Valid_0;
  wire                sA_2D_10_C_Valid_1;
  wire                sA_2D_10_C_Valid_2;
  wire                sA_2D_10_C_Valid_3;
  wire                sA_2D_10_C_Valid_4;
  wire                sA_2D_10_C_Valid_5;
  wire                sA_2D_10_C_Valid_6;
  wire                sA_2D_10_C_Valid_7;
  wire       [31:0]   sA_2D_11_MatrixC_0;
  wire       [31:0]   sA_2D_11_MatrixC_1;
  wire       [31:0]   sA_2D_11_MatrixC_2;
  wire       [31:0]   sA_2D_11_MatrixC_3;
  wire       [31:0]   sA_2D_11_MatrixC_4;
  wire       [31:0]   sA_2D_11_MatrixC_5;
  wire       [31:0]   sA_2D_11_MatrixC_6;
  wire       [31:0]   sA_2D_11_MatrixC_7;
  wire                sA_2D_11_C_Valid_0;
  wire                sA_2D_11_C_Valid_1;
  wire                sA_2D_11_C_Valid_2;
  wire                sA_2D_11_C_Valid_3;
  wire                sA_2D_11_C_Valid_4;
  wire                sA_2D_11_C_Valid_5;
  wire                sA_2D_11_C_Valid_6;
  wire                sA_2D_11_C_Valid_7;
  wire       [31:0]   sA_2D_12_MatrixC_0;
  wire       [31:0]   sA_2D_12_MatrixC_1;
  wire       [31:0]   sA_2D_12_MatrixC_2;
  wire       [31:0]   sA_2D_12_MatrixC_3;
  wire       [31:0]   sA_2D_12_MatrixC_4;
  wire       [31:0]   sA_2D_12_MatrixC_5;
  wire       [31:0]   sA_2D_12_MatrixC_6;
  wire       [31:0]   sA_2D_12_MatrixC_7;
  wire                sA_2D_12_C_Valid_0;
  wire                sA_2D_12_C_Valid_1;
  wire                sA_2D_12_C_Valid_2;
  wire                sA_2D_12_C_Valid_3;
  wire                sA_2D_12_C_Valid_4;
  wire                sA_2D_12_C_Valid_5;
  wire                sA_2D_12_C_Valid_6;
  wire                sA_2D_12_C_Valid_7;
  wire       [31:0]   sA_2D_13_MatrixC_0;
  wire       [31:0]   sA_2D_13_MatrixC_1;
  wire       [31:0]   sA_2D_13_MatrixC_2;
  wire       [31:0]   sA_2D_13_MatrixC_3;
  wire       [31:0]   sA_2D_13_MatrixC_4;
  wire       [31:0]   sA_2D_13_MatrixC_5;
  wire       [31:0]   sA_2D_13_MatrixC_6;
  wire       [31:0]   sA_2D_13_MatrixC_7;
  wire                sA_2D_13_C_Valid_0;
  wire                sA_2D_13_C_Valid_1;
  wire                sA_2D_13_C_Valid_2;
  wire                sA_2D_13_C_Valid_3;
  wire                sA_2D_13_C_Valid_4;
  wire                sA_2D_13_C_Valid_5;
  wire                sA_2D_13_C_Valid_6;
  wire                sA_2D_13_C_Valid_7;
  wire       [31:0]   sA_2D_14_MatrixC_0;
  wire       [31:0]   sA_2D_14_MatrixC_1;
  wire       [31:0]   sA_2D_14_MatrixC_2;
  wire       [31:0]   sA_2D_14_MatrixC_3;
  wire       [31:0]   sA_2D_14_MatrixC_4;
  wire       [31:0]   sA_2D_14_MatrixC_5;
  wire       [31:0]   sA_2D_14_MatrixC_6;
  wire       [31:0]   sA_2D_14_MatrixC_7;
  wire                sA_2D_14_C_Valid_0;
  wire                sA_2D_14_C_Valid_1;
  wire                sA_2D_14_C_Valid_2;
  wire                sA_2D_14_C_Valid_3;
  wire                sA_2D_14_C_Valid_4;
  wire                sA_2D_14_C_Valid_5;
  wire                sA_2D_14_C_Valid_6;
  wire                sA_2D_14_C_Valid_7;
  wire       [31:0]   sA_2D_15_MatrixC_0;
  wire       [31:0]   sA_2D_15_MatrixC_1;
  wire       [31:0]   sA_2D_15_MatrixC_2;
  wire       [31:0]   sA_2D_15_MatrixC_3;
  wire       [31:0]   sA_2D_15_MatrixC_4;
  wire       [31:0]   sA_2D_15_MatrixC_5;
  wire       [31:0]   sA_2D_15_MatrixC_6;
  wire       [31:0]   sA_2D_15_MatrixC_7;
  wire                sA_2D_15_C_Valid_0;
  wire                sA_2D_15_C_Valid_1;
  wire                sA_2D_15_C_Valid_2;
  wire                sA_2D_15_C_Valid_3;
  wire                sA_2D_15_C_Valid_4;
  wire                sA_2D_15_C_Valid_5;
  wire                sA_2D_15_C_Valid_6;
  wire                sA_2D_15_C_Valid_7;

  SA_2D sA_2D_8 (
    .io_MatrixA_0 (_zz_io_MatrixA_0[7:0]  ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1[7:0]  ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2[7:0]  ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3[7:0]  ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4[7:0]  ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5[7:0]  ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6[7:0]  ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7[7:0]  ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0[7:0]  ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1[7:0]  ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2[7:0]  ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3[7:0]  ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4[7:0]  ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5[7:0]  ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6[7:0]  ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7[7:0]  ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0       ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1       ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2       ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3       ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4       ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5       ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6       ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7       ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0       ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1       ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2       ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3       ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4       ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5       ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6       ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7       ), //i
    .io_signCount (_zz_io_signCount[15:0] ), //i
    .MatrixC_0    (sA_2D_8_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_8_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_8_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_8_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_8_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_8_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_8_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_8_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_8_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_8_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_8_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_8_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_8_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_8_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_8_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_8_C_Valid_7      ), //o
    .start        (sA_2D_8_start          ), //i
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  SA_2D sA_2D_9 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_1[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_1[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_1[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_1[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_1[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_1[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_1[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_1[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_1[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_1[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_1[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_1[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_1[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_1[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_1[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_1[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_1      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_1      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_1      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_1      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_1      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_1      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_1      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_1      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_1      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_1      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_1      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_1      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_1      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_1      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_1      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_1      ), //i
    .io_signCount (_zz_io_signCount_1[15:0]), //i
    .MatrixC_0    (sA_2D_9_MatrixC_0[31:0] ), //o
    .MatrixC_1    (sA_2D_9_MatrixC_1[31:0] ), //o
    .MatrixC_2    (sA_2D_9_MatrixC_2[31:0] ), //o
    .MatrixC_3    (sA_2D_9_MatrixC_3[31:0] ), //o
    .MatrixC_4    (sA_2D_9_MatrixC_4[31:0] ), //o
    .MatrixC_5    (sA_2D_9_MatrixC_5[31:0] ), //o
    .MatrixC_6    (sA_2D_9_MatrixC_6[31:0] ), //o
    .MatrixC_7    (sA_2D_9_MatrixC_7[31:0] ), //o
    .C_Valid_0    (sA_2D_9_C_Valid_0       ), //o
    .C_Valid_1    (sA_2D_9_C_Valid_1       ), //o
    .C_Valid_2    (sA_2D_9_C_Valid_2       ), //o
    .C_Valid_3    (sA_2D_9_C_Valid_3       ), //o
    .C_Valid_4    (sA_2D_9_C_Valid_4       ), //o
    .C_Valid_5    (sA_2D_9_C_Valid_5       ), //o
    .C_Valid_6    (sA_2D_9_C_Valid_6       ), //o
    .C_Valid_7    (sA_2D_9_C_Valid_7       ), //o
    .start        (sA_2D_9_start           ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );
  SA_2D sA_2D_10 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_2[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_2[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_2[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_2[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_2[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_2[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_2[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_2[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_2[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_2[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_2[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_2[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_2[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_2[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_2[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_2[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_2      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_2      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_2      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_2      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_2      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_2      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_2      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_2      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_2      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_2      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_2      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_2      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_2      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_2      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_2      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_2      ), //i
    .io_signCount (_zz_io_signCount_2[15:0]), //i
    .MatrixC_0    (sA_2D_10_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_10_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_10_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_10_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_10_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_10_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_10_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_10_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_10_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_10_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_10_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_10_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_10_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_10_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_10_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_10_C_Valid_7      ), //o
    .start        (sA_2D_10_start          ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );
  SA_2D sA_2D_11 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_3[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_3[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_3[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_3[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_3[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_3[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_3[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_3[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_3[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_3[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_3[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_3[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_3[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_3[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_3[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_3[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_3      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_3      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_3      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_3      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_3      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_3      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_3      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_3      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_3      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_3      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_3      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_3      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_3      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_3      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_3      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_3      ), //i
    .io_signCount (_zz_io_signCount_3[15:0]), //i
    .MatrixC_0    (sA_2D_11_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_11_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_11_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_11_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_11_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_11_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_11_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_11_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_11_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_11_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_11_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_11_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_11_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_11_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_11_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_11_C_Valid_7      ), //o
    .start        (sA_2D_11_start          ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );
  SA_2D sA_2D_12 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_4[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_4[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_4[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_4[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_4[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_4[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_4[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_4[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_4[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_4[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_4[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_4[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_4[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_4[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_4[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_4[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_4      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_4      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_4      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_4      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_4      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_4      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_4      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_4      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_4      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_4      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_4      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_4      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_4      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_4      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_4      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_4      ), //i
    .io_signCount (_zz_io_signCount_4[15:0]), //i
    .MatrixC_0    (sA_2D_12_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_12_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_12_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_12_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_12_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_12_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_12_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_12_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_12_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_12_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_12_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_12_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_12_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_12_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_12_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_12_C_Valid_7      ), //o
    .start        (sA_2D_12_start          ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );
  SA_2D sA_2D_13 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_5[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_5[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_5[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_5[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_5[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_5[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_5[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_5[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_5[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_5[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_5[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_5[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_5[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_5[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_5[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_5[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_5      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_5      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_5      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_5      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_5      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_5      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_5      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_5      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_5      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_5      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_5      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_5      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_5      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_5      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_5      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_5      ), //i
    .io_signCount (_zz_io_signCount_5[15:0]), //i
    .MatrixC_0    (sA_2D_13_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_13_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_13_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_13_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_13_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_13_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_13_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_13_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_13_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_13_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_13_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_13_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_13_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_13_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_13_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_13_C_Valid_7      ), //o
    .start        (sA_2D_13_start          ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );
  SA_2D sA_2D_14 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_6[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_6[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_6[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_6[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_6[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_6[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_6[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_6[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_6[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_6[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_6[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_6[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_6[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_6[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_6[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_6[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_6      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_6      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_6      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_6      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_6      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_6      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_6      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_6      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_6      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_6      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_6      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_6      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_6      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_6      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_6      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_6      ), //i
    .io_signCount (_zz_io_signCount_6[15:0]), //i
    .MatrixC_0    (sA_2D_14_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_14_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_14_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_14_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_14_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_14_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_14_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_14_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_14_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_14_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_14_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_14_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_14_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_14_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_14_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_14_C_Valid_7      ), //o
    .start        (sA_2D_14_start          ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );
  SA_2D sA_2D_15 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_7[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_7[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_7[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_7[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_7[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_7[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_7[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_7[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_7[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_7[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_7[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_7[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_7[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_7[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_7[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_7[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_7      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_7      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_7      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_7      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_7      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_7      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_7      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_7      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_7      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_7      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_7      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_7      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_7      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_7      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_7      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_7      ), //i
    .io_signCount (_zz_io_signCount_7[15:0]), //i
    .MatrixC_0    (sA_2D_15_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_15_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_15_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_15_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_15_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_15_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_15_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_15_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_15_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_15_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_15_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_15_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_15_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_15_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_15_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_15_C_Valid_7      ), //o
    .start        (sA_2D_15_start          ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );

endmodule

module Img2ColStreamV2 (
  output reg [63:0]   mData,
  output reg [7:0]    mValid,
  input      [63:0]   s_axis_s2mm_tdata,
  input      [7:0]    s_axis_s2mm_tkeep,
  input               s_axis_s2mm_tlast,
  output              s_axis_s2mm_tready,
  input               s_axis_s2mm_tvalid,
  input               start,
  output              Raddr_Valid,
  output              LayerEnd,
  input      [4:0]    Stride,
  input      [4:0]    Kernel_Size,
  input      [15:0]   Window_Size,
  input      [15:0]   InFeature_Size,
  input      [15:0]   InFeature_Channel,
  input      [15:0]   OutFeature_Channel,
  input      [15:0]   OutFeature_Size,
  input      [15:0]   OutCol_Count_Times,
  input      [15:0]   InCol_Count_Times,
  input      [15:0]   OutRow_Count_Times,
  input      [15:0]   OutFeature_Channel_Count_Times,
  input      [12:0]   Sliding_Size,
  input               clk,
  input               reset
);

  wire                SubModule_Fifo_Clear;
  wire       [15:0]   SubModule_Test_Generate_Period;
  wire                streamFifo_io_push_valid;
  wire                streamFifo_1_io_push_valid;
  wire                streamFifo_2_io_push_valid;
  wire                streamFifo_3_io_push_valid;
  wire                streamFifo_4_io_push_valid;
  wire                streamFifo_5_io_push_valid;
  wire                streamFifo_6_io_push_valid;
  wire                streamFifo_7_io_push_valid;
  wire                SubModule_sData_ready;
  wire       [63:0]   SubModule_mData;
  wire                SubModule_mValid;
  wire                SubModule_mLast;
  wire                SubModule_Test_Signal;
  wire                SubModule_Test_End;
  wire                SubModule_Raddr_Valid;
  wire                SubModule_LayerEnd;
  wire                SubModule_SA_Row_Cnt_Valid;
  wire                streamFifo_io_push_ready;
  wire                streamFifo_io_pop_valid;
  wire       [63:0]   streamFifo_io_pop_payload;
  wire       [4:0]    streamFifo_io_occupancy;
  wire       [4:0]    streamFifo_io_availability;
  wire                axisDataConverter_8_inStream_ready;
  wire                axisDataConverter_8_outStream_valid;
  wire       [7:0]    axisDataConverter_8_outStream_payload;
  wire                streamFifo_1_io_push_ready;
  wire                streamFifo_1_io_pop_valid;
  wire       [63:0]   streamFifo_1_io_pop_payload;
  wire       [4:0]    streamFifo_1_io_occupancy;
  wire       [4:0]    streamFifo_1_io_availability;
  wire                axisDataConverter_9_inStream_ready;
  wire                axisDataConverter_9_outStream_valid;
  wire       [7:0]    axisDataConverter_9_outStream_payload;
  wire                streamFifo_2_io_push_ready;
  wire                streamFifo_2_io_pop_valid;
  wire       [63:0]   streamFifo_2_io_pop_payload;
  wire       [4:0]    streamFifo_2_io_occupancy;
  wire       [4:0]    streamFifo_2_io_availability;
  wire                axisDataConverter_10_inStream_ready;
  wire                axisDataConverter_10_outStream_valid;
  wire       [7:0]    axisDataConverter_10_outStream_payload;
  wire                streamFifo_3_io_push_ready;
  wire                streamFifo_3_io_pop_valid;
  wire       [63:0]   streamFifo_3_io_pop_payload;
  wire       [4:0]    streamFifo_3_io_occupancy;
  wire       [4:0]    streamFifo_3_io_availability;
  wire                axisDataConverter_11_inStream_ready;
  wire                axisDataConverter_11_outStream_valid;
  wire       [7:0]    axisDataConverter_11_outStream_payload;
  wire                streamFifo_4_io_push_ready;
  wire                streamFifo_4_io_pop_valid;
  wire       [63:0]   streamFifo_4_io_pop_payload;
  wire       [4:0]    streamFifo_4_io_occupancy;
  wire       [4:0]    streamFifo_4_io_availability;
  wire                axisDataConverter_12_inStream_ready;
  wire                axisDataConverter_12_outStream_valid;
  wire       [7:0]    axisDataConverter_12_outStream_payload;
  wire                streamFifo_5_io_push_ready;
  wire                streamFifo_5_io_pop_valid;
  wire       [63:0]   streamFifo_5_io_pop_payload;
  wire       [4:0]    streamFifo_5_io_occupancy;
  wire       [4:0]    streamFifo_5_io_availability;
  wire                axisDataConverter_13_inStream_ready;
  wire                axisDataConverter_13_outStream_valid;
  wire       [7:0]    axisDataConverter_13_outStream_payload;
  wire                streamFifo_6_io_push_ready;
  wire                streamFifo_6_io_pop_valid;
  wire       [63:0]   streamFifo_6_io_pop_payload;
  wire       [4:0]    streamFifo_6_io_occupancy;
  wire       [4:0]    streamFifo_6_io_availability;
  wire                axisDataConverter_14_inStream_ready;
  wire                axisDataConverter_14_outStream_valid;
  wire       [7:0]    axisDataConverter_14_outStream_payload;
  wire                streamFifo_7_io_push_ready;
  wire                streamFifo_7_io_pop_valid;
  wire       [63:0]   streamFifo_7_io_pop_payload;
  wire       [4:0]    streamFifo_7_io_occupancy;
  wire       [4:0]    streamFifo_7_io_availability;
  wire                axisDataConverter_15_inStream_ready;
  wire                axisDataConverter_15_outStream_valid;
  wire       [7:0]    axisDataConverter_15_outStream_payload;
  reg        [7:0]    OutData_Switch;
  reg                 Switch_Reset;
  wire                TestValid_Signal_0;
  wire                TestValid_Signal_1;
  wire                TestValid_Signal_2;
  wire                TestValid_Signal_3;
  wire                TestValid_Signal_4;
  wire                TestValid_Signal_5;
  wire                TestValid_Signal_6;
  wire                TestValid_Signal_7;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_8_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_8_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_9_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_9_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_10_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_10_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_11_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_11_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_12_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_12_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_13_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_13_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_14_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_14_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_15_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_15_outStream_valid_regNext;
  reg                 SubModule_Img2Col_SubModule_LayerEnd_delay_1;
  reg                 SubModule_Img2Col_SubModule_LayerEnd_delay_2;
  reg                 SubModule_Img2Col_SubModule_LayerEnd_delay_3;

  Img2Col_Top SubModule (
    .start                          (start                               ), //i
    .sData_valid                    (s_axis_s2mm_tvalid                  ), //i
    .sData_ready                    (SubModule_sData_ready               ), //o
    .sData_payload                  (s_axis_s2mm_tdata[63:0]             ), //i
    .mData                          (SubModule_mData[63:0]               ), //o
    .mReady                         (streamFifo_io_push_ready            ), //i
    .mValid                         (SubModule_mValid                    ), //o
    .Fifo_Clear                     (SubModule_Fifo_Clear                ), //i
    .mLast                          (SubModule_mLast                     ), //o
    .Stride                         (Stride[4:0]                         ), //i
    .Kernel_Size                    (Kernel_Size[4:0]                    ), //i
    .Window_Size                    (Window_Size[15:0]                   ), //i
    .InFeature_Size                 (InFeature_Size[15:0]                ), //i
    .InFeature_Channel              (InFeature_Channel[15:0]             ), //i
    .OutFeature_Channel             (OutFeature_Channel[15:0]            ), //i
    .OutFeature_Size                (OutFeature_Size[15:0]               ), //i
    .OutCol_Count_Times             (OutCol_Count_Times[15:0]            ), //i
    .InCol_Count_Times              (InCol_Count_Times[15:0]             ), //i
    .OutRow_Count_Times             (OutRow_Count_Times[15:0]            ), //i
    .OutFeature_Channel_Count_Times (OutFeature_Channel_Count_Times[15:0]), //i
    .Sliding_Size                   (Sliding_Size[12:0]                  ), //i
    .Test_Signal                    (SubModule_Test_Signal               ), //o
    .Test_Generate_Period           (SubModule_Test_Generate_Period[15:0]), //i
    .Test_End                       (SubModule_Test_End                  ), //o
    .Raddr_Valid                    (SubModule_Raddr_Valid               ), //o
    .LayerEnd                       (SubModule_LayerEnd                  ), //o
    .SA_Row_Cnt_Valid               (SubModule_SA_Row_Cnt_Valid          ), //o
    .clk                            (clk                                 ), //i
    .reset                          (reset                               )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo (
    .io_push_valid   (streamFifo_io_push_valid          ), //i
    .io_push_ready   (streamFifo_io_push_ready          ), //o
    .io_push_payload (SubModule_mData[63:0]             ), //i
    .io_pop_valid    (streamFifo_io_pop_valid           ), //o
    .io_pop_ready    (axisDataConverter_8_inStream_ready), //i
    .io_pop_payload  (streamFifo_io_pop_payload[63:0]   ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (streamFifo_io_occupancy[4:0]      ), //o
    .io_availability (streamFifo_io_availability[4:0]   ), //o
    .clk             (clk                               ), //i
    .reset           (reset                             )  //i
  );
  AxisDataConverter axisDataConverter_8 (
    .inStream_valid    (streamFifo_io_pop_valid                   ), //i
    .inStream_ready    (axisDataConverter_8_inStream_ready        ), //o
    .inStream_payload  (streamFifo_io_pop_payload[63:0]           ), //i
    .outStream_valid   (axisDataConverter_8_outStream_valid       ), //o
    .outStream_ready   (1'b1                                      ), //i
    .outStream_payload (axisDataConverter_8_outStream_payload[7:0]), //o
    .clk               (clk                                       ), //i
    .reset             (reset                                     )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_1 (
    .io_push_valid   (streamFifo_1_io_push_valid        ), //i
    .io_push_ready   (streamFifo_1_io_push_ready        ), //o
    .io_push_payload (SubModule_mData[63:0]             ), //i
    .io_pop_valid    (streamFifo_1_io_pop_valid         ), //o
    .io_pop_ready    (axisDataConverter_9_inStream_ready), //i
    .io_pop_payload  (streamFifo_1_io_pop_payload[63:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (streamFifo_1_io_occupancy[4:0]    ), //o
    .io_availability (streamFifo_1_io_availability[4:0] ), //o
    .clk             (clk                               ), //i
    .reset           (reset                             )  //i
  );
  AxisDataConverter axisDataConverter_9 (
    .inStream_valid    (streamFifo_1_io_pop_valid                 ), //i
    .inStream_ready    (axisDataConverter_9_inStream_ready        ), //o
    .inStream_payload  (streamFifo_1_io_pop_payload[63:0]         ), //i
    .outStream_valid   (axisDataConverter_9_outStream_valid       ), //o
    .outStream_ready   (1'b1                                      ), //i
    .outStream_payload (axisDataConverter_9_outStream_payload[7:0]), //o
    .clk               (clk                                       ), //i
    .reset             (reset                                     )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_2 (
    .io_push_valid   (streamFifo_2_io_push_valid         ), //i
    .io_push_ready   (streamFifo_2_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_2_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_10_inStream_ready), //i
    .io_pop_payload  (streamFifo_2_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_2_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_2_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_10 (
    .inStream_valid    (streamFifo_2_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_10_inStream_ready        ), //o
    .inStream_payload  (streamFifo_2_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_10_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_10_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_3 (
    .io_push_valid   (streamFifo_3_io_push_valid         ), //i
    .io_push_ready   (streamFifo_3_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_3_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_11_inStream_ready), //i
    .io_pop_payload  (streamFifo_3_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_3_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_3_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_11 (
    .inStream_valid    (streamFifo_3_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_11_inStream_ready        ), //o
    .inStream_payload  (streamFifo_3_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_11_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_11_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_4 (
    .io_push_valid   (streamFifo_4_io_push_valid         ), //i
    .io_push_ready   (streamFifo_4_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_4_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_12_inStream_ready), //i
    .io_pop_payload  (streamFifo_4_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_4_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_4_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_12 (
    .inStream_valid    (streamFifo_4_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_12_inStream_ready        ), //o
    .inStream_payload  (streamFifo_4_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_12_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_12_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_5 (
    .io_push_valid   (streamFifo_5_io_push_valid         ), //i
    .io_push_ready   (streamFifo_5_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_5_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_13_inStream_ready), //i
    .io_pop_payload  (streamFifo_5_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_5_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_5_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_13 (
    .inStream_valid    (streamFifo_5_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_13_inStream_ready        ), //o
    .inStream_payload  (streamFifo_5_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_13_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_13_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_6 (
    .io_push_valid   (streamFifo_6_io_push_valid         ), //i
    .io_push_ready   (streamFifo_6_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_6_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_14_inStream_ready), //i
    .io_pop_payload  (streamFifo_6_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_6_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_6_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_14 (
    .inStream_valid    (streamFifo_6_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_14_inStream_ready        ), //o
    .inStream_payload  (streamFifo_6_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_14_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_14_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_7 (
    .io_push_valid   (streamFifo_7_io_push_valid         ), //i
    .io_push_ready   (streamFifo_7_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_7_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_15_inStream_ready), //i
    .io_pop_payload  (streamFifo_7_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_7_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_7_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_15 (
    .inStream_valid    (streamFifo_7_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_15_inStream_ready        ), //o
    .inStream_payload  (streamFifo_7_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_15_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_15_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  assign streamFifo_io_push_valid = (OutData_Switch[0] && SubModule_mValid);
  always @(*) begin
    mData[7 : 0] = SubModule_Img2Col_axisDataConverter_8_outStream_payload_regNext;
    mData[15 : 8] = SubModule_Img2Col_axisDataConverter_9_outStream_payload_regNext;
    mData[23 : 16] = SubModule_Img2Col_axisDataConverter_10_outStream_payload_regNext;
    mData[31 : 24] = SubModule_Img2Col_axisDataConverter_11_outStream_payload_regNext;
    mData[39 : 32] = SubModule_Img2Col_axisDataConverter_12_outStream_payload_regNext;
    mData[47 : 40] = SubModule_Img2Col_axisDataConverter_13_outStream_payload_regNext;
    mData[55 : 48] = SubModule_Img2Col_axisDataConverter_14_outStream_payload_regNext;
    mData[63 : 56] = SubModule_Img2Col_axisDataConverter_15_outStream_payload_regNext;
  end

  always @(*) begin
    mValid[0] = SubModule_Img2Col_axisDataConverter_8_outStream_valid_regNext;
    mValid[1] = SubModule_Img2Col_axisDataConverter_9_outStream_valid_regNext;
    mValid[2] = SubModule_Img2Col_axisDataConverter_10_outStream_valid_regNext;
    mValid[3] = SubModule_Img2Col_axisDataConverter_11_outStream_valid_regNext;
    mValid[4] = SubModule_Img2Col_axisDataConverter_12_outStream_valid_regNext;
    mValid[5] = SubModule_Img2Col_axisDataConverter_13_outStream_valid_regNext;
    mValid[6] = SubModule_Img2Col_axisDataConverter_14_outStream_valid_regNext;
    mValid[7] = SubModule_Img2Col_axisDataConverter_15_outStream_valid_regNext;
  end

  assign streamFifo_1_io_push_valid = (OutData_Switch[1] && SubModule_mValid);
  assign streamFifo_2_io_push_valid = (OutData_Switch[2] && SubModule_mValid);
  assign streamFifo_3_io_push_valid = (OutData_Switch[3] && SubModule_mValid);
  assign streamFifo_4_io_push_valid = (OutData_Switch[4] && SubModule_mValid);
  assign streamFifo_5_io_push_valid = (OutData_Switch[5] && SubModule_mValid);
  assign streamFifo_6_io_push_valid = (OutData_Switch[6] && SubModule_mValid);
  assign streamFifo_7_io_push_valid = (OutData_Switch[7] && SubModule_mValid);
  assign Raddr_Valid = axisDataConverter_8_outStream_valid;
  assign s_axis_s2mm_tready = SubModule_sData_ready;
  assign SubModule_Fifo_Clear = (! streamFifo_io_pop_valid);
  assign LayerEnd = SubModule_Img2Col_SubModule_LayerEnd_delay_3;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      OutData_Switch <= 8'h01;
    end else begin
      if(Switch_Reset) begin
        OutData_Switch <= 8'h01;
      end else begin
        if(SubModule_mValid) begin
          OutData_Switch <= {OutData_Switch[6 : 0],OutData_Switch[7 : 7]};
        end
      end
    end
  end

  always @(posedge clk) begin
    Switch_Reset <= SubModule_SA_Row_Cnt_Valid;
    SubModule_Img2Col_axisDataConverter_8_outStream_payload_regNext <= axisDataConverter_8_outStream_payload;
    SubModule_Img2Col_axisDataConverter_8_outStream_valid_regNext <= axisDataConverter_8_outStream_valid;
    SubModule_Img2Col_axisDataConverter_9_outStream_payload_regNext <= axisDataConverter_9_outStream_payload;
    SubModule_Img2Col_axisDataConverter_9_outStream_valid_regNext <= axisDataConverter_9_outStream_valid;
    SubModule_Img2Col_axisDataConverter_10_outStream_payload_regNext <= axisDataConverter_10_outStream_payload;
    SubModule_Img2Col_axisDataConverter_10_outStream_valid_regNext <= axisDataConverter_10_outStream_valid;
    SubModule_Img2Col_axisDataConverter_11_outStream_payload_regNext <= axisDataConverter_11_outStream_payload;
    SubModule_Img2Col_axisDataConverter_11_outStream_valid_regNext <= axisDataConverter_11_outStream_valid;
    SubModule_Img2Col_axisDataConverter_12_outStream_payload_regNext <= axisDataConverter_12_outStream_payload;
    SubModule_Img2Col_axisDataConverter_12_outStream_valid_regNext <= axisDataConverter_12_outStream_valid;
    SubModule_Img2Col_axisDataConverter_13_outStream_payload_regNext <= axisDataConverter_13_outStream_payload;
    SubModule_Img2Col_axisDataConverter_13_outStream_valid_regNext <= axisDataConverter_13_outStream_valid;
    SubModule_Img2Col_axisDataConverter_14_outStream_payload_regNext <= axisDataConverter_14_outStream_payload;
    SubModule_Img2Col_axisDataConverter_14_outStream_valid_regNext <= axisDataConverter_14_outStream_valid;
    SubModule_Img2Col_axisDataConverter_15_outStream_payload_regNext <= axisDataConverter_15_outStream_payload;
    SubModule_Img2Col_axisDataConverter_15_outStream_valid_regNext <= axisDataConverter_15_outStream_valid;
    SubModule_Img2Col_SubModule_LayerEnd_delay_1 <= SubModule_LayerEnd;
    SubModule_Img2Col_SubModule_LayerEnd_delay_2 <= SubModule_Img2Col_SubModule_LayerEnd_delay_1;
    SubModule_Img2Col_SubModule_LayerEnd_delay_3 <= SubModule_Img2Col_SubModule_LayerEnd_delay_2;
  end


endmodule

module Compute_DataIn_Switch (
  input      [1:0]    Switch,
  input      [63:0]   s0_axis_s2mm_tdata,
  input      [7:0]    s0_axis_s2mm_tkeep,
  input               s0_axis_s2mm_tlast,
  output reg          s0_axis_s2mm_tready,
  input               s0_axis_s2mm_tvalid,
  output reg [63:0]   m_0_axis_mm2s_tdata,
  output     [7:0]    m_0_axis_mm2s_tkeep,
  output reg          m_0_axis_mm2s_tlast,
  input               m_0_axis_mm2s_tready,
  output reg          m_0_axis_mm2s_tvalid,
  output reg [63:0]   m_1_axis_mm2s_tdata,
  output     [7:0]    m_1_axis_mm2s_tkeep,
  output reg          m_1_axis_mm2s_tlast,
  input               m_1_axis_mm2s_tready,
  output reg          m_1_axis_mm2s_tvalid
);

  wire                when_Axis_Switch_l103;
  wire                when_Axis_Switch_l103_1;

  assign m_0_axis_mm2s_tkeep = s0_axis_s2mm_tkeep;
  assign m_1_axis_mm2s_tkeep = s0_axis_s2mm_tkeep;
  always @(*) begin
    s0_axis_s2mm_tready = 1'b0;
    if(when_Axis_Switch_l103) begin
      s0_axis_s2mm_tready = m_0_axis_mm2s_tready;
    end
    if(when_Axis_Switch_l103_1) begin
      s0_axis_s2mm_tready = m_1_axis_mm2s_tready;
    end
  end

  assign when_Axis_Switch_l103 = (Switch == 2'b00);
  always @(*) begin
    if(when_Axis_Switch_l103) begin
      m_0_axis_mm2s_tdata = s0_axis_s2mm_tdata;
    end else begin
      m_0_axis_mm2s_tdata = 64'h0;
    end
  end

  always @(*) begin
    if(when_Axis_Switch_l103) begin
      m_0_axis_mm2s_tlast = s0_axis_s2mm_tlast;
    end else begin
      m_0_axis_mm2s_tlast = 1'b0;
    end
  end

  always @(*) begin
    if(when_Axis_Switch_l103) begin
      m_0_axis_mm2s_tvalid = s0_axis_s2mm_tvalid;
    end else begin
      m_0_axis_mm2s_tvalid = 1'b0;
    end
  end

  assign when_Axis_Switch_l103_1 = (Switch == 2'b01);
  always @(*) begin
    if(when_Axis_Switch_l103_1) begin
      m_1_axis_mm2s_tdata = s0_axis_s2mm_tdata;
    end else begin
      m_1_axis_mm2s_tdata = 64'h0;
    end
  end

  always @(*) begin
    if(when_Axis_Switch_l103_1) begin
      m_1_axis_mm2s_tlast = s0_axis_s2mm_tlast;
    end else begin
      m_1_axis_mm2s_tlast = 1'b0;
    end
  end

  always @(*) begin
    if(when_Axis_Switch_l103_1) begin
      m_1_axis_mm2s_tvalid = s0_axis_s2mm_tvalid;
    end else begin
      m_1_axis_mm2s_tvalid = 1'b0;
    end
  end


endmodule

module Weight_Cache (
  input               start,
  input               sData_valid,
  output              sData_ready,
  input      [63:0]   sData_payload,
  input      [15:0]   Matrix_Row,
  input      [15:0]   Matrix_Col,
  output     [7:0]    mData_0,
  output     [7:0]    mData_1,
  output     [7:0]    mData_2,
  output     [7:0]    mData_3,
  output     [7:0]    mData_4,
  output     [7:0]    mData_5,
  output     [7:0]    mData_6,
  output     [7:0]    mData_7,
  output     [7:0]    mData_8,
  output     [7:0]    mData_9,
  output     [7:0]    mData_10,
  output     [7:0]    mData_11,
  output     [7:0]    mData_12,
  output     [7:0]    mData_13,
  output     [7:0]    mData_14,
  output     [7:0]    mData_15,
  output     [7:0]    mData_16,
  output     [7:0]    mData_17,
  output     [7:0]    mData_18,
  output     [7:0]    mData_19,
  output     [7:0]    mData_20,
  output     [7:0]    mData_21,
  output     [7:0]    mData_22,
  output     [7:0]    mData_23,
  output     [7:0]    mData_24,
  output     [7:0]    mData_25,
  output     [7:0]    mData_26,
  output     [7:0]    mData_27,
  output     [7:0]    mData_28,
  output     [7:0]    mData_29,
  output     [7:0]    mData_30,
  output     [7:0]    mData_31,
  output     [7:0]    mData_32,
  output     [7:0]    mData_33,
  output     [7:0]    mData_34,
  output     [7:0]    mData_35,
  output     [7:0]    mData_36,
  output     [7:0]    mData_37,
  output     [7:0]    mData_38,
  output     [7:0]    mData_39,
  output     [7:0]    mData_40,
  output     [7:0]    mData_41,
  output     [7:0]    mData_42,
  output     [7:0]    mData_43,
  output     [7:0]    mData_44,
  output     [7:0]    mData_45,
  output     [7:0]    mData_46,
  output     [7:0]    mData_47,
  output     [7:0]    mData_48,
  output     [7:0]    mData_49,
  output     [7:0]    mData_50,
  output     [7:0]    mData_51,
  output     [7:0]    mData_52,
  output     [7:0]    mData_53,
  output     [7:0]    mData_54,
  output     [7:0]    mData_55,
  output     [7:0]    mData_56,
  output     [7:0]    mData_57,
  output     [7:0]    mData_58,
  output     [7:0]    mData_59,
  output     [7:0]    mData_60,
  output     [7:0]    mData_61,
  output     [7:0]    mData_62,
  output     [7:0]    mData_63,
  input               Raddr_Valid,
  output              Weight_Cached,
  input               LayerEnd,
  output     [63:0]   MatrixCol_Switch,
  input               clk,
  input               reset
);
  localparam WEIGHT_CACHE_STATUS_IDLE = 4'd1;
  localparam WEIGHT_CACHE_STATUS_INIT = 4'd2;
  localparam WEIGHT_CACHE_STATUS_CACHE_WEIGHT = 4'd4;
  localparam WEIGHT_CACHE_STATUS_SA_COMPUTE = 4'd8;

  wire       [10:0]   xil_SimpleDualBram_addra;
  wire                xil_SimpleDualBram_ena;
  wire       [13:0]   xil_SimpleDualBram_addrb;
  wire       [10:0]   xil_SimpleDualBram_1_addra;
  wire                xil_SimpleDualBram_1_ena;
  wire       [13:0]   xil_SimpleDualBram_1_addrb;
  wire       [10:0]   xil_SimpleDualBram_2_addra;
  wire                xil_SimpleDualBram_2_ena;
  wire       [13:0]   xil_SimpleDualBram_2_addrb;
  wire       [10:0]   xil_SimpleDualBram_3_addra;
  wire                xil_SimpleDualBram_3_ena;
  wire       [13:0]   xil_SimpleDualBram_3_addrb;
  wire       [10:0]   xil_SimpleDualBram_4_addra;
  wire                xil_SimpleDualBram_4_ena;
  wire       [13:0]   xil_SimpleDualBram_4_addrb;
  wire       [10:0]   xil_SimpleDualBram_5_addra;
  wire                xil_SimpleDualBram_5_ena;
  wire       [13:0]   xil_SimpleDualBram_5_addrb;
  wire       [10:0]   xil_SimpleDualBram_6_addra;
  wire                xil_SimpleDualBram_6_ena;
  wire       [13:0]   xil_SimpleDualBram_6_addrb;
  wire       [10:0]   xil_SimpleDualBram_7_addra;
  wire                xil_SimpleDualBram_7_ena;
  wire       [13:0]   xil_SimpleDualBram_7_addrb;
  wire       [10:0]   xil_SimpleDualBram_8_addra;
  wire                xil_SimpleDualBram_8_ena;
  wire       [13:0]   xil_SimpleDualBram_8_addrb;
  wire       [10:0]   xil_SimpleDualBram_9_addra;
  wire                xil_SimpleDualBram_9_ena;
  wire       [13:0]   xil_SimpleDualBram_9_addrb;
  wire       [10:0]   xil_SimpleDualBram_10_addra;
  wire                xil_SimpleDualBram_10_ena;
  wire       [13:0]   xil_SimpleDualBram_10_addrb;
  wire       [10:0]   xil_SimpleDualBram_11_addra;
  wire                xil_SimpleDualBram_11_ena;
  wire       [13:0]   xil_SimpleDualBram_11_addrb;
  wire       [10:0]   xil_SimpleDualBram_12_addra;
  wire                xil_SimpleDualBram_12_ena;
  wire       [13:0]   xil_SimpleDualBram_12_addrb;
  wire       [10:0]   xil_SimpleDualBram_13_addra;
  wire                xil_SimpleDualBram_13_ena;
  wire       [13:0]   xil_SimpleDualBram_13_addrb;
  wire       [10:0]   xil_SimpleDualBram_14_addra;
  wire                xil_SimpleDualBram_14_ena;
  wire       [13:0]   xil_SimpleDualBram_14_addrb;
  wire       [10:0]   xil_SimpleDualBram_15_addra;
  wire                xil_SimpleDualBram_15_ena;
  wire       [13:0]   xil_SimpleDualBram_15_addrb;
  wire       [10:0]   xil_SimpleDualBram_16_addra;
  wire                xil_SimpleDualBram_16_ena;
  wire       [13:0]   xil_SimpleDualBram_16_addrb;
  wire       [10:0]   xil_SimpleDualBram_17_addra;
  wire                xil_SimpleDualBram_17_ena;
  wire       [13:0]   xil_SimpleDualBram_17_addrb;
  wire       [10:0]   xil_SimpleDualBram_18_addra;
  wire                xil_SimpleDualBram_18_ena;
  wire       [13:0]   xil_SimpleDualBram_18_addrb;
  wire       [10:0]   xil_SimpleDualBram_19_addra;
  wire                xil_SimpleDualBram_19_ena;
  wire       [13:0]   xil_SimpleDualBram_19_addrb;
  wire       [10:0]   xil_SimpleDualBram_20_addra;
  wire                xil_SimpleDualBram_20_ena;
  wire       [13:0]   xil_SimpleDualBram_20_addrb;
  wire       [10:0]   xil_SimpleDualBram_21_addra;
  wire                xil_SimpleDualBram_21_ena;
  wire       [13:0]   xil_SimpleDualBram_21_addrb;
  wire       [10:0]   xil_SimpleDualBram_22_addra;
  wire                xil_SimpleDualBram_22_ena;
  wire       [13:0]   xil_SimpleDualBram_22_addrb;
  wire       [10:0]   xil_SimpleDualBram_23_addra;
  wire                xil_SimpleDualBram_23_ena;
  wire       [13:0]   xil_SimpleDualBram_23_addrb;
  wire       [10:0]   xil_SimpleDualBram_24_addra;
  wire                xil_SimpleDualBram_24_ena;
  wire       [13:0]   xil_SimpleDualBram_24_addrb;
  wire       [10:0]   xil_SimpleDualBram_25_addra;
  wire                xil_SimpleDualBram_25_ena;
  wire       [13:0]   xil_SimpleDualBram_25_addrb;
  wire       [10:0]   xil_SimpleDualBram_26_addra;
  wire                xil_SimpleDualBram_26_ena;
  wire       [13:0]   xil_SimpleDualBram_26_addrb;
  wire       [10:0]   xil_SimpleDualBram_27_addra;
  wire                xil_SimpleDualBram_27_ena;
  wire       [13:0]   xil_SimpleDualBram_27_addrb;
  wire       [10:0]   xil_SimpleDualBram_28_addra;
  wire                xil_SimpleDualBram_28_ena;
  wire       [13:0]   xil_SimpleDualBram_28_addrb;
  wire       [10:0]   xil_SimpleDualBram_29_addra;
  wire                xil_SimpleDualBram_29_ena;
  wire       [13:0]   xil_SimpleDualBram_29_addrb;
  wire       [10:0]   xil_SimpleDualBram_30_addra;
  wire                xil_SimpleDualBram_30_ena;
  wire       [13:0]   xil_SimpleDualBram_30_addrb;
  wire       [10:0]   xil_SimpleDualBram_31_addra;
  wire                xil_SimpleDualBram_31_ena;
  wire       [13:0]   xil_SimpleDualBram_31_addrb;
  wire       [10:0]   xil_SimpleDualBram_32_addra;
  wire                xil_SimpleDualBram_32_ena;
  wire       [13:0]   xil_SimpleDualBram_32_addrb;
  wire       [10:0]   xil_SimpleDualBram_33_addra;
  wire                xil_SimpleDualBram_33_ena;
  wire       [13:0]   xil_SimpleDualBram_33_addrb;
  wire       [10:0]   xil_SimpleDualBram_34_addra;
  wire                xil_SimpleDualBram_34_ena;
  wire       [13:0]   xil_SimpleDualBram_34_addrb;
  wire       [10:0]   xil_SimpleDualBram_35_addra;
  wire                xil_SimpleDualBram_35_ena;
  wire       [13:0]   xil_SimpleDualBram_35_addrb;
  wire       [10:0]   xil_SimpleDualBram_36_addra;
  wire                xil_SimpleDualBram_36_ena;
  wire       [13:0]   xil_SimpleDualBram_36_addrb;
  wire       [10:0]   xil_SimpleDualBram_37_addra;
  wire                xil_SimpleDualBram_37_ena;
  wire       [13:0]   xil_SimpleDualBram_37_addrb;
  wire       [10:0]   xil_SimpleDualBram_38_addra;
  wire                xil_SimpleDualBram_38_ena;
  wire       [13:0]   xil_SimpleDualBram_38_addrb;
  wire       [10:0]   xil_SimpleDualBram_39_addra;
  wire                xil_SimpleDualBram_39_ena;
  wire       [13:0]   xil_SimpleDualBram_39_addrb;
  wire       [10:0]   xil_SimpleDualBram_40_addra;
  wire                xil_SimpleDualBram_40_ena;
  wire       [13:0]   xil_SimpleDualBram_40_addrb;
  wire       [10:0]   xil_SimpleDualBram_41_addra;
  wire                xil_SimpleDualBram_41_ena;
  wire       [13:0]   xil_SimpleDualBram_41_addrb;
  wire       [10:0]   xil_SimpleDualBram_42_addra;
  wire                xil_SimpleDualBram_42_ena;
  wire       [13:0]   xil_SimpleDualBram_42_addrb;
  wire       [10:0]   xil_SimpleDualBram_43_addra;
  wire                xil_SimpleDualBram_43_ena;
  wire       [13:0]   xil_SimpleDualBram_43_addrb;
  wire       [10:0]   xil_SimpleDualBram_44_addra;
  wire                xil_SimpleDualBram_44_ena;
  wire       [13:0]   xil_SimpleDualBram_44_addrb;
  wire       [10:0]   xil_SimpleDualBram_45_addra;
  wire                xil_SimpleDualBram_45_ena;
  wire       [13:0]   xil_SimpleDualBram_45_addrb;
  wire       [10:0]   xil_SimpleDualBram_46_addra;
  wire                xil_SimpleDualBram_46_ena;
  wire       [13:0]   xil_SimpleDualBram_46_addrb;
  wire       [10:0]   xil_SimpleDualBram_47_addra;
  wire                xil_SimpleDualBram_47_ena;
  wire       [13:0]   xil_SimpleDualBram_47_addrb;
  wire       [10:0]   xil_SimpleDualBram_48_addra;
  wire                xil_SimpleDualBram_48_ena;
  wire       [13:0]   xil_SimpleDualBram_48_addrb;
  wire       [10:0]   xil_SimpleDualBram_49_addra;
  wire                xil_SimpleDualBram_49_ena;
  wire       [13:0]   xil_SimpleDualBram_49_addrb;
  wire       [10:0]   xil_SimpleDualBram_50_addra;
  wire                xil_SimpleDualBram_50_ena;
  wire       [13:0]   xil_SimpleDualBram_50_addrb;
  wire       [10:0]   xil_SimpleDualBram_51_addra;
  wire                xil_SimpleDualBram_51_ena;
  wire       [13:0]   xil_SimpleDualBram_51_addrb;
  wire       [10:0]   xil_SimpleDualBram_52_addra;
  wire                xil_SimpleDualBram_52_ena;
  wire       [13:0]   xil_SimpleDualBram_52_addrb;
  wire       [10:0]   xil_SimpleDualBram_53_addra;
  wire                xil_SimpleDualBram_53_ena;
  wire       [13:0]   xil_SimpleDualBram_53_addrb;
  wire       [10:0]   xil_SimpleDualBram_54_addra;
  wire                xil_SimpleDualBram_54_ena;
  wire       [13:0]   xil_SimpleDualBram_54_addrb;
  wire       [10:0]   xil_SimpleDualBram_55_addra;
  wire                xil_SimpleDualBram_55_ena;
  wire       [13:0]   xil_SimpleDualBram_55_addrb;
  wire       [10:0]   xil_SimpleDualBram_56_addra;
  wire                xil_SimpleDualBram_56_ena;
  wire       [13:0]   xil_SimpleDualBram_56_addrb;
  wire       [10:0]   xil_SimpleDualBram_57_addra;
  wire                xil_SimpleDualBram_57_ena;
  wire       [13:0]   xil_SimpleDualBram_57_addrb;
  wire       [10:0]   xil_SimpleDualBram_58_addra;
  wire                xil_SimpleDualBram_58_ena;
  wire       [13:0]   xil_SimpleDualBram_58_addrb;
  wire       [10:0]   xil_SimpleDualBram_59_addra;
  wire                xil_SimpleDualBram_59_ena;
  wire       [13:0]   xil_SimpleDualBram_59_addrb;
  wire       [10:0]   xil_SimpleDualBram_60_addra;
  wire                xil_SimpleDualBram_60_ena;
  wire       [13:0]   xil_SimpleDualBram_60_addrb;
  wire       [10:0]   xil_SimpleDualBram_61_addra;
  wire                xil_SimpleDualBram_61_ena;
  wire       [13:0]   xil_SimpleDualBram_61_addrb;
  wire       [10:0]   xil_SimpleDualBram_62_addra;
  wire                xil_SimpleDualBram_62_ena;
  wire       [13:0]   xil_SimpleDualBram_62_addrb;
  wire       [10:0]   xil_SimpleDualBram_63_addra;
  wire                xil_SimpleDualBram_63_ena;
  wire       [13:0]   xil_SimpleDualBram_63_addrb;
  wire       [7:0]    xil_SimpleDualBram_doutb;
  wire       [7:0]    xil_SimpleDualBram_1_doutb;
  wire       [7:0]    xil_SimpleDualBram_2_doutb;
  wire       [7:0]    xil_SimpleDualBram_3_doutb;
  wire       [7:0]    xil_SimpleDualBram_4_doutb;
  wire       [7:0]    xil_SimpleDualBram_5_doutb;
  wire       [7:0]    xil_SimpleDualBram_6_doutb;
  wire       [7:0]    xil_SimpleDualBram_7_doutb;
  wire       [7:0]    xil_SimpleDualBram_8_doutb;
  wire       [7:0]    xil_SimpleDualBram_9_doutb;
  wire       [7:0]    xil_SimpleDualBram_10_doutb;
  wire       [7:0]    xil_SimpleDualBram_11_doutb;
  wire       [7:0]    xil_SimpleDualBram_12_doutb;
  wire       [7:0]    xil_SimpleDualBram_13_doutb;
  wire       [7:0]    xil_SimpleDualBram_14_doutb;
  wire       [7:0]    xil_SimpleDualBram_15_doutb;
  wire       [7:0]    xil_SimpleDualBram_16_doutb;
  wire       [7:0]    xil_SimpleDualBram_17_doutb;
  wire       [7:0]    xil_SimpleDualBram_18_doutb;
  wire       [7:0]    xil_SimpleDualBram_19_doutb;
  wire       [7:0]    xil_SimpleDualBram_20_doutb;
  wire       [7:0]    xil_SimpleDualBram_21_doutb;
  wire       [7:0]    xil_SimpleDualBram_22_doutb;
  wire       [7:0]    xil_SimpleDualBram_23_doutb;
  wire       [7:0]    xil_SimpleDualBram_24_doutb;
  wire       [7:0]    xil_SimpleDualBram_25_doutb;
  wire       [7:0]    xil_SimpleDualBram_26_doutb;
  wire       [7:0]    xil_SimpleDualBram_27_doutb;
  wire       [7:0]    xil_SimpleDualBram_28_doutb;
  wire       [7:0]    xil_SimpleDualBram_29_doutb;
  wire       [7:0]    xil_SimpleDualBram_30_doutb;
  wire       [7:0]    xil_SimpleDualBram_31_doutb;
  wire       [7:0]    xil_SimpleDualBram_32_doutb;
  wire       [7:0]    xil_SimpleDualBram_33_doutb;
  wire       [7:0]    xil_SimpleDualBram_34_doutb;
  wire       [7:0]    xil_SimpleDualBram_35_doutb;
  wire       [7:0]    xil_SimpleDualBram_36_doutb;
  wire       [7:0]    xil_SimpleDualBram_37_doutb;
  wire       [7:0]    xil_SimpleDualBram_38_doutb;
  wire       [7:0]    xil_SimpleDualBram_39_doutb;
  wire       [7:0]    xil_SimpleDualBram_40_doutb;
  wire       [7:0]    xil_SimpleDualBram_41_doutb;
  wire       [7:0]    xil_SimpleDualBram_42_doutb;
  wire       [7:0]    xil_SimpleDualBram_43_doutb;
  wire       [7:0]    xil_SimpleDualBram_44_doutb;
  wire       [7:0]    xil_SimpleDualBram_45_doutb;
  wire       [7:0]    xil_SimpleDualBram_46_doutb;
  wire       [7:0]    xil_SimpleDualBram_47_doutb;
  wire       [7:0]    xil_SimpleDualBram_48_doutb;
  wire       [7:0]    xil_SimpleDualBram_49_doutb;
  wire       [7:0]    xil_SimpleDualBram_50_doutb;
  wire       [7:0]    xil_SimpleDualBram_51_doutb;
  wire       [7:0]    xil_SimpleDualBram_52_doutb;
  wire       [7:0]    xil_SimpleDualBram_53_doutb;
  wire       [7:0]    xil_SimpleDualBram_54_doutb;
  wire       [7:0]    xil_SimpleDualBram_55_doutb;
  wire       [7:0]    xil_SimpleDualBram_56_doutb;
  wire       [7:0]    xil_SimpleDualBram_57_doutb;
  wire       [7:0]    xil_SimpleDualBram_58_doutb;
  wire       [7:0]    xil_SimpleDualBram_59_doutb;
  wire       [7:0]    xil_SimpleDualBram_60_doutb;
  wire       [7:0]    xil_SimpleDualBram_61_doutb;
  wire       [7:0]    xil_SimpleDualBram_62_doutb;
  wire       [7:0]    xil_SimpleDualBram_63_doutb;
  wire       [15:0]   _zz_In_Row_Cnt_valid;
  wire       [12:0]   _zz_In_Row_Cnt_valid_1;
  wire       [15:0]   _zz_In_Col_Cnt_valid;
  wire       [15:0]   _zz_OutRow_Cnt_valid;
  wire       [15:0]   _zz_OutCol_Cnt_valid;
  wire       [15:0]   _zz_OutCol_Cnt_count_1;
  wire       [15:0]   _zz_Write_Row_Base_Addr;
  wire       [15:0]   _zz_addra;
  wire       [15:0]   _zz_addrb;
  wire       [0:0]    _zz_ena;
  wire       [15:0]   _zz_addra_1;
  wire       [15:0]   _zz_addrb_1;
  wire       [0:0]    _zz_ena_1;
  wire       [15:0]   _zz_addra_2;
  wire       [15:0]   _zz_addrb_2;
  wire       [0:0]    _zz_ena_2;
  wire       [15:0]   _zz_addra_3;
  wire       [15:0]   _zz_addrb_3;
  wire       [0:0]    _zz_ena_3;
  wire       [15:0]   _zz_addra_4;
  wire       [15:0]   _zz_addrb_4;
  wire       [0:0]    _zz_ena_4;
  wire       [15:0]   _zz_addra_5;
  wire       [15:0]   _zz_addrb_5;
  wire       [0:0]    _zz_ena_5;
  wire       [15:0]   _zz_addra_6;
  wire       [15:0]   _zz_addrb_6;
  wire       [0:0]    _zz_ena_6;
  wire       [15:0]   _zz_addra_7;
  wire       [15:0]   _zz_addrb_7;
  wire       [0:0]    _zz_ena_7;
  wire       [15:0]   _zz_addra_8;
  wire       [15:0]   _zz_addrb_8;
  wire       [0:0]    _zz_ena_8;
  wire       [15:0]   _zz_addra_9;
  wire       [15:0]   _zz_addrb_9;
  wire       [0:0]    _zz_ena_9;
  wire       [15:0]   _zz_addra_10;
  wire       [15:0]   _zz_addrb_10;
  wire       [0:0]    _zz_ena_10;
  wire       [15:0]   _zz_addra_11;
  wire       [15:0]   _zz_addrb_11;
  wire       [0:0]    _zz_ena_11;
  wire       [15:0]   _zz_addra_12;
  wire       [15:0]   _zz_addrb_12;
  wire       [0:0]    _zz_ena_12;
  wire       [15:0]   _zz_addra_13;
  wire       [15:0]   _zz_addrb_13;
  wire       [0:0]    _zz_ena_13;
  wire       [15:0]   _zz_addra_14;
  wire       [15:0]   _zz_addrb_14;
  wire       [0:0]    _zz_ena_14;
  wire       [15:0]   _zz_addra_15;
  wire       [15:0]   _zz_addrb_15;
  wire       [0:0]    _zz_ena_15;
  wire       [15:0]   _zz_addra_16;
  wire       [15:0]   _zz_addrb_16;
  wire       [0:0]    _zz_ena_16;
  wire       [15:0]   _zz_addra_17;
  wire       [15:0]   _zz_addrb_17;
  wire       [0:0]    _zz_ena_17;
  wire       [15:0]   _zz_addra_18;
  wire       [15:0]   _zz_addrb_18;
  wire       [0:0]    _zz_ena_18;
  wire       [15:0]   _zz_addra_19;
  wire       [15:0]   _zz_addrb_19;
  wire       [0:0]    _zz_ena_19;
  wire       [15:0]   _zz_addra_20;
  wire       [15:0]   _zz_addrb_20;
  wire       [0:0]    _zz_ena_20;
  wire       [15:0]   _zz_addra_21;
  wire       [15:0]   _zz_addrb_21;
  wire       [0:0]    _zz_ena_21;
  wire       [15:0]   _zz_addra_22;
  wire       [15:0]   _zz_addrb_22;
  wire       [0:0]    _zz_ena_22;
  wire       [15:0]   _zz_addra_23;
  wire       [15:0]   _zz_addrb_23;
  wire       [0:0]    _zz_ena_23;
  wire       [15:0]   _zz_addra_24;
  wire       [15:0]   _zz_addrb_24;
  wire       [0:0]    _zz_ena_24;
  wire       [15:0]   _zz_addra_25;
  wire       [15:0]   _zz_addrb_25;
  wire       [0:0]    _zz_ena_25;
  wire       [15:0]   _zz_addra_26;
  wire       [15:0]   _zz_addrb_26;
  wire       [0:0]    _zz_ena_26;
  wire       [15:0]   _zz_addra_27;
  wire       [15:0]   _zz_addrb_27;
  wire       [0:0]    _zz_ena_27;
  wire       [15:0]   _zz_addra_28;
  wire       [15:0]   _zz_addrb_28;
  wire       [0:0]    _zz_ena_28;
  wire       [15:0]   _zz_addra_29;
  wire       [15:0]   _zz_addrb_29;
  wire       [0:0]    _zz_ena_29;
  wire       [15:0]   _zz_addra_30;
  wire       [15:0]   _zz_addrb_30;
  wire       [0:0]    _zz_ena_30;
  wire       [15:0]   _zz_addra_31;
  wire       [15:0]   _zz_addrb_31;
  wire       [0:0]    _zz_ena_31;
  wire       [15:0]   _zz_addra_32;
  wire       [15:0]   _zz_addrb_32;
  wire       [0:0]    _zz_ena_32;
  wire       [15:0]   _zz_addra_33;
  wire       [15:0]   _zz_addrb_33;
  wire       [0:0]    _zz_ena_33;
  wire       [15:0]   _zz_addra_34;
  wire       [15:0]   _zz_addrb_34;
  wire       [0:0]    _zz_ena_34;
  wire       [15:0]   _zz_addra_35;
  wire       [15:0]   _zz_addrb_35;
  wire       [0:0]    _zz_ena_35;
  wire       [15:0]   _zz_addra_36;
  wire       [15:0]   _zz_addrb_36;
  wire       [0:0]    _zz_ena_36;
  wire       [15:0]   _zz_addra_37;
  wire       [15:0]   _zz_addrb_37;
  wire       [0:0]    _zz_ena_37;
  wire       [15:0]   _zz_addra_38;
  wire       [15:0]   _zz_addrb_38;
  wire       [0:0]    _zz_ena_38;
  wire       [15:0]   _zz_addra_39;
  wire       [15:0]   _zz_addrb_39;
  wire       [0:0]    _zz_ena_39;
  wire       [15:0]   _zz_addra_40;
  wire       [15:0]   _zz_addrb_40;
  wire       [0:0]    _zz_ena_40;
  wire       [15:0]   _zz_addra_41;
  wire       [15:0]   _zz_addrb_41;
  wire       [0:0]    _zz_ena_41;
  wire       [15:0]   _zz_addra_42;
  wire       [15:0]   _zz_addrb_42;
  wire       [0:0]    _zz_ena_42;
  wire       [15:0]   _zz_addra_43;
  wire       [15:0]   _zz_addrb_43;
  wire       [0:0]    _zz_ena_43;
  wire       [15:0]   _zz_addra_44;
  wire       [15:0]   _zz_addrb_44;
  wire       [0:0]    _zz_ena_44;
  wire       [15:0]   _zz_addra_45;
  wire       [15:0]   _zz_addrb_45;
  wire       [0:0]    _zz_ena_45;
  wire       [15:0]   _zz_addra_46;
  wire       [15:0]   _zz_addrb_46;
  wire       [0:0]    _zz_ena_46;
  wire       [15:0]   _zz_addra_47;
  wire       [15:0]   _zz_addrb_47;
  wire       [0:0]    _zz_ena_47;
  wire       [15:0]   _zz_addra_48;
  wire       [15:0]   _zz_addrb_48;
  wire       [0:0]    _zz_ena_48;
  wire       [15:0]   _zz_addra_49;
  wire       [15:0]   _zz_addrb_49;
  wire       [0:0]    _zz_ena_49;
  wire       [15:0]   _zz_addra_50;
  wire       [15:0]   _zz_addrb_50;
  wire       [0:0]    _zz_ena_50;
  wire       [15:0]   _zz_addra_51;
  wire       [15:0]   _zz_addrb_51;
  wire       [0:0]    _zz_ena_51;
  wire       [15:0]   _zz_addra_52;
  wire       [15:0]   _zz_addrb_52;
  wire       [0:0]    _zz_ena_52;
  wire       [15:0]   _zz_addra_53;
  wire       [15:0]   _zz_addrb_53;
  wire       [0:0]    _zz_ena_53;
  wire       [15:0]   _zz_addra_54;
  wire       [15:0]   _zz_addrb_54;
  wire       [0:0]    _zz_ena_54;
  wire       [15:0]   _zz_addra_55;
  wire       [15:0]   _zz_addrb_55;
  wire       [0:0]    _zz_ena_55;
  wire       [15:0]   _zz_addra_56;
  wire       [15:0]   _zz_addrb_56;
  wire       [0:0]    _zz_ena_56;
  wire       [15:0]   _zz_addra_57;
  wire       [15:0]   _zz_addrb_57;
  wire       [0:0]    _zz_ena_57;
  wire       [15:0]   _zz_addra_58;
  wire       [15:0]   _zz_addrb_58;
  wire       [0:0]    _zz_ena_58;
  wire       [15:0]   _zz_addra_59;
  wire       [15:0]   _zz_addrb_59;
  wire       [0:0]    _zz_ena_59;
  wire       [15:0]   _zz_addra_60;
  wire       [15:0]   _zz_addrb_60;
  wire       [0:0]    _zz_ena_60;
  wire       [15:0]   _zz_addra_61;
  wire       [15:0]   _zz_addrb_61;
  wire       [0:0]    _zz_ena_61;
  wire       [15:0]   _zz_addra_62;
  wire       [15:0]   _zz_addrb_62;
  wire       [0:0]    _zz_ena_62;
  wire       [15:0]   _zz_addra_63;
  wire       [15:0]   _zz_addrb_63;
  wire       [0:0]    _zz_ena_63;
  reg                 start_regNext;
  wire                when_SA3D_WeightCache_l33;
  reg        [3:0]    Fsm_currentState;
  reg        [3:0]    Fsm_nextState;
  wire                Fsm_Init_End;
  wire                Fsm_Weight_All_Cached;
  wire                Fsm_SA_Computed;
  wire                when_WaCounter_l19;
  reg        [2:0]    Init_Count_count;
  reg                 Init_Count_valid;
  wire                when_WaCounter_l14;
  reg        [63:0]   InData_Switch;
  wire       [12:0]   Matrix_In_MaxCnt;
  wire                sData_fire;
  reg        [15:0]   In_Row_Cnt_count;
  wire                In_Row_Cnt_valid;
  reg        [15:0]   In_Col_Cnt_count;
  wire                In_Col_Cnt_valid;
  reg        [15:0]   Read_Row_Base_Addr;
  reg        [15:0]   Write_Row_Base_Addr;
  wire                when_WaCounter_l40;
  reg        [15:0]   OutRow_Cnt_count;
  wire                OutRow_Cnt_valid;
  wire       [3:0]    _zz_OutCol_Cnt_count;
  reg        [15:0]   OutCol_Cnt_count;
  reg                 OutCol_Cnt_valid;
  reg        [5:0]    Col_In_8_Cnt_count;
  reg                 Col_In_8_Cnt_valid;
  wire                when_SA3D_WeightCache_l129;
  wire                when_SA3D_WeightCache_l134;
  wire                sData_fire_1;
  wire                sData_fire_2;
  wire                sData_fire_3;
  wire                sData_fire_4;
  wire                sData_fire_5;
  wire                sData_fire_6;
  wire                sData_fire_7;
  wire                sData_fire_8;
  wire                sData_fire_9;
  wire                sData_fire_10;
  wire                sData_fire_11;
  wire                sData_fire_12;
  wire                sData_fire_13;
  wire                sData_fire_14;
  wire                sData_fire_15;
  wire                sData_fire_16;
  wire                sData_fire_17;
  wire                sData_fire_18;
  wire                sData_fire_19;
  wire                sData_fire_20;
  wire                sData_fire_21;
  wire                sData_fire_22;
  wire                sData_fire_23;
  wire                sData_fire_24;
  wire                sData_fire_25;
  wire                sData_fire_26;
  wire                sData_fire_27;
  wire                sData_fire_28;
  wire                sData_fire_29;
  wire                sData_fire_30;
  wire                sData_fire_31;
  wire                sData_fire_32;
  wire                sData_fire_33;
  wire                sData_fire_34;
  wire                sData_fire_35;
  wire                sData_fire_36;
  wire                sData_fire_37;
  wire                sData_fire_38;
  wire                sData_fire_39;
  wire                sData_fire_40;
  wire                sData_fire_41;
  wire                sData_fire_42;
  wire                sData_fire_43;
  wire                sData_fire_44;
  wire                sData_fire_45;
  wire                sData_fire_46;
  wire                sData_fire_47;
  wire                sData_fire_48;
  wire                sData_fire_49;
  wire                sData_fire_50;
  wire                sData_fire_51;
  wire                sData_fire_52;
  wire                sData_fire_53;
  wire                sData_fire_54;
  wire                sData_fire_55;
  wire                sData_fire_56;
  wire                sData_fire_57;
  wire                sData_fire_58;
  wire                sData_fire_59;
  wire                sData_fire_60;
  wire                sData_fire_61;
  wire                sData_fire_62;
  wire                sData_fire_63;
  wire                sData_fire_64;
  reg        [63:0]   MatrixCol_Switch_1;
  reg        [63:0]   MatrixCol_Switch_1_regNext;
  `ifndef SYNTHESIS
  reg [95:0] Fsm_currentState_string;
  reg [95:0] Fsm_nextState_string;
  `endif


  assign _zz_In_Row_Cnt_valid_1 = (Matrix_In_MaxCnt - 13'h0001);
  assign _zz_In_Row_Cnt_valid = {3'd0, _zz_In_Row_Cnt_valid_1};
  assign _zz_In_Col_Cnt_valid = (Matrix_Col - 16'h0001);
  assign _zz_OutRow_Cnt_valid = (Matrix_Row - 16'h0001);
  assign _zz_OutCol_Cnt_valid = {12'd0, _zz_OutCol_Cnt_count};
  assign _zz_OutCol_Cnt_count_1 = {12'd0, _zz_OutCol_Cnt_count};
  assign _zz_Write_Row_Base_Addr = {3'd0, Matrix_In_MaxCnt};
  assign _zz_addra = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena = InData_Switch[0 : 0];
  assign _zz_addra_1 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_1 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_1 = InData_Switch[1 : 1];
  assign _zz_addra_2 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_2 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_2 = InData_Switch[2 : 2];
  assign _zz_addra_3 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_3 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_3 = InData_Switch[3 : 3];
  assign _zz_addra_4 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_4 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_4 = InData_Switch[4 : 4];
  assign _zz_addra_5 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_5 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_5 = InData_Switch[5 : 5];
  assign _zz_addra_6 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_6 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_6 = InData_Switch[6 : 6];
  assign _zz_addra_7 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_7 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_7 = InData_Switch[7 : 7];
  assign _zz_addra_8 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_8 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_8 = InData_Switch[8 : 8];
  assign _zz_addra_9 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_9 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_9 = InData_Switch[9 : 9];
  assign _zz_addra_10 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_10 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_10 = InData_Switch[10 : 10];
  assign _zz_addra_11 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_11 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_11 = InData_Switch[11 : 11];
  assign _zz_addra_12 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_12 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_12 = InData_Switch[12 : 12];
  assign _zz_addra_13 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_13 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_13 = InData_Switch[13 : 13];
  assign _zz_addra_14 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_14 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_14 = InData_Switch[14 : 14];
  assign _zz_addra_15 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_15 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_15 = InData_Switch[15 : 15];
  assign _zz_addra_16 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_16 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_16 = InData_Switch[16 : 16];
  assign _zz_addra_17 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_17 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_17 = InData_Switch[17 : 17];
  assign _zz_addra_18 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_18 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_18 = InData_Switch[18 : 18];
  assign _zz_addra_19 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_19 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_19 = InData_Switch[19 : 19];
  assign _zz_addra_20 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_20 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_20 = InData_Switch[20 : 20];
  assign _zz_addra_21 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_21 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_21 = InData_Switch[21 : 21];
  assign _zz_addra_22 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_22 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_22 = InData_Switch[22 : 22];
  assign _zz_addra_23 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_23 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_23 = InData_Switch[23 : 23];
  assign _zz_addra_24 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_24 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_24 = InData_Switch[24 : 24];
  assign _zz_addra_25 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_25 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_25 = InData_Switch[25 : 25];
  assign _zz_addra_26 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_26 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_26 = InData_Switch[26 : 26];
  assign _zz_addra_27 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_27 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_27 = InData_Switch[27 : 27];
  assign _zz_addra_28 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_28 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_28 = InData_Switch[28 : 28];
  assign _zz_addra_29 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_29 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_29 = InData_Switch[29 : 29];
  assign _zz_addra_30 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_30 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_30 = InData_Switch[30 : 30];
  assign _zz_addra_31 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_31 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_31 = InData_Switch[31 : 31];
  assign _zz_addra_32 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_32 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_32 = InData_Switch[32 : 32];
  assign _zz_addra_33 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_33 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_33 = InData_Switch[33 : 33];
  assign _zz_addra_34 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_34 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_34 = InData_Switch[34 : 34];
  assign _zz_addra_35 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_35 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_35 = InData_Switch[35 : 35];
  assign _zz_addra_36 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_36 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_36 = InData_Switch[36 : 36];
  assign _zz_addra_37 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_37 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_37 = InData_Switch[37 : 37];
  assign _zz_addra_38 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_38 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_38 = InData_Switch[38 : 38];
  assign _zz_addra_39 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_39 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_39 = InData_Switch[39 : 39];
  assign _zz_addra_40 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_40 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_40 = InData_Switch[40 : 40];
  assign _zz_addra_41 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_41 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_41 = InData_Switch[41 : 41];
  assign _zz_addra_42 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_42 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_42 = InData_Switch[42 : 42];
  assign _zz_addra_43 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_43 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_43 = InData_Switch[43 : 43];
  assign _zz_addra_44 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_44 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_44 = InData_Switch[44 : 44];
  assign _zz_addra_45 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_45 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_45 = InData_Switch[45 : 45];
  assign _zz_addra_46 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_46 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_46 = InData_Switch[46 : 46];
  assign _zz_addra_47 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_47 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_47 = InData_Switch[47 : 47];
  assign _zz_addra_48 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_48 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_48 = InData_Switch[48 : 48];
  assign _zz_addra_49 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_49 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_49 = InData_Switch[49 : 49];
  assign _zz_addra_50 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_50 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_50 = InData_Switch[50 : 50];
  assign _zz_addra_51 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_51 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_51 = InData_Switch[51 : 51];
  assign _zz_addra_52 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_52 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_52 = InData_Switch[52 : 52];
  assign _zz_addra_53 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_53 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_53 = InData_Switch[53 : 53];
  assign _zz_addra_54 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_54 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_54 = InData_Switch[54 : 54];
  assign _zz_addra_55 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_55 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_55 = InData_Switch[55 : 55];
  assign _zz_addra_56 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_56 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_56 = InData_Switch[56 : 56];
  assign _zz_addra_57 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_57 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_57 = InData_Switch[57 : 57];
  assign _zz_addra_58 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_58 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_58 = InData_Switch[58 : 58];
  assign _zz_addra_59 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_59 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_59 = InData_Switch[59 : 59];
  assign _zz_addra_60 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_60 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_60 = InData_Switch[60 : 60];
  assign _zz_addra_61 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_61 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_61 = InData_Switch[61 : 61];
  assign _zz_addra_62 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_62 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_62 = InData_Switch[62 : 62];
  assign _zz_addra_63 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_63 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_63 = InData_Switch[63 : 63];
  Weight_Bram xil_SimpleDualBram (
    .clka  (clk                           ), //i
    .addra (xil_SimpleDualBram_addra[10:0]), //i
    .dina  (sData_payload[63:0]           ), //i
    .ena   (xil_SimpleDualBram_ena        ), //i
    .wea   (1'b1                          ), //i
    .addrb (xil_SimpleDualBram_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_doutb[7:0] ), //o
    .clkb  (clk                           )  //i
  );
  Weight_Bram xil_SimpleDualBram_1 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_1_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_1_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_1_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_1_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_2 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_2_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_2_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_2_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_2_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_3 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_3_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_3_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_3_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_3_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_4 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_4_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_4_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_4_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_4_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_5 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_5_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_5_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_5_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_5_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_6 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_6_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_6_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_6_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_6_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_7 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_7_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_7_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_7_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_7_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_8 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_8_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_8_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_8_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_8_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_9 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_9_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_9_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_9_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_9_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_10 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_10_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_10_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_10_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_10_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_11 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_11_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_11_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_11_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_11_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_12 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_12_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_12_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_12_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_12_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_13 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_13_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_13_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_13_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_13_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_14 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_14_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_14_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_14_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_14_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_15 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_15_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_15_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_15_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_15_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_16 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_16_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_16_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_16_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_16_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_17 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_17_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_17_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_17_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_17_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_18 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_18_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_18_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_18_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_18_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_19 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_19_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_19_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_19_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_19_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_20 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_20_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_20_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_20_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_20_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_21 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_21_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_21_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_21_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_21_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_22 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_22_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_22_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_22_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_22_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_23 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_23_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_23_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_23_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_23_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_24 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_24_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_24_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_24_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_24_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_25 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_25_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_25_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_25_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_25_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_26 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_26_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_26_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_26_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_26_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_27 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_27_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_27_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_27_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_27_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_28 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_28_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_28_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_28_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_28_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_29 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_29_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_29_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_29_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_29_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_30 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_30_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_30_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_30_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_30_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_31 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_31_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_31_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_31_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_31_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_32 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_32_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_32_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_32_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_32_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_33 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_33_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_33_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_33_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_33_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_34 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_34_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_34_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_34_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_34_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_35 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_35_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_35_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_35_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_35_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_36 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_36_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_36_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_36_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_36_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_37 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_37_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_37_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_37_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_37_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_38 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_38_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_38_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_38_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_38_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_39 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_39_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_39_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_39_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_39_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_40 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_40_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_40_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_40_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_40_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_41 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_41_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_41_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_41_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_41_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_42 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_42_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_42_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_42_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_42_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_43 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_43_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_43_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_43_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_43_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_44 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_44_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_44_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_44_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_44_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_45 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_45_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_45_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_45_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_45_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_46 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_46_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_46_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_46_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_46_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_47 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_47_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_47_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_47_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_47_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_48 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_48_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_48_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_48_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_48_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_49 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_49_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_49_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_49_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_49_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_50 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_50_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_50_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_50_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_50_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_51 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_51_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_51_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_51_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_51_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_52 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_52_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_52_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_52_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_52_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_53 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_53_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_53_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_53_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_53_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_54 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_54_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_54_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_54_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_54_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_55 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_55_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_55_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_55_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_55_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_56 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_56_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_56_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_56_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_56_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_57 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_57_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_57_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_57_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_57_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_58 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_58_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_58_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_58_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_58_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_59 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_59_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_59_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_59_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_59_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_60 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_60_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_60_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_60_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_60_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_61 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_61_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_61_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_61_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_61_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_62 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_62_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_62_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_62_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_62_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_63 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_63_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_63_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_63_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_63_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      WEIGHT_CACHE_STATUS_IDLE : Fsm_currentState_string = "IDLE        ";
      WEIGHT_CACHE_STATUS_INIT : Fsm_currentState_string = "INIT        ";
      WEIGHT_CACHE_STATUS_CACHE_WEIGHT : Fsm_currentState_string = "CACHE_WEIGHT";
      WEIGHT_CACHE_STATUS_SA_COMPUTE : Fsm_currentState_string = "SA_COMPUTE  ";
      default : Fsm_currentState_string = "????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      WEIGHT_CACHE_STATUS_IDLE : Fsm_nextState_string = "IDLE        ";
      WEIGHT_CACHE_STATUS_INIT : Fsm_nextState_string = "INIT        ";
      WEIGHT_CACHE_STATUS_CACHE_WEIGHT : Fsm_nextState_string = "CACHE_WEIGHT";
      WEIGHT_CACHE_STATUS_SA_COMPUTE : Fsm_nextState_string = "SA_COMPUTE  ";
      default : Fsm_nextState_string = "????????????";
    endcase
  end
  `endif

  assign when_SA3D_WeightCache_l33 = (start && (! start_regNext));
  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & WEIGHT_CACHE_STATUS_IDLE) == WEIGHT_CACHE_STATUS_IDLE) : begin
        if(when_SA3D_WeightCache_l33) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_INIT;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_IDLE;
        end
      end
      (((Fsm_currentState) & WEIGHT_CACHE_STATUS_INIT) == WEIGHT_CACHE_STATUS_INIT) : begin
        if(Fsm_Init_End) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_CACHE_WEIGHT;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_INIT;
        end
      end
      (((Fsm_currentState) & WEIGHT_CACHE_STATUS_CACHE_WEIGHT) == WEIGHT_CACHE_STATUS_CACHE_WEIGHT) : begin
        if(Fsm_Weight_All_Cached) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_SA_COMPUTE;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_CACHE_WEIGHT;
        end
      end
      default : begin
        if(Fsm_SA_Computed) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_IDLE;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_SA_COMPUTE;
        end
      end
    endcase
  end

  assign when_WaCounter_l19 = ((Fsm_currentState & WEIGHT_CACHE_STATUS_INIT) != 4'b0000);
  assign when_WaCounter_l14 = (Init_Count_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l14) begin
      Init_Count_valid = 1'b1;
    end else begin
      Init_Count_valid = 1'b0;
    end
  end

  assign Fsm_Init_End = Init_Count_valid;
  assign Matrix_In_MaxCnt = (Matrix_Row >>> 3);
  assign sData_fire = (sData_valid && sData_ready);
  assign In_Row_Cnt_valid = ((In_Row_Cnt_count == _zz_In_Row_Cnt_valid) && sData_fire);
  assign In_Col_Cnt_valid = ((In_Col_Cnt_count == _zz_In_Col_Cnt_valid) && In_Row_Cnt_valid);
  assign when_WaCounter_l40 = (Raddr_Valid && ((Fsm_currentState & WEIGHT_CACHE_STATUS_SA_COMPUTE) != 4'b0000));
  assign OutRow_Cnt_valid = ((OutRow_Cnt_count == _zz_OutRow_Cnt_valid) && when_WaCounter_l40);
  assign _zz_OutCol_Cnt_count = 4'b1000;
  always @(*) begin
    OutCol_Cnt_valid = ((OutCol_Cnt_count <= _zz_OutCol_Cnt_valid) && OutRow_Cnt_valid);
    if(start) begin
      OutCol_Cnt_valid = 1'b0;
    end
  end

  always @(*) begin
    Col_In_8_Cnt_valid = ((Col_In_8_Cnt_count == 6'h3f) && In_Row_Cnt_valid);
    if(OutCol_Cnt_valid) begin
      Col_In_8_Cnt_valid = 1'b0;
    end
  end

  assign when_SA3D_WeightCache_l129 = ((Fsm_currentState & WEIGHT_CACHE_STATUS_INIT) != 4'b0000);
  assign when_SA3D_WeightCache_l134 = ((Fsm_currentState & WEIGHT_CACHE_STATUS_INIT) != 4'b0000);
  assign Fsm_Weight_All_Cached = In_Col_Cnt_valid;
  assign Weight_Cached = In_Col_Cnt_valid;
  assign xil_SimpleDualBram_addra = _zz_addra[10:0];
  assign xil_SimpleDualBram_addrb = _zz_addrb[13:0];
  assign sData_fire_1 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_ena = (_zz_ena[0] && sData_fire_1);
  assign mData_0 = xil_SimpleDualBram_doutb;
  assign xil_SimpleDualBram_1_addra = _zz_addra_1[10:0];
  assign xil_SimpleDualBram_1_addrb = _zz_addrb_1[13:0];
  assign sData_fire_2 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_1_ena = (_zz_ena_1[0] && sData_fire_2);
  assign mData_1 = xil_SimpleDualBram_1_doutb;
  assign xil_SimpleDualBram_2_addra = _zz_addra_2[10:0];
  assign xil_SimpleDualBram_2_addrb = _zz_addrb_2[13:0];
  assign sData_fire_3 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_2_ena = (_zz_ena_2[0] && sData_fire_3);
  assign mData_2 = xil_SimpleDualBram_2_doutb;
  assign xil_SimpleDualBram_3_addra = _zz_addra_3[10:0];
  assign xil_SimpleDualBram_3_addrb = _zz_addrb_3[13:0];
  assign sData_fire_4 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_3_ena = (_zz_ena_3[0] && sData_fire_4);
  assign mData_3 = xil_SimpleDualBram_3_doutb;
  assign xil_SimpleDualBram_4_addra = _zz_addra_4[10:0];
  assign xil_SimpleDualBram_4_addrb = _zz_addrb_4[13:0];
  assign sData_fire_5 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_4_ena = (_zz_ena_4[0] && sData_fire_5);
  assign mData_4 = xil_SimpleDualBram_4_doutb;
  assign xil_SimpleDualBram_5_addra = _zz_addra_5[10:0];
  assign xil_SimpleDualBram_5_addrb = _zz_addrb_5[13:0];
  assign sData_fire_6 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_5_ena = (_zz_ena_5[0] && sData_fire_6);
  assign mData_5 = xil_SimpleDualBram_5_doutb;
  assign xil_SimpleDualBram_6_addra = _zz_addra_6[10:0];
  assign xil_SimpleDualBram_6_addrb = _zz_addrb_6[13:0];
  assign sData_fire_7 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_6_ena = (_zz_ena_6[0] && sData_fire_7);
  assign mData_6 = xil_SimpleDualBram_6_doutb;
  assign xil_SimpleDualBram_7_addra = _zz_addra_7[10:0];
  assign xil_SimpleDualBram_7_addrb = _zz_addrb_7[13:0];
  assign sData_fire_8 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_7_ena = (_zz_ena_7[0] && sData_fire_8);
  assign mData_7 = xil_SimpleDualBram_7_doutb;
  assign xil_SimpleDualBram_8_addra = _zz_addra_8[10:0];
  assign xil_SimpleDualBram_8_addrb = _zz_addrb_8[13:0];
  assign sData_fire_9 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_8_ena = (_zz_ena_8[0] && sData_fire_9);
  assign mData_8 = xil_SimpleDualBram_8_doutb;
  assign xil_SimpleDualBram_9_addra = _zz_addra_9[10:0];
  assign xil_SimpleDualBram_9_addrb = _zz_addrb_9[13:0];
  assign sData_fire_10 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_9_ena = (_zz_ena_9[0] && sData_fire_10);
  assign mData_9 = xil_SimpleDualBram_9_doutb;
  assign xil_SimpleDualBram_10_addra = _zz_addra_10[10:0];
  assign xil_SimpleDualBram_10_addrb = _zz_addrb_10[13:0];
  assign sData_fire_11 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_10_ena = (_zz_ena_10[0] && sData_fire_11);
  assign mData_10 = xil_SimpleDualBram_10_doutb;
  assign xil_SimpleDualBram_11_addra = _zz_addra_11[10:0];
  assign xil_SimpleDualBram_11_addrb = _zz_addrb_11[13:0];
  assign sData_fire_12 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_11_ena = (_zz_ena_11[0] && sData_fire_12);
  assign mData_11 = xil_SimpleDualBram_11_doutb;
  assign xil_SimpleDualBram_12_addra = _zz_addra_12[10:0];
  assign xil_SimpleDualBram_12_addrb = _zz_addrb_12[13:0];
  assign sData_fire_13 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_12_ena = (_zz_ena_12[0] && sData_fire_13);
  assign mData_12 = xil_SimpleDualBram_12_doutb;
  assign xil_SimpleDualBram_13_addra = _zz_addra_13[10:0];
  assign xil_SimpleDualBram_13_addrb = _zz_addrb_13[13:0];
  assign sData_fire_14 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_13_ena = (_zz_ena_13[0] && sData_fire_14);
  assign mData_13 = xil_SimpleDualBram_13_doutb;
  assign xil_SimpleDualBram_14_addra = _zz_addra_14[10:0];
  assign xil_SimpleDualBram_14_addrb = _zz_addrb_14[13:0];
  assign sData_fire_15 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_14_ena = (_zz_ena_14[0] && sData_fire_15);
  assign mData_14 = xil_SimpleDualBram_14_doutb;
  assign xil_SimpleDualBram_15_addra = _zz_addra_15[10:0];
  assign xil_SimpleDualBram_15_addrb = _zz_addrb_15[13:0];
  assign sData_fire_16 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_15_ena = (_zz_ena_15[0] && sData_fire_16);
  assign mData_15 = xil_SimpleDualBram_15_doutb;
  assign xil_SimpleDualBram_16_addra = _zz_addra_16[10:0];
  assign xil_SimpleDualBram_16_addrb = _zz_addrb_16[13:0];
  assign sData_fire_17 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_16_ena = (_zz_ena_16[0] && sData_fire_17);
  assign mData_16 = xil_SimpleDualBram_16_doutb;
  assign xil_SimpleDualBram_17_addra = _zz_addra_17[10:0];
  assign xil_SimpleDualBram_17_addrb = _zz_addrb_17[13:0];
  assign sData_fire_18 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_17_ena = (_zz_ena_17[0] && sData_fire_18);
  assign mData_17 = xil_SimpleDualBram_17_doutb;
  assign xil_SimpleDualBram_18_addra = _zz_addra_18[10:0];
  assign xil_SimpleDualBram_18_addrb = _zz_addrb_18[13:0];
  assign sData_fire_19 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_18_ena = (_zz_ena_18[0] && sData_fire_19);
  assign mData_18 = xil_SimpleDualBram_18_doutb;
  assign xil_SimpleDualBram_19_addra = _zz_addra_19[10:0];
  assign xil_SimpleDualBram_19_addrb = _zz_addrb_19[13:0];
  assign sData_fire_20 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_19_ena = (_zz_ena_19[0] && sData_fire_20);
  assign mData_19 = xil_SimpleDualBram_19_doutb;
  assign xil_SimpleDualBram_20_addra = _zz_addra_20[10:0];
  assign xil_SimpleDualBram_20_addrb = _zz_addrb_20[13:0];
  assign sData_fire_21 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_20_ena = (_zz_ena_20[0] && sData_fire_21);
  assign mData_20 = xil_SimpleDualBram_20_doutb;
  assign xil_SimpleDualBram_21_addra = _zz_addra_21[10:0];
  assign xil_SimpleDualBram_21_addrb = _zz_addrb_21[13:0];
  assign sData_fire_22 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_21_ena = (_zz_ena_21[0] && sData_fire_22);
  assign mData_21 = xil_SimpleDualBram_21_doutb;
  assign xil_SimpleDualBram_22_addra = _zz_addra_22[10:0];
  assign xil_SimpleDualBram_22_addrb = _zz_addrb_22[13:0];
  assign sData_fire_23 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_22_ena = (_zz_ena_22[0] && sData_fire_23);
  assign mData_22 = xil_SimpleDualBram_22_doutb;
  assign xil_SimpleDualBram_23_addra = _zz_addra_23[10:0];
  assign xil_SimpleDualBram_23_addrb = _zz_addrb_23[13:0];
  assign sData_fire_24 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_23_ena = (_zz_ena_23[0] && sData_fire_24);
  assign mData_23 = xil_SimpleDualBram_23_doutb;
  assign xil_SimpleDualBram_24_addra = _zz_addra_24[10:0];
  assign xil_SimpleDualBram_24_addrb = _zz_addrb_24[13:0];
  assign sData_fire_25 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_24_ena = (_zz_ena_24[0] && sData_fire_25);
  assign mData_24 = xil_SimpleDualBram_24_doutb;
  assign xil_SimpleDualBram_25_addra = _zz_addra_25[10:0];
  assign xil_SimpleDualBram_25_addrb = _zz_addrb_25[13:0];
  assign sData_fire_26 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_25_ena = (_zz_ena_25[0] && sData_fire_26);
  assign mData_25 = xil_SimpleDualBram_25_doutb;
  assign xil_SimpleDualBram_26_addra = _zz_addra_26[10:0];
  assign xil_SimpleDualBram_26_addrb = _zz_addrb_26[13:0];
  assign sData_fire_27 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_26_ena = (_zz_ena_26[0] && sData_fire_27);
  assign mData_26 = xil_SimpleDualBram_26_doutb;
  assign xil_SimpleDualBram_27_addra = _zz_addra_27[10:0];
  assign xil_SimpleDualBram_27_addrb = _zz_addrb_27[13:0];
  assign sData_fire_28 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_27_ena = (_zz_ena_27[0] && sData_fire_28);
  assign mData_27 = xil_SimpleDualBram_27_doutb;
  assign xil_SimpleDualBram_28_addra = _zz_addra_28[10:0];
  assign xil_SimpleDualBram_28_addrb = _zz_addrb_28[13:0];
  assign sData_fire_29 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_28_ena = (_zz_ena_28[0] && sData_fire_29);
  assign mData_28 = xil_SimpleDualBram_28_doutb;
  assign xil_SimpleDualBram_29_addra = _zz_addra_29[10:0];
  assign xil_SimpleDualBram_29_addrb = _zz_addrb_29[13:0];
  assign sData_fire_30 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_29_ena = (_zz_ena_29[0] && sData_fire_30);
  assign mData_29 = xil_SimpleDualBram_29_doutb;
  assign xil_SimpleDualBram_30_addra = _zz_addra_30[10:0];
  assign xil_SimpleDualBram_30_addrb = _zz_addrb_30[13:0];
  assign sData_fire_31 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_30_ena = (_zz_ena_30[0] && sData_fire_31);
  assign mData_30 = xil_SimpleDualBram_30_doutb;
  assign xil_SimpleDualBram_31_addra = _zz_addra_31[10:0];
  assign xil_SimpleDualBram_31_addrb = _zz_addrb_31[13:0];
  assign sData_fire_32 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_31_ena = (_zz_ena_31[0] && sData_fire_32);
  assign mData_31 = xil_SimpleDualBram_31_doutb;
  assign xil_SimpleDualBram_32_addra = _zz_addra_32[10:0];
  assign xil_SimpleDualBram_32_addrb = _zz_addrb_32[13:0];
  assign sData_fire_33 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_32_ena = (_zz_ena_32[0] && sData_fire_33);
  assign mData_32 = xil_SimpleDualBram_32_doutb;
  assign xil_SimpleDualBram_33_addra = _zz_addra_33[10:0];
  assign xil_SimpleDualBram_33_addrb = _zz_addrb_33[13:0];
  assign sData_fire_34 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_33_ena = (_zz_ena_33[0] && sData_fire_34);
  assign mData_33 = xil_SimpleDualBram_33_doutb;
  assign xil_SimpleDualBram_34_addra = _zz_addra_34[10:0];
  assign xil_SimpleDualBram_34_addrb = _zz_addrb_34[13:0];
  assign sData_fire_35 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_34_ena = (_zz_ena_34[0] && sData_fire_35);
  assign mData_34 = xil_SimpleDualBram_34_doutb;
  assign xil_SimpleDualBram_35_addra = _zz_addra_35[10:0];
  assign xil_SimpleDualBram_35_addrb = _zz_addrb_35[13:0];
  assign sData_fire_36 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_35_ena = (_zz_ena_35[0] && sData_fire_36);
  assign mData_35 = xil_SimpleDualBram_35_doutb;
  assign xil_SimpleDualBram_36_addra = _zz_addra_36[10:0];
  assign xil_SimpleDualBram_36_addrb = _zz_addrb_36[13:0];
  assign sData_fire_37 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_36_ena = (_zz_ena_36[0] && sData_fire_37);
  assign mData_36 = xil_SimpleDualBram_36_doutb;
  assign xil_SimpleDualBram_37_addra = _zz_addra_37[10:0];
  assign xil_SimpleDualBram_37_addrb = _zz_addrb_37[13:0];
  assign sData_fire_38 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_37_ena = (_zz_ena_37[0] && sData_fire_38);
  assign mData_37 = xil_SimpleDualBram_37_doutb;
  assign xil_SimpleDualBram_38_addra = _zz_addra_38[10:0];
  assign xil_SimpleDualBram_38_addrb = _zz_addrb_38[13:0];
  assign sData_fire_39 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_38_ena = (_zz_ena_38[0] && sData_fire_39);
  assign mData_38 = xil_SimpleDualBram_38_doutb;
  assign xil_SimpleDualBram_39_addra = _zz_addra_39[10:0];
  assign xil_SimpleDualBram_39_addrb = _zz_addrb_39[13:0];
  assign sData_fire_40 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_39_ena = (_zz_ena_39[0] && sData_fire_40);
  assign mData_39 = xil_SimpleDualBram_39_doutb;
  assign xil_SimpleDualBram_40_addra = _zz_addra_40[10:0];
  assign xil_SimpleDualBram_40_addrb = _zz_addrb_40[13:0];
  assign sData_fire_41 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_40_ena = (_zz_ena_40[0] && sData_fire_41);
  assign mData_40 = xil_SimpleDualBram_40_doutb;
  assign xil_SimpleDualBram_41_addra = _zz_addra_41[10:0];
  assign xil_SimpleDualBram_41_addrb = _zz_addrb_41[13:0];
  assign sData_fire_42 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_41_ena = (_zz_ena_41[0] && sData_fire_42);
  assign mData_41 = xil_SimpleDualBram_41_doutb;
  assign xil_SimpleDualBram_42_addra = _zz_addra_42[10:0];
  assign xil_SimpleDualBram_42_addrb = _zz_addrb_42[13:0];
  assign sData_fire_43 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_42_ena = (_zz_ena_42[0] && sData_fire_43);
  assign mData_42 = xil_SimpleDualBram_42_doutb;
  assign xil_SimpleDualBram_43_addra = _zz_addra_43[10:0];
  assign xil_SimpleDualBram_43_addrb = _zz_addrb_43[13:0];
  assign sData_fire_44 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_43_ena = (_zz_ena_43[0] && sData_fire_44);
  assign mData_43 = xil_SimpleDualBram_43_doutb;
  assign xil_SimpleDualBram_44_addra = _zz_addra_44[10:0];
  assign xil_SimpleDualBram_44_addrb = _zz_addrb_44[13:0];
  assign sData_fire_45 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_44_ena = (_zz_ena_44[0] && sData_fire_45);
  assign mData_44 = xil_SimpleDualBram_44_doutb;
  assign xil_SimpleDualBram_45_addra = _zz_addra_45[10:0];
  assign xil_SimpleDualBram_45_addrb = _zz_addrb_45[13:0];
  assign sData_fire_46 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_45_ena = (_zz_ena_45[0] && sData_fire_46);
  assign mData_45 = xil_SimpleDualBram_45_doutb;
  assign xil_SimpleDualBram_46_addra = _zz_addra_46[10:0];
  assign xil_SimpleDualBram_46_addrb = _zz_addrb_46[13:0];
  assign sData_fire_47 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_46_ena = (_zz_ena_46[0] && sData_fire_47);
  assign mData_46 = xil_SimpleDualBram_46_doutb;
  assign xil_SimpleDualBram_47_addra = _zz_addra_47[10:0];
  assign xil_SimpleDualBram_47_addrb = _zz_addrb_47[13:0];
  assign sData_fire_48 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_47_ena = (_zz_ena_47[0] && sData_fire_48);
  assign mData_47 = xil_SimpleDualBram_47_doutb;
  assign xil_SimpleDualBram_48_addra = _zz_addra_48[10:0];
  assign xil_SimpleDualBram_48_addrb = _zz_addrb_48[13:0];
  assign sData_fire_49 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_48_ena = (_zz_ena_48[0] && sData_fire_49);
  assign mData_48 = xil_SimpleDualBram_48_doutb;
  assign xil_SimpleDualBram_49_addra = _zz_addra_49[10:0];
  assign xil_SimpleDualBram_49_addrb = _zz_addrb_49[13:0];
  assign sData_fire_50 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_49_ena = (_zz_ena_49[0] && sData_fire_50);
  assign mData_49 = xil_SimpleDualBram_49_doutb;
  assign xil_SimpleDualBram_50_addra = _zz_addra_50[10:0];
  assign xil_SimpleDualBram_50_addrb = _zz_addrb_50[13:0];
  assign sData_fire_51 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_50_ena = (_zz_ena_50[0] && sData_fire_51);
  assign mData_50 = xil_SimpleDualBram_50_doutb;
  assign xil_SimpleDualBram_51_addra = _zz_addra_51[10:0];
  assign xil_SimpleDualBram_51_addrb = _zz_addrb_51[13:0];
  assign sData_fire_52 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_51_ena = (_zz_ena_51[0] && sData_fire_52);
  assign mData_51 = xil_SimpleDualBram_51_doutb;
  assign xil_SimpleDualBram_52_addra = _zz_addra_52[10:0];
  assign xil_SimpleDualBram_52_addrb = _zz_addrb_52[13:0];
  assign sData_fire_53 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_52_ena = (_zz_ena_52[0] && sData_fire_53);
  assign mData_52 = xil_SimpleDualBram_52_doutb;
  assign xil_SimpleDualBram_53_addra = _zz_addra_53[10:0];
  assign xil_SimpleDualBram_53_addrb = _zz_addrb_53[13:0];
  assign sData_fire_54 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_53_ena = (_zz_ena_53[0] && sData_fire_54);
  assign mData_53 = xil_SimpleDualBram_53_doutb;
  assign xil_SimpleDualBram_54_addra = _zz_addra_54[10:0];
  assign xil_SimpleDualBram_54_addrb = _zz_addrb_54[13:0];
  assign sData_fire_55 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_54_ena = (_zz_ena_54[0] && sData_fire_55);
  assign mData_54 = xil_SimpleDualBram_54_doutb;
  assign xil_SimpleDualBram_55_addra = _zz_addra_55[10:0];
  assign xil_SimpleDualBram_55_addrb = _zz_addrb_55[13:0];
  assign sData_fire_56 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_55_ena = (_zz_ena_55[0] && sData_fire_56);
  assign mData_55 = xil_SimpleDualBram_55_doutb;
  assign xil_SimpleDualBram_56_addra = _zz_addra_56[10:0];
  assign xil_SimpleDualBram_56_addrb = _zz_addrb_56[13:0];
  assign sData_fire_57 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_56_ena = (_zz_ena_56[0] && sData_fire_57);
  assign mData_56 = xil_SimpleDualBram_56_doutb;
  assign xil_SimpleDualBram_57_addra = _zz_addra_57[10:0];
  assign xil_SimpleDualBram_57_addrb = _zz_addrb_57[13:0];
  assign sData_fire_58 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_57_ena = (_zz_ena_57[0] && sData_fire_58);
  assign mData_57 = xil_SimpleDualBram_57_doutb;
  assign xil_SimpleDualBram_58_addra = _zz_addra_58[10:0];
  assign xil_SimpleDualBram_58_addrb = _zz_addrb_58[13:0];
  assign sData_fire_59 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_58_ena = (_zz_ena_58[0] && sData_fire_59);
  assign mData_58 = xil_SimpleDualBram_58_doutb;
  assign xil_SimpleDualBram_59_addra = _zz_addra_59[10:0];
  assign xil_SimpleDualBram_59_addrb = _zz_addrb_59[13:0];
  assign sData_fire_60 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_59_ena = (_zz_ena_59[0] && sData_fire_60);
  assign mData_59 = xil_SimpleDualBram_59_doutb;
  assign xil_SimpleDualBram_60_addra = _zz_addra_60[10:0];
  assign xil_SimpleDualBram_60_addrb = _zz_addrb_60[13:0];
  assign sData_fire_61 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_60_ena = (_zz_ena_60[0] && sData_fire_61);
  assign mData_60 = xil_SimpleDualBram_60_doutb;
  assign xil_SimpleDualBram_61_addra = _zz_addra_61[10:0];
  assign xil_SimpleDualBram_61_addrb = _zz_addrb_61[13:0];
  assign sData_fire_62 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_61_ena = (_zz_ena_61[0] && sData_fire_62);
  assign mData_61 = xil_SimpleDualBram_61_doutb;
  assign xil_SimpleDualBram_62_addra = _zz_addra_62[10:0];
  assign xil_SimpleDualBram_62_addrb = _zz_addrb_62[13:0];
  assign sData_fire_63 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_62_ena = (_zz_ena_62[0] && sData_fire_63);
  assign mData_62 = xil_SimpleDualBram_62_doutb;
  assign xil_SimpleDualBram_63_addra = _zz_addra_63[10:0];
  assign xil_SimpleDualBram_63_addrb = _zz_addrb_63[13:0];
  assign sData_fire_64 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_63_ena = (_zz_ena_63[0] && sData_fire_64);
  assign mData_63 = xil_SimpleDualBram_63_doutb;
  assign sData_ready = ((Fsm_currentState & WEIGHT_CACHE_STATUS_CACHE_WEIGHT) != 4'b0000);
  assign Fsm_SA_Computed = LayerEnd;
  always @(*) begin
    case(OutCol_Cnt_count)
      16'h0001 : begin
        MatrixCol_Switch_1[0 : 0] = 1'b1;
        MatrixCol_Switch_1[63 : 1] = 63'h0;
      end
      16'h0002 : begin
        MatrixCol_Switch_1[1 : 0] = 2'b11;
        MatrixCol_Switch_1[63 : 2] = 62'h0;
      end
      16'h0003 : begin
        MatrixCol_Switch_1[2 : 0] = 3'b111;
        MatrixCol_Switch_1[63 : 3] = 61'h0;
      end
      16'h0004 : begin
        MatrixCol_Switch_1[3 : 0] = 4'b1111;
        MatrixCol_Switch_1[63 : 4] = 60'h0;
      end
      16'h0005 : begin
        MatrixCol_Switch_1[4 : 0] = 5'h1f;
        MatrixCol_Switch_1[63 : 5] = 59'h0;
      end
      16'h0006 : begin
        MatrixCol_Switch_1[5 : 0] = 6'h3f;
        MatrixCol_Switch_1[63 : 6] = 58'h0;
      end
      16'h0007 : begin
        MatrixCol_Switch_1[6 : 0] = 7'h7f;
        MatrixCol_Switch_1[63 : 7] = 57'h0;
      end
      16'h0008 : begin
        MatrixCol_Switch_1[7 : 0] = 8'hff;
        MatrixCol_Switch_1[63 : 8] = 56'h0;
      end
      16'h0009 : begin
        MatrixCol_Switch_1[8 : 0] = 9'h1ff;
        MatrixCol_Switch_1[63 : 9] = 55'h0;
      end
      16'h000a : begin
        MatrixCol_Switch_1[9 : 0] = 10'h3ff;
        MatrixCol_Switch_1[63 : 10] = 54'h0;
      end
      16'h000b : begin
        MatrixCol_Switch_1[10 : 0] = 11'h7ff;
        MatrixCol_Switch_1[63 : 11] = 53'h0;
      end
      16'h000c : begin
        MatrixCol_Switch_1[11 : 0] = 12'hfff;
        MatrixCol_Switch_1[63 : 12] = 52'h0;
      end
      16'h000d : begin
        MatrixCol_Switch_1[12 : 0] = 13'h1fff;
        MatrixCol_Switch_1[63 : 13] = 51'h0;
      end
      16'h000e : begin
        MatrixCol_Switch_1[13 : 0] = 14'h3fff;
        MatrixCol_Switch_1[63 : 14] = 50'h0;
      end
      16'h000f : begin
        MatrixCol_Switch_1[14 : 0] = 15'h7fff;
        MatrixCol_Switch_1[63 : 15] = 49'h0;
      end
      16'h0010 : begin
        MatrixCol_Switch_1[15 : 0] = 16'hffff;
        MatrixCol_Switch_1[63 : 16] = 48'h0;
      end
      16'h0011 : begin
        MatrixCol_Switch_1[16 : 0] = 17'h1ffff;
        MatrixCol_Switch_1[63 : 17] = 47'h0;
      end
      16'h0012 : begin
        MatrixCol_Switch_1[17 : 0] = 18'h3ffff;
        MatrixCol_Switch_1[63 : 18] = 46'h0;
      end
      16'h0013 : begin
        MatrixCol_Switch_1[18 : 0] = 19'h7ffff;
        MatrixCol_Switch_1[63 : 19] = 45'h0;
      end
      16'h0014 : begin
        MatrixCol_Switch_1[19 : 0] = 20'hfffff;
        MatrixCol_Switch_1[63 : 20] = 44'h0;
      end
      16'h0015 : begin
        MatrixCol_Switch_1[20 : 0] = 21'h1fffff;
        MatrixCol_Switch_1[63 : 21] = 43'h0;
      end
      16'h0016 : begin
        MatrixCol_Switch_1[21 : 0] = 22'h3fffff;
        MatrixCol_Switch_1[63 : 22] = 42'h0;
      end
      16'h0017 : begin
        MatrixCol_Switch_1[22 : 0] = 23'h7fffff;
        MatrixCol_Switch_1[63 : 23] = 41'h0;
      end
      16'h0018 : begin
        MatrixCol_Switch_1[23 : 0] = 24'hffffff;
        MatrixCol_Switch_1[63 : 24] = 40'h0;
      end
      16'h0019 : begin
        MatrixCol_Switch_1[24 : 0] = 25'h1ffffff;
        MatrixCol_Switch_1[63 : 25] = 39'h0;
      end
      16'h001a : begin
        MatrixCol_Switch_1[25 : 0] = 26'h3ffffff;
        MatrixCol_Switch_1[63 : 26] = 38'h0;
      end
      16'h001b : begin
        MatrixCol_Switch_1[26 : 0] = 27'h7ffffff;
        MatrixCol_Switch_1[63 : 27] = 37'h0;
      end
      16'h001c : begin
        MatrixCol_Switch_1[27 : 0] = 28'hfffffff;
        MatrixCol_Switch_1[63 : 28] = 36'h0;
      end
      16'h001d : begin
        MatrixCol_Switch_1[28 : 0] = 29'h1fffffff;
        MatrixCol_Switch_1[63 : 29] = 35'h0;
      end
      16'h001e : begin
        MatrixCol_Switch_1[29 : 0] = 30'h3fffffff;
        MatrixCol_Switch_1[63 : 30] = 34'h0;
      end
      16'h001f : begin
        MatrixCol_Switch_1[30 : 0] = 31'h7fffffff;
        MatrixCol_Switch_1[63 : 31] = 33'h0;
      end
      16'h0020 : begin
        MatrixCol_Switch_1[31 : 0] = 32'hffffffff;
        MatrixCol_Switch_1[63 : 32] = 32'h0;
      end
      16'h0021 : begin
        MatrixCol_Switch_1[32 : 0] = 33'h1ffffffff;
        MatrixCol_Switch_1[63 : 33] = 31'h0;
      end
      16'h0022 : begin
        MatrixCol_Switch_1[33 : 0] = 34'h3ffffffff;
        MatrixCol_Switch_1[63 : 34] = 30'h0;
      end
      16'h0023 : begin
        MatrixCol_Switch_1[34 : 0] = 35'h7ffffffff;
        MatrixCol_Switch_1[63 : 35] = 29'h0;
      end
      16'h0024 : begin
        MatrixCol_Switch_1[35 : 0] = 36'hfffffffff;
        MatrixCol_Switch_1[63 : 36] = 28'h0;
      end
      16'h0025 : begin
        MatrixCol_Switch_1[36 : 0] = 37'h1fffffffff;
        MatrixCol_Switch_1[63 : 37] = 27'h0;
      end
      16'h0026 : begin
        MatrixCol_Switch_1[37 : 0] = 38'h3fffffffff;
        MatrixCol_Switch_1[63 : 38] = 26'h0;
      end
      16'h0027 : begin
        MatrixCol_Switch_1[38 : 0] = 39'h7fffffffff;
        MatrixCol_Switch_1[63 : 39] = 25'h0;
      end
      16'h0028 : begin
        MatrixCol_Switch_1[39 : 0] = 40'hffffffffff;
        MatrixCol_Switch_1[63 : 40] = 24'h0;
      end
      16'h0029 : begin
        MatrixCol_Switch_1[40 : 0] = 41'h1ffffffffff;
        MatrixCol_Switch_1[63 : 41] = 23'h0;
      end
      16'h002a : begin
        MatrixCol_Switch_1[41 : 0] = 42'h3ffffffffff;
        MatrixCol_Switch_1[63 : 42] = 22'h0;
      end
      16'h002b : begin
        MatrixCol_Switch_1[42 : 0] = 43'h7ffffffffff;
        MatrixCol_Switch_1[63 : 43] = 21'h0;
      end
      16'h002c : begin
        MatrixCol_Switch_1[43 : 0] = 44'hfffffffffff;
        MatrixCol_Switch_1[63 : 44] = 20'h0;
      end
      16'h002d : begin
        MatrixCol_Switch_1[44 : 0] = 45'h1fffffffffff;
        MatrixCol_Switch_1[63 : 45] = 19'h0;
      end
      16'h002e : begin
        MatrixCol_Switch_1[45 : 0] = 46'h3fffffffffff;
        MatrixCol_Switch_1[63 : 46] = 18'h0;
      end
      16'h002f : begin
        MatrixCol_Switch_1[46 : 0] = 47'h7fffffffffff;
        MatrixCol_Switch_1[63 : 47] = 17'h0;
      end
      16'h0030 : begin
        MatrixCol_Switch_1[47 : 0] = 48'hffffffffffff;
        MatrixCol_Switch_1[63 : 48] = 16'h0;
      end
      16'h0031 : begin
        MatrixCol_Switch_1[48 : 0] = 49'h1ffffffffffff;
        MatrixCol_Switch_1[63 : 49] = 15'h0;
      end
      16'h0032 : begin
        MatrixCol_Switch_1[49 : 0] = 50'h3ffffffffffff;
        MatrixCol_Switch_1[63 : 50] = 14'h0;
      end
      16'h0033 : begin
        MatrixCol_Switch_1[50 : 0] = 51'h7ffffffffffff;
        MatrixCol_Switch_1[63 : 51] = 13'h0;
      end
      16'h0034 : begin
        MatrixCol_Switch_1[51 : 0] = 52'hfffffffffffff;
        MatrixCol_Switch_1[63 : 52] = 12'h0;
      end
      16'h0035 : begin
        MatrixCol_Switch_1[52 : 0] = 53'h1fffffffffffff;
        MatrixCol_Switch_1[63 : 53] = 11'h0;
      end
      16'h0036 : begin
        MatrixCol_Switch_1[53 : 0] = 54'h3fffffffffffff;
        MatrixCol_Switch_1[63 : 54] = 10'h0;
      end
      16'h0037 : begin
        MatrixCol_Switch_1[54 : 0] = 55'h7fffffffffffff;
        MatrixCol_Switch_1[63 : 55] = 9'h0;
      end
      16'h0038 : begin
        MatrixCol_Switch_1[55 : 0] = 56'hffffffffffffff;
        MatrixCol_Switch_1[63 : 56] = 8'h0;
      end
      16'h0039 : begin
        MatrixCol_Switch_1[56 : 0] = 57'h1ffffffffffffff;
        MatrixCol_Switch_1[63 : 57] = 7'h0;
      end
      16'h003a : begin
        MatrixCol_Switch_1[57 : 0] = 58'h3ffffffffffffff;
        MatrixCol_Switch_1[63 : 58] = 6'h0;
      end
      16'h003b : begin
        MatrixCol_Switch_1[58 : 0] = 59'h7ffffffffffffff;
        MatrixCol_Switch_1[63 : 59] = 5'h0;
      end
      16'h003c : begin
        MatrixCol_Switch_1[59 : 0] = 60'hfffffffffffffff;
        MatrixCol_Switch_1[63 : 60] = 4'b0000;
      end
      16'h003d : begin
        MatrixCol_Switch_1[60 : 0] = 61'h1fffffffffffffff;
        MatrixCol_Switch_1[63 : 61] = 3'b000;
      end
      16'h003e : begin
        MatrixCol_Switch_1[61 : 0] = 62'h3fffffffffffffff;
        MatrixCol_Switch_1[63 : 62] = 2'b00;
      end
      16'h003f : begin
        MatrixCol_Switch_1[62 : 0] = 63'h7fffffffffffffff;
        MatrixCol_Switch_1[63 : 63] = 1'b0;
      end
      default : begin
        MatrixCol_Switch_1 = 64'hffffffffffffffff;
      end
    endcase
  end

  assign MatrixCol_Switch = MatrixCol_Switch_1_regNext;
  always @(posedge clk) begin
    start_regNext <= start;
    MatrixCol_Switch_1_regNext <= MatrixCol_Switch_1;
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= WEIGHT_CACHE_STATUS_IDLE;
      Init_Count_count <= 3'b000;
      InData_Switch <= 64'h0000000000000001;
      In_Row_Cnt_count <= 16'h0;
      In_Col_Cnt_count <= 16'h0;
      Read_Row_Base_Addr <= 16'h0;
      Write_Row_Base_Addr <= 16'h0;
      OutRow_Cnt_count <= 16'h0;
      OutCol_Cnt_count <= Matrix_Col;
      Col_In_8_Cnt_count <= 6'h0;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l19) begin
        Init_Count_count <= (Init_Count_count + 3'b001);
        if(Init_Count_valid) begin
          Init_Count_count <= 3'b000;
        end
      end
      if(sData_fire) begin
        if(In_Row_Cnt_valid) begin
          In_Row_Cnt_count <= 16'h0;
        end else begin
          In_Row_Cnt_count <= (In_Row_Cnt_count + 16'h0001);
        end
      end
      if(In_Row_Cnt_valid) begin
        if(In_Col_Cnt_valid) begin
          In_Col_Cnt_count <= 16'h0;
        end else begin
          In_Col_Cnt_count <= (In_Col_Cnt_count + 16'h0001);
        end
      end
      if(when_WaCounter_l40) begin
        if(OutRow_Cnt_valid) begin
          OutRow_Cnt_count <= 16'h0;
        end else begin
          OutRow_Cnt_count <= (OutRow_Cnt_count + 16'h0001);
        end
      end
      if(OutRow_Cnt_valid) begin
        if(OutCol_Cnt_valid) begin
          OutCol_Cnt_count <= Matrix_Col;
        end else begin
          OutCol_Cnt_count <= (OutCol_Cnt_count - _zz_OutCol_Cnt_count_1);
        end
      end
      if(start) begin
        OutCol_Cnt_count <= Matrix_Col;
      end
      if(In_Row_Cnt_valid) begin
        if(Col_In_8_Cnt_valid) begin
          Col_In_8_Cnt_count <= 6'h0;
        end else begin
          Col_In_8_Cnt_count <= (Col_In_8_Cnt_count + 6'h01);
        end
      end
      if(OutCol_Cnt_valid) begin
        Col_In_8_Cnt_count <= 6'h0;
        Read_Row_Base_Addr <= 16'h0;
      end else begin
        if(OutRow_Cnt_valid) begin
          Read_Row_Base_Addr <= (Read_Row_Base_Addr + Matrix_Row);
        end
      end
      if(when_SA3D_WeightCache_l129) begin
        InData_Switch <= 64'h0000000000000001;
      end else begin
        if(In_Row_Cnt_valid) begin
          InData_Switch <= {InData_Switch[62 : 0],InData_Switch[63 : 63]};
        end
      end
      if(when_SA3D_WeightCache_l134) begin
        Write_Row_Base_Addr <= 16'h0;
      end else begin
        if(Col_In_8_Cnt_valid) begin
          Write_Row_Base_Addr <= (Write_Row_Base_Addr + _zz_Write_Row_Base_Addr);
        end
      end
    end
  end


endmodule

//SA_2D_7 replaced by SA_2D

//SA_2D_6 replaced by SA_2D

//SA_2D_5 replaced by SA_2D

//SA_2D_4 replaced by SA_2D

//SA_2D_3 replaced by SA_2D

//SA_2D_2 replaced by SA_2D

//SA_2D_1 replaced by SA_2D

module SA_2D (
  input      [7:0]    io_MatrixA_0,
  input      [7:0]    io_MatrixA_1,
  input      [7:0]    io_MatrixA_2,
  input      [7:0]    io_MatrixA_3,
  input      [7:0]    io_MatrixA_4,
  input      [7:0]    io_MatrixA_5,
  input      [7:0]    io_MatrixA_6,
  input      [7:0]    io_MatrixA_7,
  input      [7:0]    io_MatrixB_0,
  input      [7:0]    io_MatrixB_1,
  input      [7:0]    io_MatrixB_2,
  input      [7:0]    io_MatrixB_3,
  input      [7:0]    io_MatrixB_4,
  input      [7:0]    io_MatrixB_5,
  input      [7:0]    io_MatrixB_6,
  input      [7:0]    io_MatrixB_7,
  input               io_A_Valid_0,
  input               io_A_Valid_1,
  input               io_A_Valid_2,
  input               io_A_Valid_3,
  input               io_A_Valid_4,
  input               io_A_Valid_5,
  input               io_A_Valid_6,
  input               io_A_Valid_7,
  input               io_B_Valid_0,
  input               io_B_Valid_1,
  input               io_B_Valid_2,
  input               io_B_Valid_3,
  input               io_B_Valid_4,
  input               io_B_Valid_5,
  input               io_B_Valid_6,
  input               io_B_Valid_7,
  input      [15:0]   io_signCount,
  output reg [31:0]   MatrixC_0,
  output reg [31:0]   MatrixC_1,
  output reg [31:0]   MatrixC_2,
  output reg [31:0]   MatrixC_3,
  output reg [31:0]   MatrixC_4,
  output reg [31:0]   MatrixC_5,
  output reg [31:0]   MatrixC_6,
  output reg [31:0]   MatrixC_7,
  output              C_Valid_0,
  output              C_Valid_1,
  output              C_Valid_2,
  output              C_Valid_3,
  output              C_Valid_4,
  output              C_Valid_5,
  output              C_Valid_6,
  output              C_Valid_7,
  input               start,
  input               clk,
  input               reset
);

  wire                pE_512_valid;
  wire                pE_513_valid;
  wire                pE_514_valid;
  wire                pE_515_valid;
  wire                pE_516_valid;
  wire                pE_517_valid;
  wire                pE_518_valid;
  wire                pE_519_valid;
  wire                pE_520_valid;
  wire                pE_521_valid;
  wire                pE_522_valid;
  wire                pE_523_valid;
  wire                pE_524_valid;
  wire                pE_525_valid;
  wire                pE_526_valid;
  wire                pE_527_valid;
  wire                pE_528_valid;
  wire                pE_529_valid;
  wire                pE_530_valid;
  wire                pE_531_valid;
  wire                pE_532_valid;
  wire                pE_533_valid;
  wire                pE_534_valid;
  wire                pE_535_valid;
  wire                pE_536_valid;
  wire                pE_537_valid;
  wire                pE_538_valid;
  wire                pE_539_valid;
  wire                pE_540_valid;
  wire                pE_541_valid;
  wire                pE_542_valid;
  wire                pE_543_valid;
  wire                pE_544_valid;
  wire                pE_545_valid;
  wire                pE_546_valid;
  wire                pE_547_valid;
  wire                pE_548_valid;
  wire                pE_549_valid;
  wire                pE_550_valid;
  wire                pE_551_valid;
  wire                pE_552_valid;
  wire                pE_553_valid;
  wire                pE_554_valid;
  wire                pE_555_valid;
  wire                pE_556_valid;
  wire                pE_557_valid;
  wire                pE_558_valid;
  wire                pE_559_valid;
  wire                pE_560_valid;
  wire                pE_561_valid;
  wire                pE_562_valid;
  wire                pE_563_valid;
  wire                pE_564_valid;
  wire                pE_565_valid;
  wire                pE_566_valid;
  wire                pE_567_valid;
  wire                pE_568_valid;
  wire                pE_569_valid;
  wire                pE_570_valid;
  wire                pE_571_valid;
  wire                pE_572_valid;
  wire                pE_573_valid;
  wire                pE_574_valid;
  wire                pE_575_valid;
  wire       [7:0]    pE_512_acount;
  wire       [7:0]    pE_512_bcount;
  wire       [31:0]   pE_512_PE_OUT;
  wire                pE_512_finish;
  wire       [7:0]    pE_513_acount;
  wire       [7:0]    pE_513_bcount;
  wire       [31:0]   pE_513_PE_OUT;
  wire                pE_513_finish;
  wire       [7:0]    pE_514_acount;
  wire       [7:0]    pE_514_bcount;
  wire       [31:0]   pE_514_PE_OUT;
  wire                pE_514_finish;
  wire       [7:0]    pE_515_acount;
  wire       [7:0]    pE_515_bcount;
  wire       [31:0]   pE_515_PE_OUT;
  wire                pE_515_finish;
  wire       [7:0]    pE_516_acount;
  wire       [7:0]    pE_516_bcount;
  wire       [31:0]   pE_516_PE_OUT;
  wire                pE_516_finish;
  wire       [7:0]    pE_517_acount;
  wire       [7:0]    pE_517_bcount;
  wire       [31:0]   pE_517_PE_OUT;
  wire                pE_517_finish;
  wire       [7:0]    pE_518_acount;
  wire       [7:0]    pE_518_bcount;
  wire       [31:0]   pE_518_PE_OUT;
  wire                pE_518_finish;
  wire       [7:0]    pE_519_acount;
  wire       [7:0]    pE_519_bcount;
  wire       [31:0]   pE_519_PE_OUT;
  wire                pE_519_finish;
  wire       [7:0]    pE_520_acount;
  wire       [7:0]    pE_520_bcount;
  wire       [31:0]   pE_520_PE_OUT;
  wire                pE_520_finish;
  wire       [7:0]    pE_521_acount;
  wire       [7:0]    pE_521_bcount;
  wire       [31:0]   pE_521_PE_OUT;
  wire                pE_521_finish;
  wire       [7:0]    pE_522_acount;
  wire       [7:0]    pE_522_bcount;
  wire       [31:0]   pE_522_PE_OUT;
  wire                pE_522_finish;
  wire       [7:0]    pE_523_acount;
  wire       [7:0]    pE_523_bcount;
  wire       [31:0]   pE_523_PE_OUT;
  wire                pE_523_finish;
  wire       [7:0]    pE_524_acount;
  wire       [7:0]    pE_524_bcount;
  wire       [31:0]   pE_524_PE_OUT;
  wire                pE_524_finish;
  wire       [7:0]    pE_525_acount;
  wire       [7:0]    pE_525_bcount;
  wire       [31:0]   pE_525_PE_OUT;
  wire                pE_525_finish;
  wire       [7:0]    pE_526_acount;
  wire       [7:0]    pE_526_bcount;
  wire       [31:0]   pE_526_PE_OUT;
  wire                pE_526_finish;
  wire       [7:0]    pE_527_acount;
  wire       [7:0]    pE_527_bcount;
  wire       [31:0]   pE_527_PE_OUT;
  wire                pE_527_finish;
  wire       [7:0]    pE_528_acount;
  wire       [7:0]    pE_528_bcount;
  wire       [31:0]   pE_528_PE_OUT;
  wire                pE_528_finish;
  wire       [7:0]    pE_529_acount;
  wire       [7:0]    pE_529_bcount;
  wire       [31:0]   pE_529_PE_OUT;
  wire                pE_529_finish;
  wire       [7:0]    pE_530_acount;
  wire       [7:0]    pE_530_bcount;
  wire       [31:0]   pE_530_PE_OUT;
  wire                pE_530_finish;
  wire       [7:0]    pE_531_acount;
  wire       [7:0]    pE_531_bcount;
  wire       [31:0]   pE_531_PE_OUT;
  wire                pE_531_finish;
  wire       [7:0]    pE_532_acount;
  wire       [7:0]    pE_532_bcount;
  wire       [31:0]   pE_532_PE_OUT;
  wire                pE_532_finish;
  wire       [7:0]    pE_533_acount;
  wire       [7:0]    pE_533_bcount;
  wire       [31:0]   pE_533_PE_OUT;
  wire                pE_533_finish;
  wire       [7:0]    pE_534_acount;
  wire       [7:0]    pE_534_bcount;
  wire       [31:0]   pE_534_PE_OUT;
  wire                pE_534_finish;
  wire       [7:0]    pE_535_acount;
  wire       [7:0]    pE_535_bcount;
  wire       [31:0]   pE_535_PE_OUT;
  wire                pE_535_finish;
  wire       [7:0]    pE_536_acount;
  wire       [7:0]    pE_536_bcount;
  wire       [31:0]   pE_536_PE_OUT;
  wire                pE_536_finish;
  wire       [7:0]    pE_537_acount;
  wire       [7:0]    pE_537_bcount;
  wire       [31:0]   pE_537_PE_OUT;
  wire                pE_537_finish;
  wire       [7:0]    pE_538_acount;
  wire       [7:0]    pE_538_bcount;
  wire       [31:0]   pE_538_PE_OUT;
  wire                pE_538_finish;
  wire       [7:0]    pE_539_acount;
  wire       [7:0]    pE_539_bcount;
  wire       [31:0]   pE_539_PE_OUT;
  wire                pE_539_finish;
  wire       [7:0]    pE_540_acount;
  wire       [7:0]    pE_540_bcount;
  wire       [31:0]   pE_540_PE_OUT;
  wire                pE_540_finish;
  wire       [7:0]    pE_541_acount;
  wire       [7:0]    pE_541_bcount;
  wire       [31:0]   pE_541_PE_OUT;
  wire                pE_541_finish;
  wire       [7:0]    pE_542_acount;
  wire       [7:0]    pE_542_bcount;
  wire       [31:0]   pE_542_PE_OUT;
  wire                pE_542_finish;
  wire       [7:0]    pE_543_acount;
  wire       [7:0]    pE_543_bcount;
  wire       [31:0]   pE_543_PE_OUT;
  wire                pE_543_finish;
  wire       [7:0]    pE_544_acount;
  wire       [7:0]    pE_544_bcount;
  wire       [31:0]   pE_544_PE_OUT;
  wire                pE_544_finish;
  wire       [7:0]    pE_545_acount;
  wire       [7:0]    pE_545_bcount;
  wire       [31:0]   pE_545_PE_OUT;
  wire                pE_545_finish;
  wire       [7:0]    pE_546_acount;
  wire       [7:0]    pE_546_bcount;
  wire       [31:0]   pE_546_PE_OUT;
  wire                pE_546_finish;
  wire       [7:0]    pE_547_acount;
  wire       [7:0]    pE_547_bcount;
  wire       [31:0]   pE_547_PE_OUT;
  wire                pE_547_finish;
  wire       [7:0]    pE_548_acount;
  wire       [7:0]    pE_548_bcount;
  wire       [31:0]   pE_548_PE_OUT;
  wire                pE_548_finish;
  wire       [7:0]    pE_549_acount;
  wire       [7:0]    pE_549_bcount;
  wire       [31:0]   pE_549_PE_OUT;
  wire                pE_549_finish;
  wire       [7:0]    pE_550_acount;
  wire       [7:0]    pE_550_bcount;
  wire       [31:0]   pE_550_PE_OUT;
  wire                pE_550_finish;
  wire       [7:0]    pE_551_acount;
  wire       [7:0]    pE_551_bcount;
  wire       [31:0]   pE_551_PE_OUT;
  wire                pE_551_finish;
  wire       [7:0]    pE_552_acount;
  wire       [7:0]    pE_552_bcount;
  wire       [31:0]   pE_552_PE_OUT;
  wire                pE_552_finish;
  wire       [7:0]    pE_553_acount;
  wire       [7:0]    pE_553_bcount;
  wire       [31:0]   pE_553_PE_OUT;
  wire                pE_553_finish;
  wire       [7:0]    pE_554_acount;
  wire       [7:0]    pE_554_bcount;
  wire       [31:0]   pE_554_PE_OUT;
  wire                pE_554_finish;
  wire       [7:0]    pE_555_acount;
  wire       [7:0]    pE_555_bcount;
  wire       [31:0]   pE_555_PE_OUT;
  wire                pE_555_finish;
  wire       [7:0]    pE_556_acount;
  wire       [7:0]    pE_556_bcount;
  wire       [31:0]   pE_556_PE_OUT;
  wire                pE_556_finish;
  wire       [7:0]    pE_557_acount;
  wire       [7:0]    pE_557_bcount;
  wire       [31:0]   pE_557_PE_OUT;
  wire                pE_557_finish;
  wire       [7:0]    pE_558_acount;
  wire       [7:0]    pE_558_bcount;
  wire       [31:0]   pE_558_PE_OUT;
  wire                pE_558_finish;
  wire       [7:0]    pE_559_acount;
  wire       [7:0]    pE_559_bcount;
  wire       [31:0]   pE_559_PE_OUT;
  wire                pE_559_finish;
  wire       [7:0]    pE_560_acount;
  wire       [7:0]    pE_560_bcount;
  wire       [31:0]   pE_560_PE_OUT;
  wire                pE_560_finish;
  wire       [7:0]    pE_561_acount;
  wire       [7:0]    pE_561_bcount;
  wire       [31:0]   pE_561_PE_OUT;
  wire                pE_561_finish;
  wire       [7:0]    pE_562_acount;
  wire       [7:0]    pE_562_bcount;
  wire       [31:0]   pE_562_PE_OUT;
  wire                pE_562_finish;
  wire       [7:0]    pE_563_acount;
  wire       [7:0]    pE_563_bcount;
  wire       [31:0]   pE_563_PE_OUT;
  wire                pE_563_finish;
  wire       [7:0]    pE_564_acount;
  wire       [7:0]    pE_564_bcount;
  wire       [31:0]   pE_564_PE_OUT;
  wire                pE_564_finish;
  wire       [7:0]    pE_565_acount;
  wire       [7:0]    pE_565_bcount;
  wire       [31:0]   pE_565_PE_OUT;
  wire                pE_565_finish;
  wire       [7:0]    pE_566_acount;
  wire       [7:0]    pE_566_bcount;
  wire       [31:0]   pE_566_PE_OUT;
  wire                pE_566_finish;
  wire       [7:0]    pE_567_acount;
  wire       [7:0]    pE_567_bcount;
  wire       [31:0]   pE_567_PE_OUT;
  wire                pE_567_finish;
  wire       [7:0]    pE_568_acount;
  wire       [7:0]    pE_568_bcount;
  wire       [31:0]   pE_568_PE_OUT;
  wire                pE_568_finish;
  wire       [7:0]    pE_569_acount;
  wire       [7:0]    pE_569_bcount;
  wire       [31:0]   pE_569_PE_OUT;
  wire                pE_569_finish;
  wire       [7:0]    pE_570_acount;
  wire       [7:0]    pE_570_bcount;
  wire       [31:0]   pE_570_PE_OUT;
  wire                pE_570_finish;
  wire       [7:0]    pE_571_acount;
  wire       [7:0]    pE_571_bcount;
  wire       [31:0]   pE_571_PE_OUT;
  wire                pE_571_finish;
  wire       [7:0]    pE_572_acount;
  wire       [7:0]    pE_572_bcount;
  wire       [31:0]   pE_572_PE_OUT;
  wire                pE_572_finish;
  wire       [7:0]    pE_573_acount;
  wire       [7:0]    pE_573_bcount;
  wire       [31:0]   pE_573_PE_OUT;
  wire                pE_573_finish;
  wire       [7:0]    pE_574_acount;
  wire       [7:0]    pE_574_bcount;
  wire       [31:0]   pE_574_PE_OUT;
  wire                pE_574_finish;
  wire       [7:0]    pE_575_acount;
  wire       [7:0]    pE_575_bcount;
  wire       [31:0]   pE_575_PE_OUT;
  wire                pE_575_finish;
  reg        [7:0]    tmp;
  wire                when_SA_3D_l80;
  wire                when_SA_3D_l80_1;
  wire                when_SA_3D_l80_2;
  wire                when_SA_3D_l80_3;
  wire                when_SA_3D_l80_4;
  wire                when_SA_3D_l80_5;
  wire                when_SA_3D_l80_6;
  wire                when_SA_3D_l80_7;
  wire                when_SA_3D_l80_8;
  wire                when_SA_3D_l80_9;
  wire                when_SA_3D_l80_10;
  wire                when_SA_3D_l80_11;
  wire                when_SA_3D_l80_12;
  wire                when_SA_3D_l80_13;
  wire                when_SA_3D_l80_14;
  wire                when_SA_3D_l80_15;
  wire                when_SA_3D_l80_16;
  wire                when_SA_3D_l80_17;
  wire                when_SA_3D_l80_18;
  wire                when_SA_3D_l80_19;
  wire                when_SA_3D_l80_20;
  wire                when_SA_3D_l80_21;
  wire                when_SA_3D_l80_22;
  wire                when_SA_3D_l80_23;
  wire                when_SA_3D_l80_24;
  wire                when_SA_3D_l80_25;
  wire                when_SA_3D_l80_26;
  wire                when_SA_3D_l80_27;
  wire                when_SA_3D_l80_28;
  wire                when_SA_3D_l80_29;
  wire                when_SA_3D_l80_30;
  wire                when_SA_3D_l80_31;
  wire                when_SA_3D_l80_32;
  wire                when_SA_3D_l80_33;
  wire                when_SA_3D_l80_34;
  wire                when_SA_3D_l80_35;
  wire                when_SA_3D_l80_36;
  wire                when_SA_3D_l80_37;
  wire                when_SA_3D_l80_38;
  wire                when_SA_3D_l80_39;
  wire                when_SA_3D_l80_40;
  wire                when_SA_3D_l80_41;
  wire                when_SA_3D_l80_42;
  wire                when_SA_3D_l80_43;
  wire                when_SA_3D_l80_44;
  wire                when_SA_3D_l80_45;
  wire                when_SA_3D_l80_46;
  wire                when_SA_3D_l80_47;
  wire                when_SA_3D_l80_48;
  wire                when_SA_3D_l80_49;
  wire                when_SA_3D_l80_50;
  wire                when_SA_3D_l80_51;
  wire                when_SA_3D_l80_52;
  wire                when_SA_3D_l80_53;
  wire                when_SA_3D_l80_54;
  wire                when_SA_3D_l80_55;
  wire                when_SA_3D_l80_56;
  wire                when_SA_3D_l80_57;
  wire                when_SA_3D_l80_58;
  wire                when_SA_3D_l80_59;
  wire                when_SA_3D_l80_60;
  wire                when_SA_3D_l80_61;
  wire                when_SA_3D_l80_62;
  wire                when_SA_3D_l80_63;
  reg        [15:0]   io_signCount_regNextWhen;
  reg                 io_A_Valid_0_delay_1;
  reg                 io_A_Valid_0_delay_1_1;
  reg                 io_A_Valid_0_delay_2;
  reg                 io_A_Valid_0_delay_1_2;
  reg                 io_A_Valid_0_delay_2_1;
  reg                 io_A_Valid_0_delay_3;
  reg                 io_A_Valid_0_delay_1_3;
  reg                 io_A_Valid_0_delay_2_2;
  reg                 io_A_Valid_0_delay_3_1;
  reg                 io_A_Valid_0_delay_4;
  reg                 io_A_Valid_0_delay_1_4;
  reg                 io_A_Valid_0_delay_2_3;
  reg                 io_A_Valid_0_delay_3_2;
  reg                 io_A_Valid_0_delay_4_1;
  reg                 io_A_Valid_0_delay_5;
  reg                 io_A_Valid_0_delay_1_5;
  reg                 io_A_Valid_0_delay_2_4;
  reg                 io_A_Valid_0_delay_3_3;
  reg                 io_A_Valid_0_delay_4_2;
  reg                 io_A_Valid_0_delay_5_1;
  reg                 io_A_Valid_0_delay_6;
  reg                 io_A_Valid_0_delay_1_6;
  reg                 io_A_Valid_0_delay_2_5;
  reg                 io_A_Valid_0_delay_3_4;
  reg                 io_A_Valid_0_delay_4_3;
  reg                 io_A_Valid_0_delay_5_2;
  reg                 io_A_Valid_0_delay_6_1;
  reg                 io_A_Valid_0_delay_7;
  reg        [15:0]   io_signCount_regNextWhen_1;
  reg                 io_B_Valid_0_delay_1;
  reg                 io_A_Valid_1_delay_1;
  reg                 io_B_Valid_1_delay_1;
  reg                 io_A_Valid_1_delay_1_1;
  reg                 io_A_Valid_1_delay_2;
  reg                 io_B_Valid_2_delay_1;
  reg                 io_A_Valid_1_delay_1_2;
  reg                 io_A_Valid_1_delay_2_1;
  reg                 io_A_Valid_1_delay_3;
  reg                 io_B_Valid_3_delay_1;
  reg                 io_A_Valid_1_delay_1_3;
  reg                 io_A_Valid_1_delay_2_2;
  reg                 io_A_Valid_1_delay_3_1;
  reg                 io_A_Valid_1_delay_4;
  reg                 io_B_Valid_4_delay_1;
  reg                 io_A_Valid_1_delay_1_4;
  reg                 io_A_Valid_1_delay_2_3;
  reg                 io_A_Valid_1_delay_3_2;
  reg                 io_A_Valid_1_delay_4_1;
  reg                 io_A_Valid_1_delay_5;
  reg                 io_B_Valid_5_delay_1;
  reg                 io_A_Valid_1_delay_1_5;
  reg                 io_A_Valid_1_delay_2_4;
  reg                 io_A_Valid_1_delay_3_3;
  reg                 io_A_Valid_1_delay_4_2;
  reg                 io_A_Valid_1_delay_5_1;
  reg                 io_A_Valid_1_delay_6;
  reg                 io_B_Valid_6_delay_1;
  reg                 io_A_Valid_1_delay_1_6;
  reg                 io_A_Valid_1_delay_2_5;
  reg                 io_A_Valid_1_delay_3_4;
  reg                 io_A_Valid_1_delay_4_3;
  reg                 io_A_Valid_1_delay_5_2;
  reg                 io_A_Valid_1_delay_6_1;
  reg                 io_A_Valid_1_delay_7;
  reg                 io_B_Valid_7_delay_1;
  reg        [15:0]   io_signCount_regNextWhen_2;
  reg                 io_B_Valid_0_delay_1_1;
  reg                 io_B_Valid_0_delay_2;
  reg                 io_A_Valid_2_delay_1;
  reg                 io_B_Valid_1_delay_1_1;
  reg                 io_B_Valid_1_delay_2;
  reg                 io_A_Valid_2_delay_1_1;
  reg                 io_A_Valid_2_delay_2;
  reg                 io_B_Valid_2_delay_1_1;
  reg                 io_B_Valid_2_delay_2;
  reg                 io_A_Valid_2_delay_1_2;
  reg                 io_A_Valid_2_delay_2_1;
  reg                 io_A_Valid_2_delay_3;
  reg                 io_B_Valid_3_delay_1_1;
  reg                 io_B_Valid_3_delay_2;
  reg                 io_A_Valid_2_delay_1_3;
  reg                 io_A_Valid_2_delay_2_2;
  reg                 io_A_Valid_2_delay_3_1;
  reg                 io_A_Valid_2_delay_4;
  reg                 io_B_Valid_4_delay_1_1;
  reg                 io_B_Valid_4_delay_2;
  reg                 io_A_Valid_2_delay_1_4;
  reg                 io_A_Valid_2_delay_2_3;
  reg                 io_A_Valid_2_delay_3_2;
  reg                 io_A_Valid_2_delay_4_1;
  reg                 io_A_Valid_2_delay_5;
  reg                 io_B_Valid_5_delay_1_1;
  reg                 io_B_Valid_5_delay_2;
  reg                 io_A_Valid_2_delay_1_5;
  reg                 io_A_Valid_2_delay_2_4;
  reg                 io_A_Valid_2_delay_3_3;
  reg                 io_A_Valid_2_delay_4_2;
  reg                 io_A_Valid_2_delay_5_1;
  reg                 io_A_Valid_2_delay_6;
  reg                 io_B_Valid_6_delay_1_1;
  reg                 io_B_Valid_6_delay_2;
  reg                 io_A_Valid_2_delay_1_6;
  reg                 io_A_Valid_2_delay_2_5;
  reg                 io_A_Valid_2_delay_3_4;
  reg                 io_A_Valid_2_delay_4_3;
  reg                 io_A_Valid_2_delay_5_2;
  reg                 io_A_Valid_2_delay_6_1;
  reg                 io_A_Valid_2_delay_7;
  reg                 io_B_Valid_7_delay_1_1;
  reg                 io_B_Valid_7_delay_2;
  reg        [15:0]   io_signCount_regNextWhen_3;
  reg                 io_B_Valid_0_delay_1_2;
  reg                 io_B_Valid_0_delay_2_1;
  reg                 io_B_Valid_0_delay_3;
  reg                 io_A_Valid_3_delay_1;
  reg                 io_B_Valid_1_delay_1_2;
  reg                 io_B_Valid_1_delay_2_1;
  reg                 io_B_Valid_1_delay_3;
  reg                 io_A_Valid_3_delay_1_1;
  reg                 io_A_Valid_3_delay_2;
  reg                 io_B_Valid_2_delay_1_2;
  reg                 io_B_Valid_2_delay_2_1;
  reg                 io_B_Valid_2_delay_3;
  reg                 io_A_Valid_3_delay_1_2;
  reg                 io_A_Valid_3_delay_2_1;
  reg                 io_A_Valid_3_delay_3;
  reg                 io_B_Valid_3_delay_1_2;
  reg                 io_B_Valid_3_delay_2_1;
  reg                 io_B_Valid_3_delay_3;
  reg                 io_A_Valid_3_delay_1_3;
  reg                 io_A_Valid_3_delay_2_2;
  reg                 io_A_Valid_3_delay_3_1;
  reg                 io_A_Valid_3_delay_4;
  reg                 io_B_Valid_4_delay_1_2;
  reg                 io_B_Valid_4_delay_2_1;
  reg                 io_B_Valid_4_delay_3;
  reg                 io_A_Valid_3_delay_1_4;
  reg                 io_A_Valid_3_delay_2_3;
  reg                 io_A_Valid_3_delay_3_2;
  reg                 io_A_Valid_3_delay_4_1;
  reg                 io_A_Valid_3_delay_5;
  reg                 io_B_Valid_5_delay_1_2;
  reg                 io_B_Valid_5_delay_2_1;
  reg                 io_B_Valid_5_delay_3;
  reg                 io_A_Valid_3_delay_1_5;
  reg                 io_A_Valid_3_delay_2_4;
  reg                 io_A_Valid_3_delay_3_3;
  reg                 io_A_Valid_3_delay_4_2;
  reg                 io_A_Valid_3_delay_5_1;
  reg                 io_A_Valid_3_delay_6;
  reg                 io_B_Valid_6_delay_1_2;
  reg                 io_B_Valid_6_delay_2_1;
  reg                 io_B_Valid_6_delay_3;
  reg                 io_A_Valid_3_delay_1_6;
  reg                 io_A_Valid_3_delay_2_5;
  reg                 io_A_Valid_3_delay_3_4;
  reg                 io_A_Valid_3_delay_4_3;
  reg                 io_A_Valid_3_delay_5_2;
  reg                 io_A_Valid_3_delay_6_1;
  reg                 io_A_Valid_3_delay_7;
  reg                 io_B_Valid_7_delay_1_2;
  reg                 io_B_Valid_7_delay_2_1;
  reg                 io_B_Valid_7_delay_3;
  reg        [15:0]   io_signCount_regNextWhen_4;
  reg                 io_B_Valid_0_delay_1_3;
  reg                 io_B_Valid_0_delay_2_2;
  reg                 io_B_Valid_0_delay_3_1;
  reg                 io_B_Valid_0_delay_4;
  reg                 io_A_Valid_4_delay_1;
  reg                 io_B_Valid_1_delay_1_3;
  reg                 io_B_Valid_1_delay_2_2;
  reg                 io_B_Valid_1_delay_3_1;
  reg                 io_B_Valid_1_delay_4;
  reg                 io_A_Valid_4_delay_1_1;
  reg                 io_A_Valid_4_delay_2;
  reg                 io_B_Valid_2_delay_1_3;
  reg                 io_B_Valid_2_delay_2_2;
  reg                 io_B_Valid_2_delay_3_1;
  reg                 io_B_Valid_2_delay_4;
  reg                 io_A_Valid_4_delay_1_2;
  reg                 io_A_Valid_4_delay_2_1;
  reg                 io_A_Valid_4_delay_3;
  reg                 io_B_Valid_3_delay_1_3;
  reg                 io_B_Valid_3_delay_2_2;
  reg                 io_B_Valid_3_delay_3_1;
  reg                 io_B_Valid_3_delay_4;
  reg                 io_A_Valid_4_delay_1_3;
  reg                 io_A_Valid_4_delay_2_2;
  reg                 io_A_Valid_4_delay_3_1;
  reg                 io_A_Valid_4_delay_4;
  reg                 io_B_Valid_4_delay_1_3;
  reg                 io_B_Valid_4_delay_2_2;
  reg                 io_B_Valid_4_delay_3_1;
  reg                 io_B_Valid_4_delay_4;
  reg                 io_A_Valid_4_delay_1_4;
  reg                 io_A_Valid_4_delay_2_3;
  reg                 io_A_Valid_4_delay_3_2;
  reg                 io_A_Valid_4_delay_4_1;
  reg                 io_A_Valid_4_delay_5;
  reg                 io_B_Valid_5_delay_1_3;
  reg                 io_B_Valid_5_delay_2_2;
  reg                 io_B_Valid_5_delay_3_1;
  reg                 io_B_Valid_5_delay_4;
  reg                 io_A_Valid_4_delay_1_5;
  reg                 io_A_Valid_4_delay_2_4;
  reg                 io_A_Valid_4_delay_3_3;
  reg                 io_A_Valid_4_delay_4_2;
  reg                 io_A_Valid_4_delay_5_1;
  reg                 io_A_Valid_4_delay_6;
  reg                 io_B_Valid_6_delay_1_3;
  reg                 io_B_Valid_6_delay_2_2;
  reg                 io_B_Valid_6_delay_3_1;
  reg                 io_B_Valid_6_delay_4;
  reg                 io_A_Valid_4_delay_1_6;
  reg                 io_A_Valid_4_delay_2_5;
  reg                 io_A_Valid_4_delay_3_4;
  reg                 io_A_Valid_4_delay_4_3;
  reg                 io_A_Valid_4_delay_5_2;
  reg                 io_A_Valid_4_delay_6_1;
  reg                 io_A_Valid_4_delay_7;
  reg                 io_B_Valid_7_delay_1_3;
  reg                 io_B_Valid_7_delay_2_2;
  reg                 io_B_Valid_7_delay_3_1;
  reg                 io_B_Valid_7_delay_4;
  reg        [15:0]   io_signCount_regNextWhen_5;
  reg                 io_B_Valid_0_delay_1_4;
  reg                 io_B_Valid_0_delay_2_3;
  reg                 io_B_Valid_0_delay_3_2;
  reg                 io_B_Valid_0_delay_4_1;
  reg                 io_B_Valid_0_delay_5;
  reg                 io_A_Valid_5_delay_1;
  reg                 io_B_Valid_1_delay_1_4;
  reg                 io_B_Valid_1_delay_2_3;
  reg                 io_B_Valid_1_delay_3_2;
  reg                 io_B_Valid_1_delay_4_1;
  reg                 io_B_Valid_1_delay_5;
  reg                 io_A_Valid_5_delay_1_1;
  reg                 io_A_Valid_5_delay_2;
  reg                 io_B_Valid_2_delay_1_4;
  reg                 io_B_Valid_2_delay_2_3;
  reg                 io_B_Valid_2_delay_3_2;
  reg                 io_B_Valid_2_delay_4_1;
  reg                 io_B_Valid_2_delay_5;
  reg                 io_A_Valid_5_delay_1_2;
  reg                 io_A_Valid_5_delay_2_1;
  reg                 io_A_Valid_5_delay_3;
  reg                 io_B_Valid_3_delay_1_4;
  reg                 io_B_Valid_3_delay_2_3;
  reg                 io_B_Valid_3_delay_3_2;
  reg                 io_B_Valid_3_delay_4_1;
  reg                 io_B_Valid_3_delay_5;
  reg                 io_A_Valid_5_delay_1_3;
  reg                 io_A_Valid_5_delay_2_2;
  reg                 io_A_Valid_5_delay_3_1;
  reg                 io_A_Valid_5_delay_4;
  reg                 io_B_Valid_4_delay_1_4;
  reg                 io_B_Valid_4_delay_2_3;
  reg                 io_B_Valid_4_delay_3_2;
  reg                 io_B_Valid_4_delay_4_1;
  reg                 io_B_Valid_4_delay_5;
  reg                 io_A_Valid_5_delay_1_4;
  reg                 io_A_Valid_5_delay_2_3;
  reg                 io_A_Valid_5_delay_3_2;
  reg                 io_A_Valid_5_delay_4_1;
  reg                 io_A_Valid_5_delay_5;
  reg                 io_B_Valid_5_delay_1_4;
  reg                 io_B_Valid_5_delay_2_3;
  reg                 io_B_Valid_5_delay_3_2;
  reg                 io_B_Valid_5_delay_4_1;
  reg                 io_B_Valid_5_delay_5;
  reg                 io_A_Valid_5_delay_1_5;
  reg                 io_A_Valid_5_delay_2_4;
  reg                 io_A_Valid_5_delay_3_3;
  reg                 io_A_Valid_5_delay_4_2;
  reg                 io_A_Valid_5_delay_5_1;
  reg                 io_A_Valid_5_delay_6;
  reg                 io_B_Valid_6_delay_1_4;
  reg                 io_B_Valid_6_delay_2_3;
  reg                 io_B_Valid_6_delay_3_2;
  reg                 io_B_Valid_6_delay_4_1;
  reg                 io_B_Valid_6_delay_5;
  reg                 io_A_Valid_5_delay_1_6;
  reg                 io_A_Valid_5_delay_2_5;
  reg                 io_A_Valid_5_delay_3_4;
  reg                 io_A_Valid_5_delay_4_3;
  reg                 io_A_Valid_5_delay_5_2;
  reg                 io_A_Valid_5_delay_6_1;
  reg                 io_A_Valid_5_delay_7;
  reg                 io_B_Valid_7_delay_1_4;
  reg                 io_B_Valid_7_delay_2_3;
  reg                 io_B_Valid_7_delay_3_2;
  reg                 io_B_Valid_7_delay_4_1;
  reg                 io_B_Valid_7_delay_5;
  reg        [15:0]   io_signCount_regNextWhen_6;
  reg                 io_B_Valid_0_delay_1_5;
  reg                 io_B_Valid_0_delay_2_4;
  reg                 io_B_Valid_0_delay_3_3;
  reg                 io_B_Valid_0_delay_4_2;
  reg                 io_B_Valid_0_delay_5_1;
  reg                 io_B_Valid_0_delay_6;
  reg                 io_A_Valid_6_delay_1;
  reg                 io_B_Valid_1_delay_1_5;
  reg                 io_B_Valid_1_delay_2_4;
  reg                 io_B_Valid_1_delay_3_3;
  reg                 io_B_Valid_1_delay_4_2;
  reg                 io_B_Valid_1_delay_5_1;
  reg                 io_B_Valid_1_delay_6;
  reg                 io_A_Valid_6_delay_1_1;
  reg                 io_A_Valid_6_delay_2;
  reg                 io_B_Valid_2_delay_1_5;
  reg                 io_B_Valid_2_delay_2_4;
  reg                 io_B_Valid_2_delay_3_3;
  reg                 io_B_Valid_2_delay_4_2;
  reg                 io_B_Valid_2_delay_5_1;
  reg                 io_B_Valid_2_delay_6;
  reg                 io_A_Valid_6_delay_1_2;
  reg                 io_A_Valid_6_delay_2_1;
  reg                 io_A_Valid_6_delay_3;
  reg                 io_B_Valid_3_delay_1_5;
  reg                 io_B_Valid_3_delay_2_4;
  reg                 io_B_Valid_3_delay_3_3;
  reg                 io_B_Valid_3_delay_4_2;
  reg                 io_B_Valid_3_delay_5_1;
  reg                 io_B_Valid_3_delay_6;
  reg                 io_A_Valid_6_delay_1_3;
  reg                 io_A_Valid_6_delay_2_2;
  reg                 io_A_Valid_6_delay_3_1;
  reg                 io_A_Valid_6_delay_4;
  reg                 io_B_Valid_4_delay_1_5;
  reg                 io_B_Valid_4_delay_2_4;
  reg                 io_B_Valid_4_delay_3_3;
  reg                 io_B_Valid_4_delay_4_2;
  reg                 io_B_Valid_4_delay_5_1;
  reg                 io_B_Valid_4_delay_6;
  reg                 io_A_Valid_6_delay_1_4;
  reg                 io_A_Valid_6_delay_2_3;
  reg                 io_A_Valid_6_delay_3_2;
  reg                 io_A_Valid_6_delay_4_1;
  reg                 io_A_Valid_6_delay_5;
  reg                 io_B_Valid_5_delay_1_5;
  reg                 io_B_Valid_5_delay_2_4;
  reg                 io_B_Valid_5_delay_3_3;
  reg                 io_B_Valid_5_delay_4_2;
  reg                 io_B_Valid_5_delay_5_1;
  reg                 io_B_Valid_5_delay_6;
  reg                 io_A_Valid_6_delay_1_5;
  reg                 io_A_Valid_6_delay_2_4;
  reg                 io_A_Valid_6_delay_3_3;
  reg                 io_A_Valid_6_delay_4_2;
  reg                 io_A_Valid_6_delay_5_1;
  reg                 io_A_Valid_6_delay_6;
  reg                 io_B_Valid_6_delay_1_5;
  reg                 io_B_Valid_6_delay_2_4;
  reg                 io_B_Valid_6_delay_3_3;
  reg                 io_B_Valid_6_delay_4_2;
  reg                 io_B_Valid_6_delay_5_1;
  reg                 io_B_Valid_6_delay_6;
  reg                 io_A_Valid_6_delay_1_6;
  reg                 io_A_Valid_6_delay_2_5;
  reg                 io_A_Valid_6_delay_3_4;
  reg                 io_A_Valid_6_delay_4_3;
  reg                 io_A_Valid_6_delay_5_2;
  reg                 io_A_Valid_6_delay_6_1;
  reg                 io_A_Valid_6_delay_7;
  reg                 io_B_Valid_7_delay_1_5;
  reg                 io_B_Valid_7_delay_2_4;
  reg                 io_B_Valid_7_delay_3_3;
  reg                 io_B_Valid_7_delay_4_2;
  reg                 io_B_Valid_7_delay_5_1;
  reg                 io_B_Valid_7_delay_6;
  reg        [15:0]   io_signCount_regNextWhen_7;
  reg                 io_B_Valid_0_delay_1_6;
  reg                 io_B_Valid_0_delay_2_5;
  reg                 io_B_Valid_0_delay_3_4;
  reg                 io_B_Valid_0_delay_4_3;
  reg                 io_B_Valid_0_delay_5_2;
  reg                 io_B_Valid_0_delay_6_1;
  reg                 io_B_Valid_0_delay_7;
  reg                 io_A_Valid_7_delay_1;
  reg                 io_B_Valid_1_delay_1_6;
  reg                 io_B_Valid_1_delay_2_5;
  reg                 io_B_Valid_1_delay_3_4;
  reg                 io_B_Valid_1_delay_4_3;
  reg                 io_B_Valid_1_delay_5_2;
  reg                 io_B_Valid_1_delay_6_1;
  reg                 io_B_Valid_1_delay_7;
  reg                 io_A_Valid_7_delay_1_1;
  reg                 io_A_Valid_7_delay_2;
  reg                 io_B_Valid_2_delay_1_6;
  reg                 io_B_Valid_2_delay_2_5;
  reg                 io_B_Valid_2_delay_3_4;
  reg                 io_B_Valid_2_delay_4_3;
  reg                 io_B_Valid_2_delay_5_2;
  reg                 io_B_Valid_2_delay_6_1;
  reg                 io_B_Valid_2_delay_7;
  reg                 io_A_Valid_7_delay_1_2;
  reg                 io_A_Valid_7_delay_2_1;
  reg                 io_A_Valid_7_delay_3;
  reg                 io_B_Valid_3_delay_1_6;
  reg                 io_B_Valid_3_delay_2_5;
  reg                 io_B_Valid_3_delay_3_4;
  reg                 io_B_Valid_3_delay_4_3;
  reg                 io_B_Valid_3_delay_5_2;
  reg                 io_B_Valid_3_delay_6_1;
  reg                 io_B_Valid_3_delay_7;
  reg                 io_A_Valid_7_delay_1_3;
  reg                 io_A_Valid_7_delay_2_2;
  reg                 io_A_Valid_7_delay_3_1;
  reg                 io_A_Valid_7_delay_4;
  reg                 io_B_Valid_4_delay_1_6;
  reg                 io_B_Valid_4_delay_2_5;
  reg                 io_B_Valid_4_delay_3_4;
  reg                 io_B_Valid_4_delay_4_3;
  reg                 io_B_Valid_4_delay_5_2;
  reg                 io_B_Valid_4_delay_6_1;
  reg                 io_B_Valid_4_delay_7;
  reg                 io_A_Valid_7_delay_1_4;
  reg                 io_A_Valid_7_delay_2_3;
  reg                 io_A_Valid_7_delay_3_2;
  reg                 io_A_Valid_7_delay_4_1;
  reg                 io_A_Valid_7_delay_5;
  reg                 io_B_Valid_5_delay_1_6;
  reg                 io_B_Valid_5_delay_2_5;
  reg                 io_B_Valid_5_delay_3_4;
  reg                 io_B_Valid_5_delay_4_3;
  reg                 io_B_Valid_5_delay_5_2;
  reg                 io_B_Valid_5_delay_6_1;
  reg                 io_B_Valid_5_delay_7;
  reg                 io_A_Valid_7_delay_1_5;
  reg                 io_A_Valid_7_delay_2_4;
  reg                 io_A_Valid_7_delay_3_3;
  reg                 io_A_Valid_7_delay_4_2;
  reg                 io_A_Valid_7_delay_5_1;
  reg                 io_A_Valid_7_delay_6;
  reg                 io_B_Valid_6_delay_1_6;
  reg                 io_B_Valid_6_delay_2_5;
  reg                 io_B_Valid_6_delay_3_4;
  reg                 io_B_Valid_6_delay_4_3;
  reg                 io_B_Valid_6_delay_5_2;
  reg                 io_B_Valid_6_delay_6_1;
  reg                 io_B_Valid_6_delay_7;
  reg                 io_A_Valid_7_delay_1_6;
  reg                 io_A_Valid_7_delay_2_5;
  reg                 io_A_Valid_7_delay_3_4;
  reg                 io_A_Valid_7_delay_4_3;
  reg                 io_A_Valid_7_delay_5_2;
  reg                 io_A_Valid_7_delay_6_1;
  reg                 io_A_Valid_7_delay_7;
  reg                 io_B_Valid_7_delay_1_6;
  reg                 io_B_Valid_7_delay_2_5;
  reg                 io_B_Valid_7_delay_3_4;
  reg                 io_B_Valid_7_delay_4_3;
  reg                 io_B_Valid_7_delay_5_2;
  reg                 io_B_Valid_7_delay_6_1;
  reg                 io_B_Valid_7_delay_7;

  PE_448 pE_512 (
    .activate  (io_MatrixA_0[7:0]             ), //i
    .weight    (io_MatrixB_0[7:0]             ), //i
    .valid     (pE_512_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_512_acount[7:0]            ), //o
    .bcount    (pE_512_bcount[7:0]            ), //o
    .PE_OUT    (pE_512_PE_OUT[31:0]           ), //o
    .finish    (pE_512_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_513 (
    .activate  (pE_512_acount[7:0]            ), //i
    .weight    (io_MatrixB_1[7:0]             ), //i
    .valid     (pE_513_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_513_acount[7:0]            ), //o
    .bcount    (pE_513_bcount[7:0]            ), //o
    .PE_OUT    (pE_513_PE_OUT[31:0]           ), //o
    .finish    (pE_513_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_514 (
    .activate  (pE_513_acount[7:0]            ), //i
    .weight    (io_MatrixB_2[7:0]             ), //i
    .valid     (pE_514_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_514_acount[7:0]            ), //o
    .bcount    (pE_514_bcount[7:0]            ), //o
    .PE_OUT    (pE_514_PE_OUT[31:0]           ), //o
    .finish    (pE_514_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_515 (
    .activate  (pE_514_acount[7:0]            ), //i
    .weight    (io_MatrixB_3[7:0]             ), //i
    .valid     (pE_515_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_515_acount[7:0]            ), //o
    .bcount    (pE_515_bcount[7:0]            ), //o
    .PE_OUT    (pE_515_PE_OUT[31:0]           ), //o
    .finish    (pE_515_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_516 (
    .activate  (pE_515_acount[7:0]            ), //i
    .weight    (io_MatrixB_4[7:0]             ), //i
    .valid     (pE_516_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_516_acount[7:0]            ), //o
    .bcount    (pE_516_bcount[7:0]            ), //o
    .PE_OUT    (pE_516_PE_OUT[31:0]           ), //o
    .finish    (pE_516_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_517 (
    .activate  (pE_516_acount[7:0]            ), //i
    .weight    (io_MatrixB_5[7:0]             ), //i
    .valid     (pE_517_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_517_acount[7:0]            ), //o
    .bcount    (pE_517_bcount[7:0]            ), //o
    .PE_OUT    (pE_517_PE_OUT[31:0]           ), //o
    .finish    (pE_517_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_518 (
    .activate  (pE_517_acount[7:0]            ), //i
    .weight    (io_MatrixB_6[7:0]             ), //i
    .valid     (pE_518_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_518_acount[7:0]            ), //o
    .bcount    (pE_518_bcount[7:0]            ), //o
    .PE_OUT    (pE_518_PE_OUT[31:0]           ), //o
    .finish    (pE_518_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_519 (
    .activate  (pE_518_acount[7:0]            ), //i
    .weight    (io_MatrixB_7[7:0]             ), //i
    .valid     (pE_519_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_519_acount[7:0]            ), //o
    .bcount    (pE_519_bcount[7:0]            ), //o
    .PE_OUT    (pE_519_PE_OUT[31:0]           ), //o
    .finish    (pE_519_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_520 (
    .activate  (pE_520_acount[7:0]              ), //i
    .weight    (pE_512_bcount[7:0]              ), //i
    .valid     (pE_520_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_520_acount[7:0]              ), //o
    .bcount    (pE_520_bcount[7:0]              ), //o
    .PE_OUT    (pE_520_PE_OUT[31:0]             ), //o
    .finish    (pE_520_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_521 (
    .activate  (pE_512_acount[7:0]              ), //i
    .weight    (pE_512_bcount[7:0]              ), //i
    .valid     (pE_521_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_521_acount[7:0]              ), //o
    .bcount    (pE_521_bcount[7:0]              ), //o
    .PE_OUT    (pE_521_PE_OUT[31:0]             ), //o
    .finish    (pE_521_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_522 (
    .activate  (pE_513_acount[7:0]              ), //i
    .weight    (pE_513_bcount[7:0]              ), //i
    .valid     (pE_522_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_522_acount[7:0]              ), //o
    .bcount    (pE_522_bcount[7:0]              ), //o
    .PE_OUT    (pE_522_PE_OUT[31:0]             ), //o
    .finish    (pE_522_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_523 (
    .activate  (pE_514_acount[7:0]              ), //i
    .weight    (pE_514_bcount[7:0]              ), //i
    .valid     (pE_523_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_523_acount[7:0]              ), //o
    .bcount    (pE_523_bcount[7:0]              ), //o
    .PE_OUT    (pE_523_PE_OUT[31:0]             ), //o
    .finish    (pE_523_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_524 (
    .activate  (pE_515_acount[7:0]              ), //i
    .weight    (pE_515_bcount[7:0]              ), //i
    .valid     (pE_524_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_524_acount[7:0]              ), //o
    .bcount    (pE_524_bcount[7:0]              ), //o
    .PE_OUT    (pE_524_PE_OUT[31:0]             ), //o
    .finish    (pE_524_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_525 (
    .activate  (pE_516_acount[7:0]              ), //i
    .weight    (pE_516_bcount[7:0]              ), //i
    .valid     (pE_525_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_525_acount[7:0]              ), //o
    .bcount    (pE_525_bcount[7:0]              ), //o
    .PE_OUT    (pE_525_PE_OUT[31:0]             ), //o
    .finish    (pE_525_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_526 (
    .activate  (pE_517_acount[7:0]              ), //i
    .weight    (pE_517_bcount[7:0]              ), //i
    .valid     (pE_526_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_526_acount[7:0]              ), //o
    .bcount    (pE_526_bcount[7:0]              ), //o
    .PE_OUT    (pE_526_PE_OUT[31:0]             ), //o
    .finish    (pE_526_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_527 (
    .activate  (pE_518_acount[7:0]              ), //i
    .weight    (pE_518_bcount[7:0]              ), //i
    .valid     (pE_527_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_527_acount[7:0]              ), //o
    .bcount    (pE_527_bcount[7:0]              ), //o
    .PE_OUT    (pE_527_PE_OUT[31:0]             ), //o
    .finish    (pE_527_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_528 (
    .activate  (pE_528_acount[7:0]              ), //i
    .weight    (pE_520_bcount[7:0]              ), //i
    .valid     (pE_528_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_528_acount[7:0]              ), //o
    .bcount    (pE_528_bcount[7:0]              ), //o
    .PE_OUT    (pE_528_PE_OUT[31:0]             ), //o
    .finish    (pE_528_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_529 (
    .activate  (pE_520_acount[7:0]              ), //i
    .weight    (pE_520_bcount[7:0]              ), //i
    .valid     (pE_529_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_529_acount[7:0]              ), //o
    .bcount    (pE_529_bcount[7:0]              ), //o
    .PE_OUT    (pE_529_PE_OUT[31:0]             ), //o
    .finish    (pE_529_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_530 (
    .activate  (pE_521_acount[7:0]              ), //i
    .weight    (pE_521_bcount[7:0]              ), //i
    .valid     (pE_530_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_530_acount[7:0]              ), //o
    .bcount    (pE_530_bcount[7:0]              ), //o
    .PE_OUT    (pE_530_PE_OUT[31:0]             ), //o
    .finish    (pE_530_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_531 (
    .activate  (pE_522_acount[7:0]              ), //i
    .weight    (pE_522_bcount[7:0]              ), //i
    .valid     (pE_531_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_531_acount[7:0]              ), //o
    .bcount    (pE_531_bcount[7:0]              ), //o
    .PE_OUT    (pE_531_PE_OUT[31:0]             ), //o
    .finish    (pE_531_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_532 (
    .activate  (pE_523_acount[7:0]              ), //i
    .weight    (pE_523_bcount[7:0]              ), //i
    .valid     (pE_532_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_532_acount[7:0]              ), //o
    .bcount    (pE_532_bcount[7:0]              ), //o
    .PE_OUT    (pE_532_PE_OUT[31:0]             ), //o
    .finish    (pE_532_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_533 (
    .activate  (pE_524_acount[7:0]              ), //i
    .weight    (pE_524_bcount[7:0]              ), //i
    .valid     (pE_533_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_533_acount[7:0]              ), //o
    .bcount    (pE_533_bcount[7:0]              ), //o
    .PE_OUT    (pE_533_PE_OUT[31:0]             ), //o
    .finish    (pE_533_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_534 (
    .activate  (pE_525_acount[7:0]              ), //i
    .weight    (pE_525_bcount[7:0]              ), //i
    .valid     (pE_534_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_534_acount[7:0]              ), //o
    .bcount    (pE_534_bcount[7:0]              ), //o
    .PE_OUT    (pE_534_PE_OUT[31:0]             ), //o
    .finish    (pE_534_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_535 (
    .activate  (pE_526_acount[7:0]              ), //i
    .weight    (pE_526_bcount[7:0]              ), //i
    .valid     (pE_535_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_535_acount[7:0]              ), //o
    .bcount    (pE_535_bcount[7:0]              ), //o
    .PE_OUT    (pE_535_PE_OUT[31:0]             ), //o
    .finish    (pE_535_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_536 (
    .activate  (pE_536_acount[7:0]              ), //i
    .weight    (pE_528_bcount[7:0]              ), //i
    .valid     (pE_536_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_536_acount[7:0]              ), //o
    .bcount    (pE_536_bcount[7:0]              ), //o
    .PE_OUT    (pE_536_PE_OUT[31:0]             ), //o
    .finish    (pE_536_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_537 (
    .activate  (pE_528_acount[7:0]              ), //i
    .weight    (pE_528_bcount[7:0]              ), //i
    .valid     (pE_537_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_537_acount[7:0]              ), //o
    .bcount    (pE_537_bcount[7:0]              ), //o
    .PE_OUT    (pE_537_PE_OUT[31:0]             ), //o
    .finish    (pE_537_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_538 (
    .activate  (pE_529_acount[7:0]              ), //i
    .weight    (pE_529_bcount[7:0]              ), //i
    .valid     (pE_538_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_538_acount[7:0]              ), //o
    .bcount    (pE_538_bcount[7:0]              ), //o
    .PE_OUT    (pE_538_PE_OUT[31:0]             ), //o
    .finish    (pE_538_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_539 (
    .activate  (pE_530_acount[7:0]              ), //i
    .weight    (pE_530_bcount[7:0]              ), //i
    .valid     (pE_539_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_539_acount[7:0]              ), //o
    .bcount    (pE_539_bcount[7:0]              ), //o
    .PE_OUT    (pE_539_PE_OUT[31:0]             ), //o
    .finish    (pE_539_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_540 (
    .activate  (pE_531_acount[7:0]              ), //i
    .weight    (pE_531_bcount[7:0]              ), //i
    .valid     (pE_540_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_540_acount[7:0]              ), //o
    .bcount    (pE_540_bcount[7:0]              ), //o
    .PE_OUT    (pE_540_PE_OUT[31:0]             ), //o
    .finish    (pE_540_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_541 (
    .activate  (pE_532_acount[7:0]              ), //i
    .weight    (pE_532_bcount[7:0]              ), //i
    .valid     (pE_541_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_541_acount[7:0]              ), //o
    .bcount    (pE_541_bcount[7:0]              ), //o
    .PE_OUT    (pE_541_PE_OUT[31:0]             ), //o
    .finish    (pE_541_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_542 (
    .activate  (pE_533_acount[7:0]              ), //i
    .weight    (pE_533_bcount[7:0]              ), //i
    .valid     (pE_542_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_542_acount[7:0]              ), //o
    .bcount    (pE_542_bcount[7:0]              ), //o
    .PE_OUT    (pE_542_PE_OUT[31:0]             ), //o
    .finish    (pE_542_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_543 (
    .activate  (pE_534_acount[7:0]              ), //i
    .weight    (pE_534_bcount[7:0]              ), //i
    .valid     (pE_543_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_543_acount[7:0]              ), //o
    .bcount    (pE_543_bcount[7:0]              ), //o
    .PE_OUT    (pE_543_PE_OUT[31:0]             ), //o
    .finish    (pE_543_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_544 (
    .activate  (pE_544_acount[7:0]              ), //i
    .weight    (pE_536_bcount[7:0]              ), //i
    .valid     (pE_544_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_544_acount[7:0]              ), //o
    .bcount    (pE_544_bcount[7:0]              ), //o
    .PE_OUT    (pE_544_PE_OUT[31:0]             ), //o
    .finish    (pE_544_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_545 (
    .activate  (pE_536_acount[7:0]              ), //i
    .weight    (pE_536_bcount[7:0]              ), //i
    .valid     (pE_545_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_545_acount[7:0]              ), //o
    .bcount    (pE_545_bcount[7:0]              ), //o
    .PE_OUT    (pE_545_PE_OUT[31:0]             ), //o
    .finish    (pE_545_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_546 (
    .activate  (pE_537_acount[7:0]              ), //i
    .weight    (pE_537_bcount[7:0]              ), //i
    .valid     (pE_546_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_546_acount[7:0]              ), //o
    .bcount    (pE_546_bcount[7:0]              ), //o
    .PE_OUT    (pE_546_PE_OUT[31:0]             ), //o
    .finish    (pE_546_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_547 (
    .activate  (pE_538_acount[7:0]              ), //i
    .weight    (pE_538_bcount[7:0]              ), //i
    .valid     (pE_547_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_547_acount[7:0]              ), //o
    .bcount    (pE_547_bcount[7:0]              ), //o
    .PE_OUT    (pE_547_PE_OUT[31:0]             ), //o
    .finish    (pE_547_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_548 (
    .activate  (pE_539_acount[7:0]              ), //i
    .weight    (pE_539_bcount[7:0]              ), //i
    .valid     (pE_548_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_548_acount[7:0]              ), //o
    .bcount    (pE_548_bcount[7:0]              ), //o
    .PE_OUT    (pE_548_PE_OUT[31:0]             ), //o
    .finish    (pE_548_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_549 (
    .activate  (pE_540_acount[7:0]              ), //i
    .weight    (pE_540_bcount[7:0]              ), //i
    .valid     (pE_549_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_549_acount[7:0]              ), //o
    .bcount    (pE_549_bcount[7:0]              ), //o
    .PE_OUT    (pE_549_PE_OUT[31:0]             ), //o
    .finish    (pE_549_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_550 (
    .activate  (pE_541_acount[7:0]              ), //i
    .weight    (pE_541_bcount[7:0]              ), //i
    .valid     (pE_550_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_550_acount[7:0]              ), //o
    .bcount    (pE_550_bcount[7:0]              ), //o
    .PE_OUT    (pE_550_PE_OUT[31:0]             ), //o
    .finish    (pE_550_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_551 (
    .activate  (pE_542_acount[7:0]              ), //i
    .weight    (pE_542_bcount[7:0]              ), //i
    .valid     (pE_551_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_551_acount[7:0]              ), //o
    .bcount    (pE_551_bcount[7:0]              ), //o
    .PE_OUT    (pE_551_PE_OUT[31:0]             ), //o
    .finish    (pE_551_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_552 (
    .activate  (pE_552_acount[7:0]              ), //i
    .weight    (pE_544_bcount[7:0]              ), //i
    .valid     (pE_552_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_552_acount[7:0]              ), //o
    .bcount    (pE_552_bcount[7:0]              ), //o
    .PE_OUT    (pE_552_PE_OUT[31:0]             ), //o
    .finish    (pE_552_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_553 (
    .activate  (pE_544_acount[7:0]              ), //i
    .weight    (pE_544_bcount[7:0]              ), //i
    .valid     (pE_553_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_553_acount[7:0]              ), //o
    .bcount    (pE_553_bcount[7:0]              ), //o
    .PE_OUT    (pE_553_PE_OUT[31:0]             ), //o
    .finish    (pE_553_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_554 (
    .activate  (pE_545_acount[7:0]              ), //i
    .weight    (pE_545_bcount[7:0]              ), //i
    .valid     (pE_554_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_554_acount[7:0]              ), //o
    .bcount    (pE_554_bcount[7:0]              ), //o
    .PE_OUT    (pE_554_PE_OUT[31:0]             ), //o
    .finish    (pE_554_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_555 (
    .activate  (pE_546_acount[7:0]              ), //i
    .weight    (pE_546_bcount[7:0]              ), //i
    .valid     (pE_555_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_555_acount[7:0]              ), //o
    .bcount    (pE_555_bcount[7:0]              ), //o
    .PE_OUT    (pE_555_PE_OUT[31:0]             ), //o
    .finish    (pE_555_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_556 (
    .activate  (pE_547_acount[7:0]              ), //i
    .weight    (pE_547_bcount[7:0]              ), //i
    .valid     (pE_556_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_556_acount[7:0]              ), //o
    .bcount    (pE_556_bcount[7:0]              ), //o
    .PE_OUT    (pE_556_PE_OUT[31:0]             ), //o
    .finish    (pE_556_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_557 (
    .activate  (pE_548_acount[7:0]              ), //i
    .weight    (pE_548_bcount[7:0]              ), //i
    .valid     (pE_557_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_557_acount[7:0]              ), //o
    .bcount    (pE_557_bcount[7:0]              ), //o
    .PE_OUT    (pE_557_PE_OUT[31:0]             ), //o
    .finish    (pE_557_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_558 (
    .activate  (pE_549_acount[7:0]              ), //i
    .weight    (pE_549_bcount[7:0]              ), //i
    .valid     (pE_558_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_558_acount[7:0]              ), //o
    .bcount    (pE_558_bcount[7:0]              ), //o
    .PE_OUT    (pE_558_PE_OUT[31:0]             ), //o
    .finish    (pE_558_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_559 (
    .activate  (pE_550_acount[7:0]              ), //i
    .weight    (pE_550_bcount[7:0]              ), //i
    .valid     (pE_559_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_559_acount[7:0]              ), //o
    .bcount    (pE_559_bcount[7:0]              ), //o
    .PE_OUT    (pE_559_PE_OUT[31:0]             ), //o
    .finish    (pE_559_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_560 (
    .activate  (pE_560_acount[7:0]              ), //i
    .weight    (pE_552_bcount[7:0]              ), //i
    .valid     (pE_560_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_560_acount[7:0]              ), //o
    .bcount    (pE_560_bcount[7:0]              ), //o
    .PE_OUT    (pE_560_PE_OUT[31:0]             ), //o
    .finish    (pE_560_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_561 (
    .activate  (pE_552_acount[7:0]              ), //i
    .weight    (pE_552_bcount[7:0]              ), //i
    .valid     (pE_561_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_561_acount[7:0]              ), //o
    .bcount    (pE_561_bcount[7:0]              ), //o
    .PE_OUT    (pE_561_PE_OUT[31:0]             ), //o
    .finish    (pE_561_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_562 (
    .activate  (pE_553_acount[7:0]              ), //i
    .weight    (pE_553_bcount[7:0]              ), //i
    .valid     (pE_562_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_562_acount[7:0]              ), //o
    .bcount    (pE_562_bcount[7:0]              ), //o
    .PE_OUT    (pE_562_PE_OUT[31:0]             ), //o
    .finish    (pE_562_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_563 (
    .activate  (pE_554_acount[7:0]              ), //i
    .weight    (pE_554_bcount[7:0]              ), //i
    .valid     (pE_563_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_563_acount[7:0]              ), //o
    .bcount    (pE_563_bcount[7:0]              ), //o
    .PE_OUT    (pE_563_PE_OUT[31:0]             ), //o
    .finish    (pE_563_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_564 (
    .activate  (pE_555_acount[7:0]              ), //i
    .weight    (pE_555_bcount[7:0]              ), //i
    .valid     (pE_564_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_564_acount[7:0]              ), //o
    .bcount    (pE_564_bcount[7:0]              ), //o
    .PE_OUT    (pE_564_PE_OUT[31:0]             ), //o
    .finish    (pE_564_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_565 (
    .activate  (pE_556_acount[7:0]              ), //i
    .weight    (pE_556_bcount[7:0]              ), //i
    .valid     (pE_565_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_565_acount[7:0]              ), //o
    .bcount    (pE_565_bcount[7:0]              ), //o
    .PE_OUT    (pE_565_PE_OUT[31:0]             ), //o
    .finish    (pE_565_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_566 (
    .activate  (pE_557_acount[7:0]              ), //i
    .weight    (pE_557_bcount[7:0]              ), //i
    .valid     (pE_566_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_566_acount[7:0]              ), //o
    .bcount    (pE_566_bcount[7:0]              ), //o
    .PE_OUT    (pE_566_PE_OUT[31:0]             ), //o
    .finish    (pE_566_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_567 (
    .activate  (pE_558_acount[7:0]              ), //i
    .weight    (pE_558_bcount[7:0]              ), //i
    .valid     (pE_567_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_567_acount[7:0]              ), //o
    .bcount    (pE_567_bcount[7:0]              ), //o
    .PE_OUT    (pE_567_PE_OUT[31:0]             ), //o
    .finish    (pE_567_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_568 (
    .activate  (pE_568_acount[7:0]              ), //i
    .weight    (pE_560_bcount[7:0]              ), //i
    .valid     (pE_568_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_568_acount[7:0]              ), //o
    .bcount    (pE_568_bcount[7:0]              ), //o
    .PE_OUT    (pE_568_PE_OUT[31:0]             ), //o
    .finish    (pE_568_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_569 (
    .activate  (pE_560_acount[7:0]              ), //i
    .weight    (pE_560_bcount[7:0]              ), //i
    .valid     (pE_569_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_569_acount[7:0]              ), //o
    .bcount    (pE_569_bcount[7:0]              ), //o
    .PE_OUT    (pE_569_PE_OUT[31:0]             ), //o
    .finish    (pE_569_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_570 (
    .activate  (pE_561_acount[7:0]              ), //i
    .weight    (pE_561_bcount[7:0]              ), //i
    .valid     (pE_570_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_570_acount[7:0]              ), //o
    .bcount    (pE_570_bcount[7:0]              ), //o
    .PE_OUT    (pE_570_PE_OUT[31:0]             ), //o
    .finish    (pE_570_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_571 (
    .activate  (pE_562_acount[7:0]              ), //i
    .weight    (pE_562_bcount[7:0]              ), //i
    .valid     (pE_571_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_571_acount[7:0]              ), //o
    .bcount    (pE_571_bcount[7:0]              ), //o
    .PE_OUT    (pE_571_PE_OUT[31:0]             ), //o
    .finish    (pE_571_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_572 (
    .activate  (pE_563_acount[7:0]              ), //i
    .weight    (pE_563_bcount[7:0]              ), //i
    .valid     (pE_572_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_572_acount[7:0]              ), //o
    .bcount    (pE_572_bcount[7:0]              ), //o
    .PE_OUT    (pE_572_PE_OUT[31:0]             ), //o
    .finish    (pE_572_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_573 (
    .activate  (pE_564_acount[7:0]              ), //i
    .weight    (pE_564_bcount[7:0]              ), //i
    .valid     (pE_573_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_573_acount[7:0]              ), //o
    .bcount    (pE_573_bcount[7:0]              ), //o
    .PE_OUT    (pE_573_PE_OUT[31:0]             ), //o
    .finish    (pE_573_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_574 (
    .activate  (pE_565_acount[7:0]              ), //i
    .weight    (pE_565_bcount[7:0]              ), //i
    .valid     (pE_574_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_574_acount[7:0]              ), //o
    .bcount    (pE_574_bcount[7:0]              ), //o
    .PE_OUT    (pE_574_PE_OUT[31:0]             ), //o
    .finish    (pE_574_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_575 (
    .activate  (pE_566_acount[7:0]              ), //i
    .weight    (pE_566_bcount[7:0]              ), //i
    .valid     (pE_575_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_575_acount[7:0]              ), //o
    .bcount    (pE_575_bcount[7:0]              ), //o
    .PE_OUT    (pE_575_PE_OUT[31:0]             ), //o
    .finish    (pE_575_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  always @(*) begin
    MatrixC_0 = 32'h0;
    if(when_SA_3D_l80) begin
      MatrixC_0 = pE_512_PE_OUT;
    end
    if(when_SA_3D_l80_1) begin
      MatrixC_0 = pE_513_PE_OUT;
    end
    if(when_SA_3D_l80_2) begin
      MatrixC_0 = pE_514_PE_OUT;
    end
    if(when_SA_3D_l80_3) begin
      MatrixC_0 = pE_515_PE_OUT;
    end
    if(when_SA_3D_l80_4) begin
      MatrixC_0 = pE_516_PE_OUT;
    end
    if(when_SA_3D_l80_5) begin
      MatrixC_0 = pE_517_PE_OUT;
    end
    if(when_SA_3D_l80_6) begin
      MatrixC_0 = pE_518_PE_OUT;
    end
    if(when_SA_3D_l80_7) begin
      MatrixC_0 = pE_519_PE_OUT;
    end
  end

  always @(*) begin
    tmp[0] = pE_512_valid;
    tmp[0] = pE_513_valid;
    tmp[0] = pE_514_valid;
    tmp[0] = pE_515_valid;
    tmp[0] = pE_516_valid;
    tmp[0] = pE_517_valid;
    tmp[0] = pE_518_valid;
    tmp[0] = pE_519_valid;
    tmp[1] = pE_520_valid;
    tmp[1] = pE_521_valid;
    tmp[1] = pE_522_valid;
    tmp[1] = pE_523_valid;
    tmp[1] = pE_524_valid;
    tmp[1] = pE_525_valid;
    tmp[1] = pE_526_valid;
    tmp[1] = pE_527_valid;
    tmp[2] = pE_528_valid;
    tmp[2] = pE_529_valid;
    tmp[2] = pE_530_valid;
    tmp[2] = pE_531_valid;
    tmp[2] = pE_532_valid;
    tmp[2] = pE_533_valid;
    tmp[2] = pE_534_valid;
    tmp[2] = pE_535_valid;
    tmp[3] = pE_536_valid;
    tmp[3] = pE_537_valid;
    tmp[3] = pE_538_valid;
    tmp[3] = pE_539_valid;
    tmp[3] = pE_540_valid;
    tmp[3] = pE_541_valid;
    tmp[3] = pE_542_valid;
    tmp[3] = pE_543_valid;
    tmp[4] = pE_544_valid;
    tmp[4] = pE_545_valid;
    tmp[4] = pE_546_valid;
    tmp[4] = pE_547_valid;
    tmp[4] = pE_548_valid;
    tmp[4] = pE_549_valid;
    tmp[4] = pE_550_valid;
    tmp[4] = pE_551_valid;
    tmp[5] = pE_552_valid;
    tmp[5] = pE_553_valid;
    tmp[5] = pE_554_valid;
    tmp[5] = pE_555_valid;
    tmp[5] = pE_556_valid;
    tmp[5] = pE_557_valid;
    tmp[5] = pE_558_valid;
    tmp[5] = pE_559_valid;
    tmp[6] = pE_560_valid;
    tmp[6] = pE_561_valid;
    tmp[6] = pE_562_valid;
    tmp[6] = pE_563_valid;
    tmp[6] = pE_564_valid;
    tmp[6] = pE_565_valid;
    tmp[6] = pE_566_valid;
    tmp[6] = pE_567_valid;
    tmp[7] = pE_568_valid;
    tmp[7] = pE_569_valid;
    tmp[7] = pE_570_valid;
    tmp[7] = pE_571_valid;
    tmp[7] = pE_572_valid;
    tmp[7] = pE_573_valid;
    tmp[7] = pE_574_valid;
    tmp[7] = pE_575_valid;
  end

  assign when_SA_3D_l80 = tmp[0];
  assign when_SA_3D_l80_1 = tmp[1];
  assign when_SA_3D_l80_2 = tmp[2];
  assign when_SA_3D_l80_3 = tmp[3];
  assign when_SA_3D_l80_4 = tmp[4];
  assign when_SA_3D_l80_5 = tmp[5];
  assign when_SA_3D_l80_6 = tmp[6];
  assign when_SA_3D_l80_7 = tmp[7];
  assign C_Valid_0 = (|tmp);
  always @(*) begin
    MatrixC_1 = 32'h0;
    if(when_SA_3D_l80_8) begin
      MatrixC_1 = pE_520_PE_OUT;
    end
    if(when_SA_3D_l80_9) begin
      MatrixC_1 = pE_521_PE_OUT;
    end
    if(when_SA_3D_l80_10) begin
      MatrixC_1 = pE_522_PE_OUT;
    end
    if(when_SA_3D_l80_11) begin
      MatrixC_1 = pE_523_PE_OUT;
    end
    if(when_SA_3D_l80_12) begin
      MatrixC_1 = pE_524_PE_OUT;
    end
    if(when_SA_3D_l80_13) begin
      MatrixC_1 = pE_525_PE_OUT;
    end
    if(when_SA_3D_l80_14) begin
      MatrixC_1 = pE_526_PE_OUT;
    end
    if(when_SA_3D_l80_15) begin
      MatrixC_1 = pE_527_PE_OUT;
    end
  end

  assign when_SA_3D_l80_8 = tmp[0];
  assign when_SA_3D_l80_9 = tmp[1];
  assign when_SA_3D_l80_10 = tmp[2];
  assign when_SA_3D_l80_11 = tmp[3];
  assign when_SA_3D_l80_12 = tmp[4];
  assign when_SA_3D_l80_13 = tmp[5];
  assign when_SA_3D_l80_14 = tmp[6];
  assign when_SA_3D_l80_15 = tmp[7];
  assign C_Valid_1 = (|tmp);
  always @(*) begin
    MatrixC_2 = 32'h0;
    if(when_SA_3D_l80_16) begin
      MatrixC_2 = pE_528_PE_OUT;
    end
    if(when_SA_3D_l80_17) begin
      MatrixC_2 = pE_529_PE_OUT;
    end
    if(when_SA_3D_l80_18) begin
      MatrixC_2 = pE_530_PE_OUT;
    end
    if(when_SA_3D_l80_19) begin
      MatrixC_2 = pE_531_PE_OUT;
    end
    if(when_SA_3D_l80_20) begin
      MatrixC_2 = pE_532_PE_OUT;
    end
    if(when_SA_3D_l80_21) begin
      MatrixC_2 = pE_533_PE_OUT;
    end
    if(when_SA_3D_l80_22) begin
      MatrixC_2 = pE_534_PE_OUT;
    end
    if(when_SA_3D_l80_23) begin
      MatrixC_2 = pE_535_PE_OUT;
    end
  end

  assign when_SA_3D_l80_16 = tmp[0];
  assign when_SA_3D_l80_17 = tmp[1];
  assign when_SA_3D_l80_18 = tmp[2];
  assign when_SA_3D_l80_19 = tmp[3];
  assign when_SA_3D_l80_20 = tmp[4];
  assign when_SA_3D_l80_21 = tmp[5];
  assign when_SA_3D_l80_22 = tmp[6];
  assign when_SA_3D_l80_23 = tmp[7];
  assign C_Valid_2 = (|tmp);
  always @(*) begin
    MatrixC_3 = 32'h0;
    if(when_SA_3D_l80_24) begin
      MatrixC_3 = pE_536_PE_OUT;
    end
    if(when_SA_3D_l80_25) begin
      MatrixC_3 = pE_537_PE_OUT;
    end
    if(when_SA_3D_l80_26) begin
      MatrixC_3 = pE_538_PE_OUT;
    end
    if(when_SA_3D_l80_27) begin
      MatrixC_3 = pE_539_PE_OUT;
    end
    if(when_SA_3D_l80_28) begin
      MatrixC_3 = pE_540_PE_OUT;
    end
    if(when_SA_3D_l80_29) begin
      MatrixC_3 = pE_541_PE_OUT;
    end
    if(when_SA_3D_l80_30) begin
      MatrixC_3 = pE_542_PE_OUT;
    end
    if(when_SA_3D_l80_31) begin
      MatrixC_3 = pE_543_PE_OUT;
    end
  end

  assign when_SA_3D_l80_24 = tmp[0];
  assign when_SA_3D_l80_25 = tmp[1];
  assign when_SA_3D_l80_26 = tmp[2];
  assign when_SA_3D_l80_27 = tmp[3];
  assign when_SA_3D_l80_28 = tmp[4];
  assign when_SA_3D_l80_29 = tmp[5];
  assign when_SA_3D_l80_30 = tmp[6];
  assign when_SA_3D_l80_31 = tmp[7];
  assign C_Valid_3 = (|tmp);
  always @(*) begin
    MatrixC_4 = 32'h0;
    if(when_SA_3D_l80_32) begin
      MatrixC_4 = pE_544_PE_OUT;
    end
    if(when_SA_3D_l80_33) begin
      MatrixC_4 = pE_545_PE_OUT;
    end
    if(when_SA_3D_l80_34) begin
      MatrixC_4 = pE_546_PE_OUT;
    end
    if(when_SA_3D_l80_35) begin
      MatrixC_4 = pE_547_PE_OUT;
    end
    if(when_SA_3D_l80_36) begin
      MatrixC_4 = pE_548_PE_OUT;
    end
    if(when_SA_3D_l80_37) begin
      MatrixC_4 = pE_549_PE_OUT;
    end
    if(when_SA_3D_l80_38) begin
      MatrixC_4 = pE_550_PE_OUT;
    end
    if(when_SA_3D_l80_39) begin
      MatrixC_4 = pE_551_PE_OUT;
    end
  end

  assign when_SA_3D_l80_32 = tmp[0];
  assign when_SA_3D_l80_33 = tmp[1];
  assign when_SA_3D_l80_34 = tmp[2];
  assign when_SA_3D_l80_35 = tmp[3];
  assign when_SA_3D_l80_36 = tmp[4];
  assign when_SA_3D_l80_37 = tmp[5];
  assign when_SA_3D_l80_38 = tmp[6];
  assign when_SA_3D_l80_39 = tmp[7];
  assign C_Valid_4 = (|tmp);
  always @(*) begin
    MatrixC_5 = 32'h0;
    if(when_SA_3D_l80_40) begin
      MatrixC_5 = pE_552_PE_OUT;
    end
    if(when_SA_3D_l80_41) begin
      MatrixC_5 = pE_553_PE_OUT;
    end
    if(when_SA_3D_l80_42) begin
      MatrixC_5 = pE_554_PE_OUT;
    end
    if(when_SA_3D_l80_43) begin
      MatrixC_5 = pE_555_PE_OUT;
    end
    if(when_SA_3D_l80_44) begin
      MatrixC_5 = pE_556_PE_OUT;
    end
    if(when_SA_3D_l80_45) begin
      MatrixC_5 = pE_557_PE_OUT;
    end
    if(when_SA_3D_l80_46) begin
      MatrixC_5 = pE_558_PE_OUT;
    end
    if(when_SA_3D_l80_47) begin
      MatrixC_5 = pE_559_PE_OUT;
    end
  end

  assign when_SA_3D_l80_40 = tmp[0];
  assign when_SA_3D_l80_41 = tmp[1];
  assign when_SA_3D_l80_42 = tmp[2];
  assign when_SA_3D_l80_43 = tmp[3];
  assign when_SA_3D_l80_44 = tmp[4];
  assign when_SA_3D_l80_45 = tmp[5];
  assign when_SA_3D_l80_46 = tmp[6];
  assign when_SA_3D_l80_47 = tmp[7];
  assign C_Valid_5 = (|tmp);
  always @(*) begin
    MatrixC_6 = 32'h0;
    if(when_SA_3D_l80_48) begin
      MatrixC_6 = pE_560_PE_OUT;
    end
    if(when_SA_3D_l80_49) begin
      MatrixC_6 = pE_561_PE_OUT;
    end
    if(when_SA_3D_l80_50) begin
      MatrixC_6 = pE_562_PE_OUT;
    end
    if(when_SA_3D_l80_51) begin
      MatrixC_6 = pE_563_PE_OUT;
    end
    if(when_SA_3D_l80_52) begin
      MatrixC_6 = pE_564_PE_OUT;
    end
    if(when_SA_3D_l80_53) begin
      MatrixC_6 = pE_565_PE_OUT;
    end
    if(when_SA_3D_l80_54) begin
      MatrixC_6 = pE_566_PE_OUT;
    end
    if(when_SA_3D_l80_55) begin
      MatrixC_6 = pE_567_PE_OUT;
    end
  end

  assign when_SA_3D_l80_48 = tmp[0];
  assign when_SA_3D_l80_49 = tmp[1];
  assign when_SA_3D_l80_50 = tmp[2];
  assign when_SA_3D_l80_51 = tmp[3];
  assign when_SA_3D_l80_52 = tmp[4];
  assign when_SA_3D_l80_53 = tmp[5];
  assign when_SA_3D_l80_54 = tmp[6];
  assign when_SA_3D_l80_55 = tmp[7];
  assign C_Valid_6 = (|tmp);
  always @(*) begin
    MatrixC_7 = 32'h0;
    if(when_SA_3D_l80_56) begin
      MatrixC_7 = pE_568_PE_OUT;
    end
    if(when_SA_3D_l80_57) begin
      MatrixC_7 = pE_569_PE_OUT;
    end
    if(when_SA_3D_l80_58) begin
      MatrixC_7 = pE_570_PE_OUT;
    end
    if(when_SA_3D_l80_59) begin
      MatrixC_7 = pE_571_PE_OUT;
    end
    if(when_SA_3D_l80_60) begin
      MatrixC_7 = pE_572_PE_OUT;
    end
    if(when_SA_3D_l80_61) begin
      MatrixC_7 = pE_573_PE_OUT;
    end
    if(when_SA_3D_l80_62) begin
      MatrixC_7 = pE_574_PE_OUT;
    end
    if(when_SA_3D_l80_63) begin
      MatrixC_7 = pE_575_PE_OUT;
    end
  end

  assign when_SA_3D_l80_56 = tmp[0];
  assign when_SA_3D_l80_57 = tmp[1];
  assign when_SA_3D_l80_58 = tmp[2];
  assign when_SA_3D_l80_59 = tmp[3];
  assign when_SA_3D_l80_60 = tmp[4];
  assign when_SA_3D_l80_61 = tmp[5];
  assign when_SA_3D_l80_62 = tmp[6];
  assign when_SA_3D_l80_63 = tmp[7];
  assign C_Valid_7 = (|tmp);
  assign pE_512_valid = (io_A_Valid_0 && io_B_Valid_0);
  assign pE_513_valid = (io_A_Valid_0_delay_1 && io_B_Valid_1);
  assign pE_514_valid = (io_A_Valid_0_delay_2 && io_B_Valid_2);
  assign pE_515_valid = (io_A_Valid_0_delay_3 && io_B_Valid_3);
  assign pE_516_valid = (io_A_Valid_0_delay_4 && io_B_Valid_4);
  assign pE_517_valid = (io_A_Valid_0_delay_5 && io_B_Valid_5);
  assign pE_518_valid = (io_A_Valid_0_delay_6 && io_B_Valid_6);
  assign pE_519_valid = (io_A_Valid_0_delay_7 && io_B_Valid_7);
  assign pE_520_valid = (io_A_Valid_1 && io_B_Valid_0_delay_1);
  assign pE_521_valid = (io_A_Valid_1_delay_1 && io_B_Valid_1_delay_1);
  assign pE_522_valid = (io_A_Valid_1_delay_2 && io_B_Valid_2_delay_1);
  assign pE_523_valid = (io_A_Valid_1_delay_3 && io_B_Valid_3_delay_1);
  assign pE_524_valid = (io_A_Valid_1_delay_4 && io_B_Valid_4_delay_1);
  assign pE_525_valid = (io_A_Valid_1_delay_5 && io_B_Valid_5_delay_1);
  assign pE_526_valid = (io_A_Valid_1_delay_6 && io_B_Valid_6_delay_1);
  assign pE_527_valid = (io_A_Valid_1_delay_7 && io_B_Valid_7_delay_1);
  assign pE_528_valid = (io_A_Valid_2 && io_B_Valid_0_delay_2);
  assign pE_529_valid = (io_A_Valid_2_delay_1 && io_B_Valid_1_delay_2);
  assign pE_530_valid = (io_A_Valid_2_delay_2 && io_B_Valid_2_delay_2);
  assign pE_531_valid = (io_A_Valid_2_delay_3 && io_B_Valid_3_delay_2);
  assign pE_532_valid = (io_A_Valid_2_delay_4 && io_B_Valid_4_delay_2);
  assign pE_533_valid = (io_A_Valid_2_delay_5 && io_B_Valid_5_delay_2);
  assign pE_534_valid = (io_A_Valid_2_delay_6 && io_B_Valid_6_delay_2);
  assign pE_535_valid = (io_A_Valid_2_delay_7 && io_B_Valid_7_delay_2);
  assign pE_536_valid = (io_A_Valid_3 && io_B_Valid_0_delay_3);
  assign pE_537_valid = (io_A_Valid_3_delay_1 && io_B_Valid_1_delay_3);
  assign pE_538_valid = (io_A_Valid_3_delay_2 && io_B_Valid_2_delay_3);
  assign pE_539_valid = (io_A_Valid_3_delay_3 && io_B_Valid_3_delay_3);
  assign pE_540_valid = (io_A_Valid_3_delay_4 && io_B_Valid_4_delay_3);
  assign pE_541_valid = (io_A_Valid_3_delay_5 && io_B_Valid_5_delay_3);
  assign pE_542_valid = (io_A_Valid_3_delay_6 && io_B_Valid_6_delay_3);
  assign pE_543_valid = (io_A_Valid_3_delay_7 && io_B_Valid_7_delay_3);
  assign pE_544_valid = (io_A_Valid_4 && io_B_Valid_0_delay_4);
  assign pE_545_valid = (io_A_Valid_4_delay_1 && io_B_Valid_1_delay_4);
  assign pE_546_valid = (io_A_Valid_4_delay_2 && io_B_Valid_2_delay_4);
  assign pE_547_valid = (io_A_Valid_4_delay_3 && io_B_Valid_3_delay_4);
  assign pE_548_valid = (io_A_Valid_4_delay_4 && io_B_Valid_4_delay_4);
  assign pE_549_valid = (io_A_Valid_4_delay_5 && io_B_Valid_5_delay_4);
  assign pE_550_valid = (io_A_Valid_4_delay_6 && io_B_Valid_6_delay_4);
  assign pE_551_valid = (io_A_Valid_4_delay_7 && io_B_Valid_7_delay_4);
  assign pE_552_valid = (io_A_Valid_5 && io_B_Valid_0_delay_5);
  assign pE_553_valid = (io_A_Valid_5_delay_1 && io_B_Valid_1_delay_5);
  assign pE_554_valid = (io_A_Valid_5_delay_2 && io_B_Valid_2_delay_5);
  assign pE_555_valid = (io_A_Valid_5_delay_3 && io_B_Valid_3_delay_5);
  assign pE_556_valid = (io_A_Valid_5_delay_4 && io_B_Valid_4_delay_5);
  assign pE_557_valid = (io_A_Valid_5_delay_5 && io_B_Valid_5_delay_5);
  assign pE_558_valid = (io_A_Valid_5_delay_6 && io_B_Valid_6_delay_5);
  assign pE_559_valid = (io_A_Valid_5_delay_7 && io_B_Valid_7_delay_5);
  assign pE_560_valid = (io_A_Valid_6 && io_B_Valid_0_delay_6);
  assign pE_561_valid = (io_A_Valid_6_delay_1 && io_B_Valid_1_delay_6);
  assign pE_562_valid = (io_A_Valid_6_delay_2 && io_B_Valid_2_delay_6);
  assign pE_563_valid = (io_A_Valid_6_delay_3 && io_B_Valid_3_delay_6);
  assign pE_564_valid = (io_A_Valid_6_delay_4 && io_B_Valid_4_delay_6);
  assign pE_565_valid = (io_A_Valid_6_delay_5 && io_B_Valid_5_delay_6);
  assign pE_566_valid = (io_A_Valid_6_delay_6 && io_B_Valid_6_delay_6);
  assign pE_567_valid = (io_A_Valid_6_delay_7 && io_B_Valid_7_delay_6);
  assign pE_568_valid = (io_A_Valid_7 && io_B_Valid_0_delay_7);
  assign pE_569_valid = (io_A_Valid_7_delay_1 && io_B_Valid_1_delay_7);
  assign pE_570_valid = (io_A_Valid_7_delay_2 && io_B_Valid_2_delay_7);
  assign pE_571_valid = (io_A_Valid_7_delay_3 && io_B_Valid_3_delay_7);
  assign pE_572_valid = (io_A_Valid_7_delay_4 && io_B_Valid_4_delay_7);
  assign pE_573_valid = (io_A_Valid_7_delay_5 && io_B_Valid_5_delay_7);
  assign pE_574_valid = (io_A_Valid_7_delay_6 && io_B_Valid_6_delay_7);
  assign pE_575_valid = (io_A_Valid_7_delay_7 && io_B_Valid_7_delay_7);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      io_signCount_regNextWhen <= 16'h0;
      io_signCount_regNextWhen_1 <= 16'h0;
      io_signCount_regNextWhen_2 <= 16'h0;
      io_signCount_regNextWhen_3 <= 16'h0;
      io_signCount_regNextWhen_4 <= 16'h0;
      io_signCount_regNextWhen_5 <= 16'h0;
      io_signCount_regNextWhen_6 <= 16'h0;
      io_signCount_regNextWhen_7 <= 16'h0;
    end else begin
      if(start) begin
        io_signCount_regNextWhen <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_1 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_2 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_3 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_4 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_5 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_6 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_7 <= io_signCount;
      end
    end
  end

  always @(posedge clk) begin
    io_A_Valid_0_delay_1 <= io_A_Valid_0;
    io_A_Valid_0_delay_1_1 <= io_A_Valid_0;
    io_A_Valid_0_delay_2 <= io_A_Valid_0_delay_1_1;
    io_A_Valid_0_delay_1_2 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_1 <= io_A_Valid_0_delay_1_2;
    io_A_Valid_0_delay_3 <= io_A_Valid_0_delay_2_1;
    io_A_Valid_0_delay_1_3 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_2 <= io_A_Valid_0_delay_1_3;
    io_A_Valid_0_delay_3_1 <= io_A_Valid_0_delay_2_2;
    io_A_Valid_0_delay_4 <= io_A_Valid_0_delay_3_1;
    io_A_Valid_0_delay_1_4 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_3 <= io_A_Valid_0_delay_1_4;
    io_A_Valid_0_delay_3_2 <= io_A_Valid_0_delay_2_3;
    io_A_Valid_0_delay_4_1 <= io_A_Valid_0_delay_3_2;
    io_A_Valid_0_delay_5 <= io_A_Valid_0_delay_4_1;
    io_A_Valid_0_delay_1_5 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_4 <= io_A_Valid_0_delay_1_5;
    io_A_Valid_0_delay_3_3 <= io_A_Valid_0_delay_2_4;
    io_A_Valid_0_delay_4_2 <= io_A_Valid_0_delay_3_3;
    io_A_Valid_0_delay_5_1 <= io_A_Valid_0_delay_4_2;
    io_A_Valid_0_delay_6 <= io_A_Valid_0_delay_5_1;
    io_A_Valid_0_delay_1_6 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_5 <= io_A_Valid_0_delay_1_6;
    io_A_Valid_0_delay_3_4 <= io_A_Valid_0_delay_2_5;
    io_A_Valid_0_delay_4_3 <= io_A_Valid_0_delay_3_4;
    io_A_Valid_0_delay_5_2 <= io_A_Valid_0_delay_4_3;
    io_A_Valid_0_delay_6_1 <= io_A_Valid_0_delay_5_2;
    io_A_Valid_0_delay_7 <= io_A_Valid_0_delay_6_1;
    io_B_Valid_0_delay_1 <= io_B_Valid_0;
    io_A_Valid_1_delay_1 <= io_A_Valid_1;
    io_B_Valid_1_delay_1 <= io_B_Valid_1;
    io_A_Valid_1_delay_1_1 <= io_A_Valid_1;
    io_A_Valid_1_delay_2 <= io_A_Valid_1_delay_1_1;
    io_B_Valid_2_delay_1 <= io_B_Valid_2;
    io_A_Valid_1_delay_1_2 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_1 <= io_A_Valid_1_delay_1_2;
    io_A_Valid_1_delay_3 <= io_A_Valid_1_delay_2_1;
    io_B_Valid_3_delay_1 <= io_B_Valid_3;
    io_A_Valid_1_delay_1_3 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_2 <= io_A_Valid_1_delay_1_3;
    io_A_Valid_1_delay_3_1 <= io_A_Valid_1_delay_2_2;
    io_A_Valid_1_delay_4 <= io_A_Valid_1_delay_3_1;
    io_B_Valid_4_delay_1 <= io_B_Valid_4;
    io_A_Valid_1_delay_1_4 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_3 <= io_A_Valid_1_delay_1_4;
    io_A_Valid_1_delay_3_2 <= io_A_Valid_1_delay_2_3;
    io_A_Valid_1_delay_4_1 <= io_A_Valid_1_delay_3_2;
    io_A_Valid_1_delay_5 <= io_A_Valid_1_delay_4_1;
    io_B_Valid_5_delay_1 <= io_B_Valid_5;
    io_A_Valid_1_delay_1_5 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_4 <= io_A_Valid_1_delay_1_5;
    io_A_Valid_1_delay_3_3 <= io_A_Valid_1_delay_2_4;
    io_A_Valid_1_delay_4_2 <= io_A_Valid_1_delay_3_3;
    io_A_Valid_1_delay_5_1 <= io_A_Valid_1_delay_4_2;
    io_A_Valid_1_delay_6 <= io_A_Valid_1_delay_5_1;
    io_B_Valid_6_delay_1 <= io_B_Valid_6;
    io_A_Valid_1_delay_1_6 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_5 <= io_A_Valid_1_delay_1_6;
    io_A_Valid_1_delay_3_4 <= io_A_Valid_1_delay_2_5;
    io_A_Valid_1_delay_4_3 <= io_A_Valid_1_delay_3_4;
    io_A_Valid_1_delay_5_2 <= io_A_Valid_1_delay_4_3;
    io_A_Valid_1_delay_6_1 <= io_A_Valid_1_delay_5_2;
    io_A_Valid_1_delay_7 <= io_A_Valid_1_delay_6_1;
    io_B_Valid_7_delay_1 <= io_B_Valid_7;
    io_B_Valid_0_delay_1_1 <= io_B_Valid_0;
    io_B_Valid_0_delay_2 <= io_B_Valid_0_delay_1_1;
    io_A_Valid_2_delay_1 <= io_A_Valid_2;
    io_B_Valid_1_delay_1_1 <= io_B_Valid_1;
    io_B_Valid_1_delay_2 <= io_B_Valid_1_delay_1_1;
    io_A_Valid_2_delay_1_1 <= io_A_Valid_2;
    io_A_Valid_2_delay_2 <= io_A_Valid_2_delay_1_1;
    io_B_Valid_2_delay_1_1 <= io_B_Valid_2;
    io_B_Valid_2_delay_2 <= io_B_Valid_2_delay_1_1;
    io_A_Valid_2_delay_1_2 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_1 <= io_A_Valid_2_delay_1_2;
    io_A_Valid_2_delay_3 <= io_A_Valid_2_delay_2_1;
    io_B_Valid_3_delay_1_1 <= io_B_Valid_3;
    io_B_Valid_3_delay_2 <= io_B_Valid_3_delay_1_1;
    io_A_Valid_2_delay_1_3 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_2 <= io_A_Valid_2_delay_1_3;
    io_A_Valid_2_delay_3_1 <= io_A_Valid_2_delay_2_2;
    io_A_Valid_2_delay_4 <= io_A_Valid_2_delay_3_1;
    io_B_Valid_4_delay_1_1 <= io_B_Valid_4;
    io_B_Valid_4_delay_2 <= io_B_Valid_4_delay_1_1;
    io_A_Valid_2_delay_1_4 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_3 <= io_A_Valid_2_delay_1_4;
    io_A_Valid_2_delay_3_2 <= io_A_Valid_2_delay_2_3;
    io_A_Valid_2_delay_4_1 <= io_A_Valid_2_delay_3_2;
    io_A_Valid_2_delay_5 <= io_A_Valid_2_delay_4_1;
    io_B_Valid_5_delay_1_1 <= io_B_Valid_5;
    io_B_Valid_5_delay_2 <= io_B_Valid_5_delay_1_1;
    io_A_Valid_2_delay_1_5 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_4 <= io_A_Valid_2_delay_1_5;
    io_A_Valid_2_delay_3_3 <= io_A_Valid_2_delay_2_4;
    io_A_Valid_2_delay_4_2 <= io_A_Valid_2_delay_3_3;
    io_A_Valid_2_delay_5_1 <= io_A_Valid_2_delay_4_2;
    io_A_Valid_2_delay_6 <= io_A_Valid_2_delay_5_1;
    io_B_Valid_6_delay_1_1 <= io_B_Valid_6;
    io_B_Valid_6_delay_2 <= io_B_Valid_6_delay_1_1;
    io_A_Valid_2_delay_1_6 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_5 <= io_A_Valid_2_delay_1_6;
    io_A_Valid_2_delay_3_4 <= io_A_Valid_2_delay_2_5;
    io_A_Valid_2_delay_4_3 <= io_A_Valid_2_delay_3_4;
    io_A_Valid_2_delay_5_2 <= io_A_Valid_2_delay_4_3;
    io_A_Valid_2_delay_6_1 <= io_A_Valid_2_delay_5_2;
    io_A_Valid_2_delay_7 <= io_A_Valid_2_delay_6_1;
    io_B_Valid_7_delay_1_1 <= io_B_Valid_7;
    io_B_Valid_7_delay_2 <= io_B_Valid_7_delay_1_1;
    io_B_Valid_0_delay_1_2 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_1 <= io_B_Valid_0_delay_1_2;
    io_B_Valid_0_delay_3 <= io_B_Valid_0_delay_2_1;
    io_A_Valid_3_delay_1 <= io_A_Valid_3;
    io_B_Valid_1_delay_1_2 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_1 <= io_B_Valid_1_delay_1_2;
    io_B_Valid_1_delay_3 <= io_B_Valid_1_delay_2_1;
    io_A_Valid_3_delay_1_1 <= io_A_Valid_3;
    io_A_Valid_3_delay_2 <= io_A_Valid_3_delay_1_1;
    io_B_Valid_2_delay_1_2 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_1 <= io_B_Valid_2_delay_1_2;
    io_B_Valid_2_delay_3 <= io_B_Valid_2_delay_2_1;
    io_A_Valid_3_delay_1_2 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_1 <= io_A_Valid_3_delay_1_2;
    io_A_Valid_3_delay_3 <= io_A_Valid_3_delay_2_1;
    io_B_Valid_3_delay_1_2 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_1 <= io_B_Valid_3_delay_1_2;
    io_B_Valid_3_delay_3 <= io_B_Valid_3_delay_2_1;
    io_A_Valid_3_delay_1_3 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_2 <= io_A_Valid_3_delay_1_3;
    io_A_Valid_3_delay_3_1 <= io_A_Valid_3_delay_2_2;
    io_A_Valid_3_delay_4 <= io_A_Valid_3_delay_3_1;
    io_B_Valid_4_delay_1_2 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_1 <= io_B_Valid_4_delay_1_2;
    io_B_Valid_4_delay_3 <= io_B_Valid_4_delay_2_1;
    io_A_Valid_3_delay_1_4 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_3 <= io_A_Valid_3_delay_1_4;
    io_A_Valid_3_delay_3_2 <= io_A_Valid_3_delay_2_3;
    io_A_Valid_3_delay_4_1 <= io_A_Valid_3_delay_3_2;
    io_A_Valid_3_delay_5 <= io_A_Valid_3_delay_4_1;
    io_B_Valid_5_delay_1_2 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_1 <= io_B_Valid_5_delay_1_2;
    io_B_Valid_5_delay_3 <= io_B_Valid_5_delay_2_1;
    io_A_Valid_3_delay_1_5 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_4 <= io_A_Valid_3_delay_1_5;
    io_A_Valid_3_delay_3_3 <= io_A_Valid_3_delay_2_4;
    io_A_Valid_3_delay_4_2 <= io_A_Valid_3_delay_3_3;
    io_A_Valid_3_delay_5_1 <= io_A_Valid_3_delay_4_2;
    io_A_Valid_3_delay_6 <= io_A_Valid_3_delay_5_1;
    io_B_Valid_6_delay_1_2 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_1 <= io_B_Valid_6_delay_1_2;
    io_B_Valid_6_delay_3 <= io_B_Valid_6_delay_2_1;
    io_A_Valid_3_delay_1_6 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_5 <= io_A_Valid_3_delay_1_6;
    io_A_Valid_3_delay_3_4 <= io_A_Valid_3_delay_2_5;
    io_A_Valid_3_delay_4_3 <= io_A_Valid_3_delay_3_4;
    io_A_Valid_3_delay_5_2 <= io_A_Valid_3_delay_4_3;
    io_A_Valid_3_delay_6_1 <= io_A_Valid_3_delay_5_2;
    io_A_Valid_3_delay_7 <= io_A_Valid_3_delay_6_1;
    io_B_Valid_7_delay_1_2 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_1 <= io_B_Valid_7_delay_1_2;
    io_B_Valid_7_delay_3 <= io_B_Valid_7_delay_2_1;
    io_B_Valid_0_delay_1_3 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_2 <= io_B_Valid_0_delay_1_3;
    io_B_Valid_0_delay_3_1 <= io_B_Valid_0_delay_2_2;
    io_B_Valid_0_delay_4 <= io_B_Valid_0_delay_3_1;
    io_A_Valid_4_delay_1 <= io_A_Valid_4;
    io_B_Valid_1_delay_1_3 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_2 <= io_B_Valid_1_delay_1_3;
    io_B_Valid_1_delay_3_1 <= io_B_Valid_1_delay_2_2;
    io_B_Valid_1_delay_4 <= io_B_Valid_1_delay_3_1;
    io_A_Valid_4_delay_1_1 <= io_A_Valid_4;
    io_A_Valid_4_delay_2 <= io_A_Valid_4_delay_1_1;
    io_B_Valid_2_delay_1_3 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_2 <= io_B_Valid_2_delay_1_3;
    io_B_Valid_2_delay_3_1 <= io_B_Valid_2_delay_2_2;
    io_B_Valid_2_delay_4 <= io_B_Valid_2_delay_3_1;
    io_A_Valid_4_delay_1_2 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_1 <= io_A_Valid_4_delay_1_2;
    io_A_Valid_4_delay_3 <= io_A_Valid_4_delay_2_1;
    io_B_Valid_3_delay_1_3 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_2 <= io_B_Valid_3_delay_1_3;
    io_B_Valid_3_delay_3_1 <= io_B_Valid_3_delay_2_2;
    io_B_Valid_3_delay_4 <= io_B_Valid_3_delay_3_1;
    io_A_Valid_4_delay_1_3 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_2 <= io_A_Valid_4_delay_1_3;
    io_A_Valid_4_delay_3_1 <= io_A_Valid_4_delay_2_2;
    io_A_Valid_4_delay_4 <= io_A_Valid_4_delay_3_1;
    io_B_Valid_4_delay_1_3 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_2 <= io_B_Valid_4_delay_1_3;
    io_B_Valid_4_delay_3_1 <= io_B_Valid_4_delay_2_2;
    io_B_Valid_4_delay_4 <= io_B_Valid_4_delay_3_1;
    io_A_Valid_4_delay_1_4 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_3 <= io_A_Valid_4_delay_1_4;
    io_A_Valid_4_delay_3_2 <= io_A_Valid_4_delay_2_3;
    io_A_Valid_4_delay_4_1 <= io_A_Valid_4_delay_3_2;
    io_A_Valid_4_delay_5 <= io_A_Valid_4_delay_4_1;
    io_B_Valid_5_delay_1_3 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_2 <= io_B_Valid_5_delay_1_3;
    io_B_Valid_5_delay_3_1 <= io_B_Valid_5_delay_2_2;
    io_B_Valid_5_delay_4 <= io_B_Valid_5_delay_3_1;
    io_A_Valid_4_delay_1_5 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_4 <= io_A_Valid_4_delay_1_5;
    io_A_Valid_4_delay_3_3 <= io_A_Valid_4_delay_2_4;
    io_A_Valid_4_delay_4_2 <= io_A_Valid_4_delay_3_3;
    io_A_Valid_4_delay_5_1 <= io_A_Valid_4_delay_4_2;
    io_A_Valid_4_delay_6 <= io_A_Valid_4_delay_5_1;
    io_B_Valid_6_delay_1_3 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_2 <= io_B_Valid_6_delay_1_3;
    io_B_Valid_6_delay_3_1 <= io_B_Valid_6_delay_2_2;
    io_B_Valid_6_delay_4 <= io_B_Valid_6_delay_3_1;
    io_A_Valid_4_delay_1_6 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_5 <= io_A_Valid_4_delay_1_6;
    io_A_Valid_4_delay_3_4 <= io_A_Valid_4_delay_2_5;
    io_A_Valid_4_delay_4_3 <= io_A_Valid_4_delay_3_4;
    io_A_Valid_4_delay_5_2 <= io_A_Valid_4_delay_4_3;
    io_A_Valid_4_delay_6_1 <= io_A_Valid_4_delay_5_2;
    io_A_Valid_4_delay_7 <= io_A_Valid_4_delay_6_1;
    io_B_Valid_7_delay_1_3 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_2 <= io_B_Valid_7_delay_1_3;
    io_B_Valid_7_delay_3_1 <= io_B_Valid_7_delay_2_2;
    io_B_Valid_7_delay_4 <= io_B_Valid_7_delay_3_1;
    io_B_Valid_0_delay_1_4 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_3 <= io_B_Valid_0_delay_1_4;
    io_B_Valid_0_delay_3_2 <= io_B_Valid_0_delay_2_3;
    io_B_Valid_0_delay_4_1 <= io_B_Valid_0_delay_3_2;
    io_B_Valid_0_delay_5 <= io_B_Valid_0_delay_4_1;
    io_A_Valid_5_delay_1 <= io_A_Valid_5;
    io_B_Valid_1_delay_1_4 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_3 <= io_B_Valid_1_delay_1_4;
    io_B_Valid_1_delay_3_2 <= io_B_Valid_1_delay_2_3;
    io_B_Valid_1_delay_4_1 <= io_B_Valid_1_delay_3_2;
    io_B_Valid_1_delay_5 <= io_B_Valid_1_delay_4_1;
    io_A_Valid_5_delay_1_1 <= io_A_Valid_5;
    io_A_Valid_5_delay_2 <= io_A_Valid_5_delay_1_1;
    io_B_Valid_2_delay_1_4 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_3 <= io_B_Valid_2_delay_1_4;
    io_B_Valid_2_delay_3_2 <= io_B_Valid_2_delay_2_3;
    io_B_Valid_2_delay_4_1 <= io_B_Valid_2_delay_3_2;
    io_B_Valid_2_delay_5 <= io_B_Valid_2_delay_4_1;
    io_A_Valid_5_delay_1_2 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_1 <= io_A_Valid_5_delay_1_2;
    io_A_Valid_5_delay_3 <= io_A_Valid_5_delay_2_1;
    io_B_Valid_3_delay_1_4 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_3 <= io_B_Valid_3_delay_1_4;
    io_B_Valid_3_delay_3_2 <= io_B_Valid_3_delay_2_3;
    io_B_Valid_3_delay_4_1 <= io_B_Valid_3_delay_3_2;
    io_B_Valid_3_delay_5 <= io_B_Valid_3_delay_4_1;
    io_A_Valid_5_delay_1_3 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_2 <= io_A_Valid_5_delay_1_3;
    io_A_Valid_5_delay_3_1 <= io_A_Valid_5_delay_2_2;
    io_A_Valid_5_delay_4 <= io_A_Valid_5_delay_3_1;
    io_B_Valid_4_delay_1_4 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_3 <= io_B_Valid_4_delay_1_4;
    io_B_Valid_4_delay_3_2 <= io_B_Valid_4_delay_2_3;
    io_B_Valid_4_delay_4_1 <= io_B_Valid_4_delay_3_2;
    io_B_Valid_4_delay_5 <= io_B_Valid_4_delay_4_1;
    io_A_Valid_5_delay_1_4 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_3 <= io_A_Valid_5_delay_1_4;
    io_A_Valid_5_delay_3_2 <= io_A_Valid_5_delay_2_3;
    io_A_Valid_5_delay_4_1 <= io_A_Valid_5_delay_3_2;
    io_A_Valid_5_delay_5 <= io_A_Valid_5_delay_4_1;
    io_B_Valid_5_delay_1_4 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_3 <= io_B_Valid_5_delay_1_4;
    io_B_Valid_5_delay_3_2 <= io_B_Valid_5_delay_2_3;
    io_B_Valid_5_delay_4_1 <= io_B_Valid_5_delay_3_2;
    io_B_Valid_5_delay_5 <= io_B_Valid_5_delay_4_1;
    io_A_Valid_5_delay_1_5 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_4 <= io_A_Valid_5_delay_1_5;
    io_A_Valid_5_delay_3_3 <= io_A_Valid_5_delay_2_4;
    io_A_Valid_5_delay_4_2 <= io_A_Valid_5_delay_3_3;
    io_A_Valid_5_delay_5_1 <= io_A_Valid_5_delay_4_2;
    io_A_Valid_5_delay_6 <= io_A_Valid_5_delay_5_1;
    io_B_Valid_6_delay_1_4 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_3 <= io_B_Valid_6_delay_1_4;
    io_B_Valid_6_delay_3_2 <= io_B_Valid_6_delay_2_3;
    io_B_Valid_6_delay_4_1 <= io_B_Valid_6_delay_3_2;
    io_B_Valid_6_delay_5 <= io_B_Valid_6_delay_4_1;
    io_A_Valid_5_delay_1_6 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_5 <= io_A_Valid_5_delay_1_6;
    io_A_Valid_5_delay_3_4 <= io_A_Valid_5_delay_2_5;
    io_A_Valid_5_delay_4_3 <= io_A_Valid_5_delay_3_4;
    io_A_Valid_5_delay_5_2 <= io_A_Valid_5_delay_4_3;
    io_A_Valid_5_delay_6_1 <= io_A_Valid_5_delay_5_2;
    io_A_Valid_5_delay_7 <= io_A_Valid_5_delay_6_1;
    io_B_Valid_7_delay_1_4 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_3 <= io_B_Valid_7_delay_1_4;
    io_B_Valid_7_delay_3_2 <= io_B_Valid_7_delay_2_3;
    io_B_Valid_7_delay_4_1 <= io_B_Valid_7_delay_3_2;
    io_B_Valid_7_delay_5 <= io_B_Valid_7_delay_4_1;
    io_B_Valid_0_delay_1_5 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_4 <= io_B_Valid_0_delay_1_5;
    io_B_Valid_0_delay_3_3 <= io_B_Valid_0_delay_2_4;
    io_B_Valid_0_delay_4_2 <= io_B_Valid_0_delay_3_3;
    io_B_Valid_0_delay_5_1 <= io_B_Valid_0_delay_4_2;
    io_B_Valid_0_delay_6 <= io_B_Valid_0_delay_5_1;
    io_A_Valid_6_delay_1 <= io_A_Valid_6;
    io_B_Valid_1_delay_1_5 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_4 <= io_B_Valid_1_delay_1_5;
    io_B_Valid_1_delay_3_3 <= io_B_Valid_1_delay_2_4;
    io_B_Valid_1_delay_4_2 <= io_B_Valid_1_delay_3_3;
    io_B_Valid_1_delay_5_1 <= io_B_Valid_1_delay_4_2;
    io_B_Valid_1_delay_6 <= io_B_Valid_1_delay_5_1;
    io_A_Valid_6_delay_1_1 <= io_A_Valid_6;
    io_A_Valid_6_delay_2 <= io_A_Valid_6_delay_1_1;
    io_B_Valid_2_delay_1_5 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_4 <= io_B_Valid_2_delay_1_5;
    io_B_Valid_2_delay_3_3 <= io_B_Valid_2_delay_2_4;
    io_B_Valid_2_delay_4_2 <= io_B_Valid_2_delay_3_3;
    io_B_Valid_2_delay_5_1 <= io_B_Valid_2_delay_4_2;
    io_B_Valid_2_delay_6 <= io_B_Valid_2_delay_5_1;
    io_A_Valid_6_delay_1_2 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_1 <= io_A_Valid_6_delay_1_2;
    io_A_Valid_6_delay_3 <= io_A_Valid_6_delay_2_1;
    io_B_Valid_3_delay_1_5 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_4 <= io_B_Valid_3_delay_1_5;
    io_B_Valid_3_delay_3_3 <= io_B_Valid_3_delay_2_4;
    io_B_Valid_3_delay_4_2 <= io_B_Valid_3_delay_3_3;
    io_B_Valid_3_delay_5_1 <= io_B_Valid_3_delay_4_2;
    io_B_Valid_3_delay_6 <= io_B_Valid_3_delay_5_1;
    io_A_Valid_6_delay_1_3 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_2 <= io_A_Valid_6_delay_1_3;
    io_A_Valid_6_delay_3_1 <= io_A_Valid_6_delay_2_2;
    io_A_Valid_6_delay_4 <= io_A_Valid_6_delay_3_1;
    io_B_Valid_4_delay_1_5 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_4 <= io_B_Valid_4_delay_1_5;
    io_B_Valid_4_delay_3_3 <= io_B_Valid_4_delay_2_4;
    io_B_Valid_4_delay_4_2 <= io_B_Valid_4_delay_3_3;
    io_B_Valid_4_delay_5_1 <= io_B_Valid_4_delay_4_2;
    io_B_Valid_4_delay_6 <= io_B_Valid_4_delay_5_1;
    io_A_Valid_6_delay_1_4 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_3 <= io_A_Valid_6_delay_1_4;
    io_A_Valid_6_delay_3_2 <= io_A_Valid_6_delay_2_3;
    io_A_Valid_6_delay_4_1 <= io_A_Valid_6_delay_3_2;
    io_A_Valid_6_delay_5 <= io_A_Valid_6_delay_4_1;
    io_B_Valid_5_delay_1_5 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_4 <= io_B_Valid_5_delay_1_5;
    io_B_Valid_5_delay_3_3 <= io_B_Valid_5_delay_2_4;
    io_B_Valid_5_delay_4_2 <= io_B_Valid_5_delay_3_3;
    io_B_Valid_5_delay_5_1 <= io_B_Valid_5_delay_4_2;
    io_B_Valid_5_delay_6 <= io_B_Valid_5_delay_5_1;
    io_A_Valid_6_delay_1_5 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_4 <= io_A_Valid_6_delay_1_5;
    io_A_Valid_6_delay_3_3 <= io_A_Valid_6_delay_2_4;
    io_A_Valid_6_delay_4_2 <= io_A_Valid_6_delay_3_3;
    io_A_Valid_6_delay_5_1 <= io_A_Valid_6_delay_4_2;
    io_A_Valid_6_delay_6 <= io_A_Valid_6_delay_5_1;
    io_B_Valid_6_delay_1_5 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_4 <= io_B_Valid_6_delay_1_5;
    io_B_Valid_6_delay_3_3 <= io_B_Valid_6_delay_2_4;
    io_B_Valid_6_delay_4_2 <= io_B_Valid_6_delay_3_3;
    io_B_Valid_6_delay_5_1 <= io_B_Valid_6_delay_4_2;
    io_B_Valid_6_delay_6 <= io_B_Valid_6_delay_5_1;
    io_A_Valid_6_delay_1_6 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_5 <= io_A_Valid_6_delay_1_6;
    io_A_Valid_6_delay_3_4 <= io_A_Valid_6_delay_2_5;
    io_A_Valid_6_delay_4_3 <= io_A_Valid_6_delay_3_4;
    io_A_Valid_6_delay_5_2 <= io_A_Valid_6_delay_4_3;
    io_A_Valid_6_delay_6_1 <= io_A_Valid_6_delay_5_2;
    io_A_Valid_6_delay_7 <= io_A_Valid_6_delay_6_1;
    io_B_Valid_7_delay_1_5 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_4 <= io_B_Valid_7_delay_1_5;
    io_B_Valid_7_delay_3_3 <= io_B_Valid_7_delay_2_4;
    io_B_Valid_7_delay_4_2 <= io_B_Valid_7_delay_3_3;
    io_B_Valid_7_delay_5_1 <= io_B_Valid_7_delay_4_2;
    io_B_Valid_7_delay_6 <= io_B_Valid_7_delay_5_1;
    io_B_Valid_0_delay_1_6 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_5 <= io_B_Valid_0_delay_1_6;
    io_B_Valid_0_delay_3_4 <= io_B_Valid_0_delay_2_5;
    io_B_Valid_0_delay_4_3 <= io_B_Valid_0_delay_3_4;
    io_B_Valid_0_delay_5_2 <= io_B_Valid_0_delay_4_3;
    io_B_Valid_0_delay_6_1 <= io_B_Valid_0_delay_5_2;
    io_B_Valid_0_delay_7 <= io_B_Valid_0_delay_6_1;
    io_A_Valid_7_delay_1 <= io_A_Valid_7;
    io_B_Valid_1_delay_1_6 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_5 <= io_B_Valid_1_delay_1_6;
    io_B_Valid_1_delay_3_4 <= io_B_Valid_1_delay_2_5;
    io_B_Valid_1_delay_4_3 <= io_B_Valid_1_delay_3_4;
    io_B_Valid_1_delay_5_2 <= io_B_Valid_1_delay_4_3;
    io_B_Valid_1_delay_6_1 <= io_B_Valid_1_delay_5_2;
    io_B_Valid_1_delay_7 <= io_B_Valid_1_delay_6_1;
    io_A_Valid_7_delay_1_1 <= io_A_Valid_7;
    io_A_Valid_7_delay_2 <= io_A_Valid_7_delay_1_1;
    io_B_Valid_2_delay_1_6 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_5 <= io_B_Valid_2_delay_1_6;
    io_B_Valid_2_delay_3_4 <= io_B_Valid_2_delay_2_5;
    io_B_Valid_2_delay_4_3 <= io_B_Valid_2_delay_3_4;
    io_B_Valid_2_delay_5_2 <= io_B_Valid_2_delay_4_3;
    io_B_Valid_2_delay_6_1 <= io_B_Valid_2_delay_5_2;
    io_B_Valid_2_delay_7 <= io_B_Valid_2_delay_6_1;
    io_A_Valid_7_delay_1_2 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_1 <= io_A_Valid_7_delay_1_2;
    io_A_Valid_7_delay_3 <= io_A_Valid_7_delay_2_1;
    io_B_Valid_3_delay_1_6 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_5 <= io_B_Valid_3_delay_1_6;
    io_B_Valid_3_delay_3_4 <= io_B_Valid_3_delay_2_5;
    io_B_Valid_3_delay_4_3 <= io_B_Valid_3_delay_3_4;
    io_B_Valid_3_delay_5_2 <= io_B_Valid_3_delay_4_3;
    io_B_Valid_3_delay_6_1 <= io_B_Valid_3_delay_5_2;
    io_B_Valid_3_delay_7 <= io_B_Valid_3_delay_6_1;
    io_A_Valid_7_delay_1_3 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_2 <= io_A_Valid_7_delay_1_3;
    io_A_Valid_7_delay_3_1 <= io_A_Valid_7_delay_2_2;
    io_A_Valid_7_delay_4 <= io_A_Valid_7_delay_3_1;
    io_B_Valid_4_delay_1_6 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_5 <= io_B_Valid_4_delay_1_6;
    io_B_Valid_4_delay_3_4 <= io_B_Valid_4_delay_2_5;
    io_B_Valid_4_delay_4_3 <= io_B_Valid_4_delay_3_4;
    io_B_Valid_4_delay_5_2 <= io_B_Valid_4_delay_4_3;
    io_B_Valid_4_delay_6_1 <= io_B_Valid_4_delay_5_2;
    io_B_Valid_4_delay_7 <= io_B_Valid_4_delay_6_1;
    io_A_Valid_7_delay_1_4 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_3 <= io_A_Valid_7_delay_1_4;
    io_A_Valid_7_delay_3_2 <= io_A_Valid_7_delay_2_3;
    io_A_Valid_7_delay_4_1 <= io_A_Valid_7_delay_3_2;
    io_A_Valid_7_delay_5 <= io_A_Valid_7_delay_4_1;
    io_B_Valid_5_delay_1_6 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_5 <= io_B_Valid_5_delay_1_6;
    io_B_Valid_5_delay_3_4 <= io_B_Valid_5_delay_2_5;
    io_B_Valid_5_delay_4_3 <= io_B_Valid_5_delay_3_4;
    io_B_Valid_5_delay_5_2 <= io_B_Valid_5_delay_4_3;
    io_B_Valid_5_delay_6_1 <= io_B_Valid_5_delay_5_2;
    io_B_Valid_5_delay_7 <= io_B_Valid_5_delay_6_1;
    io_A_Valid_7_delay_1_5 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_4 <= io_A_Valid_7_delay_1_5;
    io_A_Valid_7_delay_3_3 <= io_A_Valid_7_delay_2_4;
    io_A_Valid_7_delay_4_2 <= io_A_Valid_7_delay_3_3;
    io_A_Valid_7_delay_5_1 <= io_A_Valid_7_delay_4_2;
    io_A_Valid_7_delay_6 <= io_A_Valid_7_delay_5_1;
    io_B_Valid_6_delay_1_6 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_5 <= io_B_Valid_6_delay_1_6;
    io_B_Valid_6_delay_3_4 <= io_B_Valid_6_delay_2_5;
    io_B_Valid_6_delay_4_3 <= io_B_Valid_6_delay_3_4;
    io_B_Valid_6_delay_5_2 <= io_B_Valid_6_delay_4_3;
    io_B_Valid_6_delay_6_1 <= io_B_Valid_6_delay_5_2;
    io_B_Valid_6_delay_7 <= io_B_Valid_6_delay_6_1;
    io_A_Valid_7_delay_1_6 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_5 <= io_A_Valid_7_delay_1_6;
    io_A_Valid_7_delay_3_4 <= io_A_Valid_7_delay_2_5;
    io_A_Valid_7_delay_4_3 <= io_A_Valid_7_delay_3_4;
    io_A_Valid_7_delay_5_2 <= io_A_Valid_7_delay_4_3;
    io_A_Valid_7_delay_6_1 <= io_A_Valid_7_delay_5_2;
    io_A_Valid_7_delay_7 <= io_A_Valid_7_delay_6_1;
    io_B_Valid_7_delay_1_6 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_5 <= io_B_Valid_7_delay_1_6;
    io_B_Valid_7_delay_3_4 <= io_B_Valid_7_delay_2_5;
    io_B_Valid_7_delay_4_3 <= io_B_Valid_7_delay_3_4;
    io_B_Valid_7_delay_5_2 <= io_B_Valid_7_delay_4_3;
    io_B_Valid_7_delay_6_1 <= io_B_Valid_7_delay_5_2;
    io_B_Valid_7_delay_7 <= io_B_Valid_7_delay_6_1;
  end


endmodule

//AxisDataConverter_7 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

//AxisDataConverter_6 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

//AxisDataConverter_5 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

//AxisDataConverter_4 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

//AxisDataConverter_3 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

//AxisDataConverter_2 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

//AxisDataConverter_1 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

module AxisDataConverter (
  input               inStream_valid,
  output              inStream_ready,
  input      [63:0]   inStream_payload,
  output              outStream_valid,
  input               outStream_ready,
  output     [7:0]    outStream_payload,
  input               clk,
  input               reset
);

  wire       [2:0]    _zz__zz_outStream_payload_1;
  wire       [0:0]    _zz__zz_outStream_payload_1_1;
  wire       [63:0]   _zz__zz_outStream_payload_3;
  reg        [7:0]    _zz_outStream_payload_4;
  wire                outStream_fire;
  reg                 _zz_outStream_payload;
  reg        [2:0]    _zz_outStream_payload_1;
  reg        [2:0]    _zz_outStream_payload_2;
  wire                _zz_inStream_ready;
  wire       [63:0]   _zz_outStream_payload_3;

  assign _zz__zz_outStream_payload_1_1 = _zz_outStream_payload;
  assign _zz__zz_outStream_payload_1 = {2'd0, _zz__zz_outStream_payload_1_1};
  assign _zz__zz_outStream_payload_3 = inStream_payload;
  always @(*) begin
    case(_zz_outStream_payload_2)
      3'b000 : _zz_outStream_payload_4 = _zz_outStream_payload_3[7 : 0];
      3'b001 : _zz_outStream_payload_4 = _zz_outStream_payload_3[15 : 8];
      3'b010 : _zz_outStream_payload_4 = _zz_outStream_payload_3[23 : 16];
      3'b011 : _zz_outStream_payload_4 = _zz_outStream_payload_3[31 : 24];
      3'b100 : _zz_outStream_payload_4 = _zz_outStream_payload_3[39 : 32];
      3'b101 : _zz_outStream_payload_4 = _zz_outStream_payload_3[47 : 40];
      3'b110 : _zz_outStream_payload_4 = _zz_outStream_payload_3[55 : 48];
      default : _zz_outStream_payload_4 = _zz_outStream_payload_3[63 : 56];
    endcase
  end

  assign outStream_fire = (outStream_valid && outStream_ready);
  always @(*) begin
    _zz_outStream_payload = 1'b0;
    if(outStream_fire) begin
      _zz_outStream_payload = 1'b1;
    end
  end

  assign _zz_inStream_ready = (_zz_outStream_payload_2 == 3'b111);
  always @(*) begin
    _zz_outStream_payload_1 = (_zz_outStream_payload_2 + _zz__zz_outStream_payload_1);
    if(1'b0) begin
      _zz_outStream_payload_1 = 3'b000;
    end
  end

  assign outStream_valid = inStream_valid;
  assign _zz_outStream_payload_3 = _zz__zz_outStream_payload_3;
  assign outStream_payload = _zz_outStream_payload_4;
  assign inStream_ready = (outStream_ready && _zz_inStream_ready);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _zz_outStream_payload_2 <= 3'b000;
    end else begin
      _zz_outStream_payload_2 <= _zz_outStream_payload_1;
    end
  end


endmodule

module Img2Col_WidthConverter_Fifo (
  input               io_push_valid,
  output              io_push_ready,
  input      [63:0]   io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [63:0]   io_pop_payload,
  input               io_flush,
  output     [4:0]    io_occupancy,
  output     [4:0]    io_availability,
  input               clk,
  input               reset
);

  reg        [63:0]   _zz_logic_ram_port0;
  wire       [3:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [3:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [63:0]   _zz_logic_ram_port_1;
  wire       [3:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [3:0]    logic_pushPtr_valueNext;
  reg        [3:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [3:0]    logic_popPtr_valueNext;
  reg        [3:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1122;
  wire       [3:0]    logic_ptrDif;
  reg [63:0] logic_ram [0:15];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {3'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {3'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  assign _zz_logic_ram_port_1 = io_push_payload;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 4'b1111);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 4'b0000;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 4'b1111);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 4'b0000;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1122 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_pushPtr_value <= 4'b0000;
      logic_popPtr_value <= 4'b0000;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1122) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module Img2Col_Top (
  input               start,
  input               sData_valid,
  output              sData_ready,
  input      [63:0]   sData_payload,
  output     [63:0]   mData,
  input               mReady,
  output              mValid,
  input               Fifo_Clear,
  output              mLast,
  input      [4:0]    Stride,
  input      [4:0]    Kernel_Size,
  input      [15:0]   Window_Size,
  input      [15:0]   InFeature_Size,
  input      [15:0]   InFeature_Channel,
  input      [15:0]   OutFeature_Channel,
  input      [15:0]   OutFeature_Size,
  input      [15:0]   OutCol_Count_Times,
  input      [15:0]   InCol_Count_Times,
  input      [15:0]   OutRow_Count_Times,
  input      [15:0]   OutFeature_Channel_Count_Times,
  input      [12:0]   Sliding_Size,
  output              Test_Signal,
  input      [15:0]   Test_Generate_Period,
  output              Test_End,
  output              Raddr_Valid,
  output              LayerEnd,
  output              SA_Row_Cnt_Valid,
  input               clk,
  input               reset
);
  localparam IMG2COL_ENUM_IDLE = 7'd1;
  localparam IMG2COL_ENUM_INIT = 7'd2;
  localparam IMG2COL_ENUM_INIT_ADDR = 7'd4;
  localparam IMG2COL_ENUM_DATA_CACHE = 7'd8;
  localparam IMG2COL_ENUM_WAIT_COMPUTE = 7'd16;
  localparam IMG2COL_ENUM_UPDATE_ADDR = 7'd32;
  localparam IMG2COL_ENUM_START_COMPUTE = 7'd64;

  reg                 AddrFifo_io_push_valid;
  reg                 AddrFifo_io_pop_ready;
  wire                AddrFifo_io_flush;
  reg                 RaddrFifo0_io_push_valid;
  reg        [15:0]   RaddrFifo0_io_push_payload;
  reg                 RaddrFifo0_io_pop_ready;
  wire                RaddrFifo0_io_flush;
  wire                Img2Col_SubModule_start;
  wire                Img2Col_SubModule_NewAddrIn_valid;
  wire       [13:0]   DGB_addra;
  wire       [13:0]   DGB_addrb;
  wire                AddrFifo_io_push_ready;
  wire                AddrFifo_io_pop_valid;
  wire       [15:0]   AddrFifo_io_pop_payload;
  wire       [5:0]    AddrFifo_io_occupancy;
  wire       [5:0]    AddrFifo_io_availability;
  wire                RaddrFifo0_io_push_ready;
  wire                RaddrFifo0_io_pop_valid;
  wire       [15:0]   RaddrFifo0_io_pop_payload;
  wire       [5:0]    RaddrFifo0_io_occupancy;
  wire       [5:0]    RaddrFifo0_io_availability;
  wire                Img2Col_SubModule_NewAddrIn_ready;
  wire                Img2Col_SubModule_SA_Idle;
  wire       [15:0]   Img2Col_SubModule_Raddr;
  wire                Img2Col_SubModule_Raddr_Valid;
  wire                Img2Col_SubModule_SA_End;
  wire                Img2Col_SubModule_AddrReceived;
  wire                Img2Col_SubModule_SA_Row_Cnt_Valid;
  wire       [63:0]   DGB_doutb;
  wire       [4:0]    _zz_Addr_Init_Cnt_valid;
  wire       [4:0]    _zz_Addr_Init_Cnt_valid_1;
  wire       [15:0]   _zz_In_Col_Cnt_valid;
  wire       [4:0]    _zz_Row_Cache_Cnt_valid;
  wire       [15:0]   _zz_In_Row_Cnt_valid;
  wire       [15:0]   _zz_when_Data_Generate_V2_l217;
  wire       [4:0]    _zz_when_Data_Generate_V2_l217_1;
  wire       [15:0]   _zz_Out_Row_Cnt_valid;
  wire       [15:0]   _zz_Test_Valid;
  reg                 start_regNext;
  wire                when_Data_Generate_V2_l59;
  reg        [6:0]    Fsm_currentState;
  reg        [6:0]    Fsm_nextState;
  wire                Fsm_Init_End;
  wire                Fsm_Addr_Inited;
  wire                Fsm_Data_Cached;
  wire                Fsm_Addr_Updated;
  wire                Fsm_SA_Ready;
  wire                Fsm_Cache_End;
  wire                Fsm_Layer_End;
  wire                when_WaCounter_l19;
  reg        [2:0]    Init_Count_count;
  reg                 Init_Count_valid;
  wire                when_WaCounter_l14;
  wire                when_WaCounter_l40;
  reg        [4:0]    Addr_Init_Cnt_count;
  wire                Addr_Init_Cnt_valid;
  reg        [15:0]   WaddrOffset;
  wire                when_Data_Generate_V2_l170;
  wire                when_Data_Generate_V2_l175;
  wire                SubModule_AddrFifo_io_pop_fire;
  wire                when_Data_Generate_V2_l179;
  wire                when_Data_Generate_V2_l183;
  reg        [15:0]   Raddr_Initialization;
  wire                when_Data_Generate_V2_l193;
  wire                when_Data_Generate_V2_l197;
  reg        [4:0]    Cache_Row_Num;
  reg        [4:0]    Raddr_Updata_Cnt_Num;
  wire                sData_fire;
  reg        [15:0]   In_Col_Cnt_count;
  wire                In_Col_Cnt_valid;
  reg        [4:0]    Row_Cache_Cnt_count;
  wire                Row_Cache_Cnt_valid;
  reg        [15:0]   In_Row_Cnt_count;
  wire                In_Row_Cnt_valid;
  wire                when_Data_Generate_V2_l217;
  reg                 CacheEnd_Flag;
  wire                when_Data_Generate_V2_l228;
  wire                Img2ColOutput_Module_Ready_Receive_Addr;
  wire                when_Data_Generate_V2_l245;
  wire                SubModule_RaddrFifo0_io_pop_fire;
  reg        [15:0]   Out_Row_Cnt_count;
  wire                Out_Row_Cnt_valid;
  wire       [15:0]   Waddr;
  wire                sData_fire_1;
  reg                 SubModule_Img2Col_SubModule_Raddr_Valid_regNext;
  reg                 Out_Row_Cnt_valid_regNext;
  reg        [15:0]   Out_Row_Cnt_count_regNext;
  wire                Test_Valid;
  reg                 Test_Valid_regNext;
  `ifndef SYNTHESIS
  reg [103:0] Fsm_currentState_string;
  reg [103:0] Fsm_nextState_string;
  `endif


  assign _zz_Addr_Init_Cnt_valid = (_zz_Addr_Init_Cnt_valid_1 - 5'h01);
  assign _zz_Addr_Init_Cnt_valid_1 = (Kernel_Size + Stride);
  assign _zz_In_Col_Cnt_valid = (InCol_Count_Times - 16'h0001);
  assign _zz_Row_Cache_Cnt_valid = (Cache_Row_Num - 5'h01);
  assign _zz_In_Row_Cnt_valid = (InFeature_Size - 16'h0001);
  assign _zz_when_Data_Generate_V2_l217_1 = (Kernel_Size - 5'h01);
  assign _zz_when_Data_Generate_V2_l217 = {11'd0, _zz_when_Data_Generate_V2_l217_1};
  assign _zz_Out_Row_Cnt_valid = (OutRow_Count_Times - 16'h0001);
  assign _zz_Test_Valid = (Test_Generate_Period - 16'h0001);
  WaddrOffset_Fifo_2 AddrFifo (
    .io_push_valid   (AddrFifo_io_push_valid       ), //i
    .io_push_ready   (AddrFifo_io_push_ready       ), //o
    .io_push_payload (WaddrOffset[15:0]            ), //i
    .io_pop_valid    (AddrFifo_io_pop_valid        ), //o
    .io_pop_ready    (AddrFifo_io_pop_ready        ), //i
    .io_pop_payload  (AddrFifo_io_pop_payload[15:0]), //o
    .io_flush        (AddrFifo_io_flush            ), //i
    .io_occupancy    (AddrFifo_io_occupancy[5:0]   ), //o
    .io_availability (AddrFifo_io_availability[5:0]), //o
    .clk             (clk                          ), //i
    .reset           (reset                        )  //i
  );
  WaddrOffset_Fifo_2 RaddrFifo0 (
    .io_push_valid   (RaddrFifo0_io_push_valid        ), //i
    .io_push_ready   (RaddrFifo0_io_push_ready        ), //o
    .io_push_payload (RaddrFifo0_io_push_payload[15:0]), //i
    .io_pop_valid    (RaddrFifo0_io_pop_valid         ), //o
    .io_pop_ready    (RaddrFifo0_io_pop_ready         ), //i
    .io_pop_payload  (RaddrFifo0_io_pop_payload[15:0] ), //o
    .io_flush        (RaddrFifo0_io_flush             ), //i
    .io_occupancy    (RaddrFifo0_io_occupancy[5:0]    ), //o
    .io_availability (RaddrFifo0_io_availability[5:0] ), //o
    .clk             (clk                             ), //i
    .reset           (reset                           )  //i
  );
  Img2Col_OutPut Img2Col_SubModule (
    .start                          (Img2Col_SubModule_start             ), //i
    .NewAddrIn_valid                (Img2Col_SubModule_NewAddrIn_valid   ), //i
    .NewAddrIn_ready                (Img2Col_SubModule_NewAddrIn_ready   ), //o
    .NewAddrIn_payload              (RaddrFifo0_io_pop_payload[15:0]     ), //i
    .SA_Idle                        (Img2Col_SubModule_SA_Idle           ), //o
    .Raddr                          (Img2Col_SubModule_Raddr[15:0]       ), //o
    .Raddr_Valid                    (Img2Col_SubModule_Raddr_Valid       ), //o
    .SA_End                         (Img2Col_SubModule_SA_End            ), //o
    .Stride                         (Stride[4:0]                         ), //i
    .Kernel_Size                    (Kernel_Size[4:0]                    ), //i
    .Window_Size                    (Window_Size[15:0]                   ), //i
    .InFeature_Size                 (InFeature_Size[15:0]                ), //i
    .InFeature_Channel              (InFeature_Channel[15:0]             ), //i
    .OutFeature_Channel             (OutFeature_Channel[15:0]            ), //i
    .OutFeature_Size                (OutFeature_Size[15:0]               ), //i
    .OutCol_Count_Times             (OutCol_Count_Times[15:0]            ), //i
    .InCol_Count_Times              (InCol_Count_Times[15:0]             ), //i
    .OutFeature_Channel_Count_Times (OutFeature_Channel_Count_Times[15:0]), //i
    .Sliding_Size                   (Sliding_Size[12:0]                  ), //i
    .mReady                         (mReady                              ), //i
    .Fifo_Clear                     (Fifo_Clear                          ), //i
    .AddrReceived                   (Img2Col_SubModule_AddrReceived      ), //o
    .LayerEnd                       (Fsm_Layer_End                       ), //i
    .SA_Row_Cnt_Valid               (Img2Col_SubModule_SA_Row_Cnt_Valid  ), //o
    .clk                            (clk                                 ), //i
    .reset                          (reset                               )  //i
  );
  DataGen_Bram DGB (
    .clka  (clk                ), //i
    .addra (DGB_addra[13:0]    ), //i
    .dina  (sData_payload[63:0]), //i
    .ena   (sData_fire_1       ), //i
    .wea   (1'b1               ), //i
    .addrb (DGB_addrb[13:0]    ), //i
    .doutb (DGB_doutb[63:0]    ), //o
    .clkb  (clk                )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      IMG2COL_ENUM_IDLE : Fsm_currentState_string = "IDLE         ";
      IMG2COL_ENUM_INIT : Fsm_currentState_string = "INIT         ";
      IMG2COL_ENUM_INIT_ADDR : Fsm_currentState_string = "INIT_ADDR    ";
      IMG2COL_ENUM_DATA_CACHE : Fsm_currentState_string = "DATA_CACHE   ";
      IMG2COL_ENUM_WAIT_COMPUTE : Fsm_currentState_string = "WAIT_COMPUTE ";
      IMG2COL_ENUM_UPDATE_ADDR : Fsm_currentState_string = "UPDATE_ADDR  ";
      IMG2COL_ENUM_START_COMPUTE : Fsm_currentState_string = "START_COMPUTE";
      default : Fsm_currentState_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      IMG2COL_ENUM_IDLE : Fsm_nextState_string = "IDLE         ";
      IMG2COL_ENUM_INIT : Fsm_nextState_string = "INIT         ";
      IMG2COL_ENUM_INIT_ADDR : Fsm_nextState_string = "INIT_ADDR    ";
      IMG2COL_ENUM_DATA_CACHE : Fsm_nextState_string = "DATA_CACHE   ";
      IMG2COL_ENUM_WAIT_COMPUTE : Fsm_nextState_string = "WAIT_COMPUTE ";
      IMG2COL_ENUM_UPDATE_ADDR : Fsm_nextState_string = "UPDATE_ADDR  ";
      IMG2COL_ENUM_START_COMPUTE : Fsm_nextState_string = "START_COMPUTE";
      default : Fsm_nextState_string = "?????????????";
    endcase
  end
  `endif

  assign when_Data_Generate_V2_l59 = (start && (! start_regNext));
  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & IMG2COL_ENUM_IDLE) == IMG2COL_ENUM_IDLE) : begin
        if(when_Data_Generate_V2_l59) begin
          Fsm_nextState = IMG2COL_ENUM_INIT;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_IDLE;
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_INIT) == IMG2COL_ENUM_INIT) : begin
        if(Fsm_Init_End) begin
          Fsm_nextState = IMG2COL_ENUM_INIT_ADDR;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_INIT;
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_INIT_ADDR) == IMG2COL_ENUM_INIT_ADDR) : begin
        if(Fsm_Addr_Inited) begin
          Fsm_nextState = IMG2COL_ENUM_DATA_CACHE;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_INIT_ADDR;
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_DATA_CACHE) == IMG2COL_ENUM_DATA_CACHE) : begin
        if(Fsm_Data_Cached) begin
          Fsm_nextState = IMG2COL_ENUM_WAIT_COMPUTE;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_DATA_CACHE;
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_WAIT_COMPUTE) == IMG2COL_ENUM_WAIT_COMPUTE) : begin
        if(Fsm_Layer_End) begin
          Fsm_nextState = IMG2COL_ENUM_IDLE;
        end else begin
          if(Fsm_SA_Ready) begin
            Fsm_nextState = IMG2COL_ENUM_UPDATE_ADDR;
          end else begin
            Fsm_nextState = IMG2COL_ENUM_WAIT_COMPUTE;
          end
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_UPDATE_ADDR) == IMG2COL_ENUM_UPDATE_ADDR) : begin
        if(Fsm_Addr_Updated) begin
          Fsm_nextState = IMG2COL_ENUM_START_COMPUTE;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_UPDATE_ADDR;
        end
      end
      default : begin
        if(Fsm_Layer_End) begin
          Fsm_nextState = IMG2COL_ENUM_IDLE;
        end else begin
          if(Fsm_Cache_End) begin
            Fsm_nextState = IMG2COL_ENUM_WAIT_COMPUTE;
          end else begin
            Fsm_nextState = IMG2COL_ENUM_DATA_CACHE;
          end
        end
      end
    endcase
  end

  assign when_WaCounter_l19 = ((Fsm_currentState & IMG2COL_ENUM_INIT) != 7'b0000000);
  assign when_WaCounter_l14 = (Init_Count_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l14) begin
      Init_Count_valid = 1'b1;
    end else begin
      Init_Count_valid = 1'b0;
    end
  end

  assign Fsm_Init_End = Init_Count_valid;
  assign when_WaCounter_l40 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign Addr_Init_Cnt_valid = ((Addr_Init_Cnt_count == _zz_Addr_Init_Cnt_valid) && when_WaCounter_l40);
  assign Fsm_Addr_Inited = Addr_Init_Cnt_valid;
  always @(*) begin
    AddrFifo_io_push_valid = 1'b0;
    if(when_Data_Generate_V2_l170) begin
      AddrFifo_io_push_valid = 1'b1;
    end
    if(In_Col_Cnt_valid) begin
      AddrFifo_io_push_valid = 1'b1;
    end
  end

  always @(*) begin
    AddrFifo_io_pop_ready = 1'b0;
    if(when_Data_Generate_V2_l183) begin
      AddrFifo_io_pop_ready = 1'b1;
    end
    if(In_Col_Cnt_valid) begin
      AddrFifo_io_pop_ready = 1'b1;
    end
  end

  assign when_Data_Generate_V2_l170 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign when_Data_Generate_V2_l175 = ((Fsm_currentState & IMG2COL_ENUM_INIT) != 7'b0000000);
  assign SubModule_AddrFifo_io_pop_fire = (AddrFifo_io_pop_valid && AddrFifo_io_pop_ready);
  assign when_Data_Generate_V2_l179 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign when_Data_Generate_V2_l183 = (((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000) && ((Fsm_nextState & IMG2COL_ENUM_DATA_CACHE) != 7'b0000000));
  always @(*) begin
    RaddrFifo0_io_push_valid = 1'b0;
    if(when_Data_Generate_V2_l193) begin
      RaddrFifo0_io_push_valid = 1'b1;
    end
    if(when_Data_Generate_V2_l245) begin
      RaddrFifo0_io_push_valid = SubModule_RaddrFifo0_io_pop_fire;
    end
  end

  always @(*) begin
    RaddrFifo0_io_pop_ready = 1'b0;
    if(when_Data_Generate_V2_l245) begin
      RaddrFifo0_io_pop_ready = Img2ColOutput_Module_Ready_Receive_Addr;
    end
  end

  always @(*) begin
    RaddrFifo0_io_push_payload = RaddrFifo0_io_pop_payload;
    if(when_Data_Generate_V2_l193) begin
      RaddrFifo0_io_push_payload = Raddr_Initialization;
    end
    if(when_Data_Generate_V2_l245) begin
      RaddrFifo0_io_push_payload = RaddrFifo0_io_pop_payload;
    end
  end

  assign when_Data_Generate_V2_l193 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign when_Data_Generate_V2_l197 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign sData_fire = (sData_valid && sData_ready);
  assign In_Col_Cnt_valid = ((In_Col_Cnt_count == _zz_In_Col_Cnt_valid) && sData_fire);
  assign Row_Cache_Cnt_valid = ((Row_Cache_Cnt_count == _zz_Row_Cache_Cnt_valid) && In_Col_Cnt_valid);
  assign In_Row_Cnt_valid = ((In_Row_Cnt_count == _zz_In_Row_Cnt_valid) && In_Col_Cnt_valid);
  assign when_Data_Generate_V2_l217 = (_zz_when_Data_Generate_V2_l217 < In_Row_Cnt_count);
  always @(*) begin
    if(when_Data_Generate_V2_l217) begin
      Cache_Row_Num = Stride;
    end else begin
      Cache_Row_Num = Kernel_Size;
    end
  end

  always @(*) begin
    if(when_Data_Generate_V2_l217) begin
      Raddr_Updata_Cnt_Num = Stride;
    end else begin
      Raddr_Updata_Cnt_Num = Kernel_Size;
    end
  end

  assign Fsm_Data_Cached = Row_Cache_Cnt_valid;
  assign when_Data_Generate_V2_l228 = ((Fsm_currentState & IMG2COL_ENUM_IDLE) != 7'b0000000);
  assign Fsm_Cache_End = CacheEnd_Flag;
  assign sData_ready = ((Fsm_currentState & IMG2COL_ENUM_DATA_CACHE) != 7'b0000000);
  assign when_Data_Generate_V2_l245 = ((Fsm_currentState & IMG2COL_ENUM_UPDATE_ADDR) != 7'b0000000);
  assign SubModule_RaddrFifo0_io_pop_fire = (RaddrFifo0_io_pop_valid && RaddrFifo0_io_pop_ready);
  assign Img2Col_SubModule_start = ((Fsm_currentState & IMG2COL_ENUM_UPDATE_ADDR) != 7'b0000000);
  assign Fsm_SA_Ready = Img2Col_SubModule_SA_Idle;
  assign Img2ColOutput_Module_Ready_Receive_Addr = Img2Col_SubModule_NewAddrIn_ready;
  assign Img2Col_SubModule_NewAddrIn_valid = ((Fsm_currentState & IMG2COL_ENUM_UPDATE_ADDR) != 7'b0000000);
  assign SA_Row_Cnt_Valid = Img2Col_SubModule_SA_Row_Cnt_Valid;
  assign LayerEnd = Fsm_Layer_End;
  assign Fsm_Addr_Updated = Img2Col_SubModule_AddrReceived;
  assign Out_Row_Cnt_valid = ((Out_Row_Cnt_count == _zz_Out_Row_Cnt_valid) && Img2Col_SubModule_SA_End);
  assign Fsm_Layer_End = Out_Row_Cnt_valid;
  assign Waddr = (WaddrOffset + In_Col_Cnt_count);
  assign DGB_addra = Waddr[13:0];
  assign sData_fire_1 = (sData_valid && sData_ready);
  assign DGB_addrb = Img2Col_SubModule_Raddr[13:0];
  assign mData = DGB_doutb;
  assign mValid = SubModule_Img2Col_SubModule_Raddr_Valid_regNext;
  assign mLast = Out_Row_Cnt_valid_regNext;
  assign Test_Valid = (_zz_Test_Valid == Out_Row_Cnt_count_regNext);
  assign Test_Signal = Test_Valid;
  assign Test_End = ((! Test_Valid) && Test_Valid_regNext);
  assign AddrFifo_io_flush = ((Fsm_nextState & IMG2COL_ENUM_IDLE) != 7'b0000000);
  assign RaddrFifo0_io_flush = ((Fsm_nextState & IMG2COL_ENUM_IDLE) != 7'b0000000);
  assign Raddr_Valid = Img2Col_SubModule_Raddr_Valid;
  always @(posedge clk) begin
    start_regNext <= start;
    SubModule_Img2Col_SubModule_Raddr_Valid_regNext <= Img2Col_SubModule_Raddr_Valid;
    Out_Row_Cnt_valid_regNext <= Out_Row_Cnt_valid;
    Out_Row_Cnt_count_regNext <= Out_Row_Cnt_count;
    Test_Valid_regNext <= Test_Valid;
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= IMG2COL_ENUM_IDLE;
      Init_Count_count <= 3'b000;
      Addr_Init_Cnt_count <= 5'h0;
      WaddrOffset <= 16'h0;
      Raddr_Initialization <= 16'h0;
      In_Col_Cnt_count <= 16'h0;
      Row_Cache_Cnt_count <= 5'h0;
      In_Row_Cnt_count <= 16'h0;
      CacheEnd_Flag <= 1'b0;
      Out_Row_Cnt_count <= 16'h0;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l19) begin
        Init_Count_count <= (Init_Count_count + 3'b001);
        if(Init_Count_valid) begin
          Init_Count_count <= 3'b000;
        end
      end
      if(when_WaCounter_l40) begin
        if(Addr_Init_Cnt_valid) begin
          Addr_Init_Cnt_count <= 5'h0;
        end else begin
          Addr_Init_Cnt_count <= (Addr_Init_Cnt_count + 5'h01);
        end
      end
      if(when_Data_Generate_V2_l175) begin
        WaddrOffset <= 16'h0;
      end else begin
        if(SubModule_AddrFifo_io_pop_fire) begin
          WaddrOffset <= AddrFifo_io_pop_payload;
        end else begin
          if(when_Data_Generate_V2_l179) begin
            WaddrOffset <= (WaddrOffset + InCol_Count_Times);
          end
        end
      end
      if(when_Data_Generate_V2_l197) begin
        Raddr_Initialization <= (Raddr_Initialization + InCol_Count_Times);
      end else begin
        Raddr_Initialization <= 16'h0;
      end
      if(sData_fire) begin
        if(In_Col_Cnt_valid) begin
          In_Col_Cnt_count <= 16'h0;
        end else begin
          In_Col_Cnt_count <= (In_Col_Cnt_count + 16'h0001);
        end
      end
      if(In_Col_Cnt_valid) begin
        if(Row_Cache_Cnt_valid) begin
          Row_Cache_Cnt_count <= 5'h0;
        end else begin
          Row_Cache_Cnt_count <= (Row_Cache_Cnt_count + 5'h01);
        end
      end
      if(In_Col_Cnt_valid) begin
        if(In_Row_Cnt_valid) begin
          In_Row_Cnt_count <= 16'h0;
        end else begin
          In_Row_Cnt_count <= (In_Row_Cnt_count + 16'h0001);
        end
      end
      if(In_Row_Cnt_valid) begin
        CacheEnd_Flag <= 1'b1;
      end else begin
        if(when_Data_Generate_V2_l228) begin
          CacheEnd_Flag <= 1'b0;
        end
      end
      if(Img2Col_SubModule_SA_End) begin
        if(Out_Row_Cnt_valid) begin
          Out_Row_Cnt_count <= 16'h0;
        end else begin
          Out_Row_Cnt_count <= (Out_Row_Cnt_count + 16'h0001);
        end
      end
    end
  end


endmodule

//PE_63 replaced by PE_448

//PE_62 replaced by PE_448

//PE_61 replaced by PE_448

//PE_60 replaced by PE_448

//PE_59 replaced by PE_448

//PE_58 replaced by PE_448

//PE_57 replaced by PE_448

//PE_56 replaced by PE_448

//PE_55 replaced by PE_448

//PE_54 replaced by PE_448

//PE_53 replaced by PE_448

//PE_52 replaced by PE_448

//PE_51 replaced by PE_448

//PE_50 replaced by PE_448

//PE_49 replaced by PE_448

//PE_48 replaced by PE_448

//PE_47 replaced by PE_448

//PE_46 replaced by PE_448

//PE_45 replaced by PE_448

//PE_44 replaced by PE_448

//PE_43 replaced by PE_448

//PE_42 replaced by PE_448

//PE_41 replaced by PE_448

//PE_40 replaced by PE_448

//PE_39 replaced by PE_448

//PE_38 replaced by PE_448

//PE_37 replaced by PE_448

//PE_36 replaced by PE_448

//PE_35 replaced by PE_448

//PE_34 replaced by PE_448

//PE_33 replaced by PE_448

//PE_32 replaced by PE_448

//PE_31 replaced by PE_448

//PE_30 replaced by PE_448

//PE_29 replaced by PE_448

//PE_28 replaced by PE_448

//PE_27 replaced by PE_448

//PE_26 replaced by PE_448

//PE_25 replaced by PE_448

//PE_24 replaced by PE_448

//PE_23 replaced by PE_448

//PE_22 replaced by PE_448

//PE_21 replaced by PE_448

//PE_20 replaced by PE_448

//PE_19 replaced by PE_448

//PE_18 replaced by PE_448

//PE_17 replaced by PE_448

//PE_16 replaced by PE_448

//PE_15 replaced by PE_448

//PE_14 replaced by PE_448

//PE_13 replaced by PE_448

//PE_12 replaced by PE_448

//PE_11 replaced by PE_448

//PE_10 replaced by PE_448

//PE_9 replaced by PE_448

//PE_8 replaced by PE_448

//PE_7 replaced by PE_448

//PE_6 replaced by PE_448

//PE_5 replaced by PE_448

//PE_4 replaced by PE_448

//PE_3 replaced by PE_448

//PE_2 replaced by PE_448

//PE_1 replaced by PE_448

//PE replaced by PE_448

//PE_127 replaced by PE_448

//PE_126 replaced by PE_448

//PE_125 replaced by PE_448

//PE_124 replaced by PE_448

//PE_123 replaced by PE_448

//PE_122 replaced by PE_448

//PE_121 replaced by PE_448

//PE_120 replaced by PE_448

//PE_119 replaced by PE_448

//PE_118 replaced by PE_448

//PE_117 replaced by PE_448

//PE_116 replaced by PE_448

//PE_115 replaced by PE_448

//PE_114 replaced by PE_448

//PE_113 replaced by PE_448

//PE_112 replaced by PE_448

//PE_111 replaced by PE_448

//PE_110 replaced by PE_448

//PE_109 replaced by PE_448

//PE_108 replaced by PE_448

//PE_107 replaced by PE_448

//PE_106 replaced by PE_448

//PE_105 replaced by PE_448

//PE_104 replaced by PE_448

//PE_103 replaced by PE_448

//PE_102 replaced by PE_448

//PE_101 replaced by PE_448

//PE_100 replaced by PE_448

//PE_99 replaced by PE_448

//PE_98 replaced by PE_448

//PE_97 replaced by PE_448

//PE_96 replaced by PE_448

//PE_95 replaced by PE_448

//PE_94 replaced by PE_448

//PE_93 replaced by PE_448

//PE_92 replaced by PE_448

//PE_91 replaced by PE_448

//PE_90 replaced by PE_448

//PE_89 replaced by PE_448

//PE_88 replaced by PE_448

//PE_87 replaced by PE_448

//PE_86 replaced by PE_448

//PE_85 replaced by PE_448

//PE_84 replaced by PE_448

//PE_83 replaced by PE_448

//PE_82 replaced by PE_448

//PE_81 replaced by PE_448

//PE_80 replaced by PE_448

//PE_79 replaced by PE_448

//PE_78 replaced by PE_448

//PE_77 replaced by PE_448

//PE_76 replaced by PE_448

//PE_75 replaced by PE_448

//PE_74 replaced by PE_448

//PE_73 replaced by PE_448

//PE_72 replaced by PE_448

//PE_71 replaced by PE_448

//PE_70 replaced by PE_448

//PE_69 replaced by PE_448

//PE_68 replaced by PE_448

//PE_67 replaced by PE_448

//PE_66 replaced by PE_448

//PE_65 replaced by PE_448

//PE_64 replaced by PE_448

//PE_191 replaced by PE_448

//PE_190 replaced by PE_448

//PE_189 replaced by PE_448

//PE_188 replaced by PE_448

//PE_187 replaced by PE_448

//PE_186 replaced by PE_448

//PE_185 replaced by PE_448

//PE_184 replaced by PE_448

//PE_183 replaced by PE_448

//PE_182 replaced by PE_448

//PE_181 replaced by PE_448

//PE_180 replaced by PE_448

//PE_179 replaced by PE_448

//PE_178 replaced by PE_448

//PE_177 replaced by PE_448

//PE_176 replaced by PE_448

//PE_175 replaced by PE_448

//PE_174 replaced by PE_448

//PE_173 replaced by PE_448

//PE_172 replaced by PE_448

//PE_171 replaced by PE_448

//PE_170 replaced by PE_448

//PE_169 replaced by PE_448

//PE_168 replaced by PE_448

//PE_167 replaced by PE_448

//PE_166 replaced by PE_448

//PE_165 replaced by PE_448

//PE_164 replaced by PE_448

//PE_163 replaced by PE_448

//PE_162 replaced by PE_448

//PE_161 replaced by PE_448

//PE_160 replaced by PE_448

//PE_159 replaced by PE_448

//PE_158 replaced by PE_448

//PE_157 replaced by PE_448

//PE_156 replaced by PE_448

//PE_155 replaced by PE_448

//PE_154 replaced by PE_448

//PE_153 replaced by PE_448

//PE_152 replaced by PE_448

//PE_151 replaced by PE_448

//PE_150 replaced by PE_448

//PE_149 replaced by PE_448

//PE_148 replaced by PE_448

//PE_147 replaced by PE_448

//PE_146 replaced by PE_448

//PE_145 replaced by PE_448

//PE_144 replaced by PE_448

//PE_143 replaced by PE_448

//PE_142 replaced by PE_448

//PE_141 replaced by PE_448

//PE_140 replaced by PE_448

//PE_139 replaced by PE_448

//PE_138 replaced by PE_448

//PE_137 replaced by PE_448

//PE_136 replaced by PE_448

//PE_135 replaced by PE_448

//PE_134 replaced by PE_448

//PE_133 replaced by PE_448

//PE_132 replaced by PE_448

//PE_131 replaced by PE_448

//PE_130 replaced by PE_448

//PE_129 replaced by PE_448

//PE_128 replaced by PE_448

//PE_255 replaced by PE_448

//PE_254 replaced by PE_448

//PE_253 replaced by PE_448

//PE_252 replaced by PE_448

//PE_251 replaced by PE_448

//PE_250 replaced by PE_448

//PE_249 replaced by PE_448

//PE_248 replaced by PE_448

//PE_247 replaced by PE_448

//PE_246 replaced by PE_448

//PE_245 replaced by PE_448

//PE_244 replaced by PE_448

//PE_243 replaced by PE_448

//PE_242 replaced by PE_448

//PE_241 replaced by PE_448

//PE_240 replaced by PE_448

//PE_239 replaced by PE_448

//PE_238 replaced by PE_448

//PE_237 replaced by PE_448

//PE_236 replaced by PE_448

//PE_235 replaced by PE_448

//PE_234 replaced by PE_448

//PE_233 replaced by PE_448

//PE_232 replaced by PE_448

//PE_231 replaced by PE_448

//PE_230 replaced by PE_448

//PE_229 replaced by PE_448

//PE_228 replaced by PE_448

//PE_227 replaced by PE_448

//PE_226 replaced by PE_448

//PE_225 replaced by PE_448

//PE_224 replaced by PE_448

//PE_223 replaced by PE_448

//PE_222 replaced by PE_448

//PE_221 replaced by PE_448

//PE_220 replaced by PE_448

//PE_219 replaced by PE_448

//PE_218 replaced by PE_448

//PE_217 replaced by PE_448

//PE_216 replaced by PE_448

//PE_215 replaced by PE_448

//PE_214 replaced by PE_448

//PE_213 replaced by PE_448

//PE_212 replaced by PE_448

//PE_211 replaced by PE_448

//PE_210 replaced by PE_448

//PE_209 replaced by PE_448

//PE_208 replaced by PE_448

//PE_207 replaced by PE_448

//PE_206 replaced by PE_448

//PE_205 replaced by PE_448

//PE_204 replaced by PE_448

//PE_203 replaced by PE_448

//PE_202 replaced by PE_448

//PE_201 replaced by PE_448

//PE_200 replaced by PE_448

//PE_199 replaced by PE_448

//PE_198 replaced by PE_448

//PE_197 replaced by PE_448

//PE_196 replaced by PE_448

//PE_195 replaced by PE_448

//PE_194 replaced by PE_448

//PE_193 replaced by PE_448

//PE_192 replaced by PE_448

//PE_319 replaced by PE_448

//PE_318 replaced by PE_448

//PE_317 replaced by PE_448

//PE_316 replaced by PE_448

//PE_315 replaced by PE_448

//PE_314 replaced by PE_448

//PE_313 replaced by PE_448

//PE_312 replaced by PE_448

//PE_311 replaced by PE_448

//PE_310 replaced by PE_448

//PE_309 replaced by PE_448

//PE_308 replaced by PE_448

//PE_307 replaced by PE_448

//PE_306 replaced by PE_448

//PE_305 replaced by PE_448

//PE_304 replaced by PE_448

//PE_303 replaced by PE_448

//PE_302 replaced by PE_448

//PE_301 replaced by PE_448

//PE_300 replaced by PE_448

//PE_299 replaced by PE_448

//PE_298 replaced by PE_448

//PE_297 replaced by PE_448

//PE_296 replaced by PE_448

//PE_295 replaced by PE_448

//PE_294 replaced by PE_448

//PE_293 replaced by PE_448

//PE_292 replaced by PE_448

//PE_291 replaced by PE_448

//PE_290 replaced by PE_448

//PE_289 replaced by PE_448

//PE_288 replaced by PE_448

//PE_287 replaced by PE_448

//PE_286 replaced by PE_448

//PE_285 replaced by PE_448

//PE_284 replaced by PE_448

//PE_283 replaced by PE_448

//PE_282 replaced by PE_448

//PE_281 replaced by PE_448

//PE_280 replaced by PE_448

//PE_279 replaced by PE_448

//PE_278 replaced by PE_448

//PE_277 replaced by PE_448

//PE_276 replaced by PE_448

//PE_275 replaced by PE_448

//PE_274 replaced by PE_448

//PE_273 replaced by PE_448

//PE_272 replaced by PE_448

//PE_271 replaced by PE_448

//PE_270 replaced by PE_448

//PE_269 replaced by PE_448

//PE_268 replaced by PE_448

//PE_267 replaced by PE_448

//PE_266 replaced by PE_448

//PE_265 replaced by PE_448

//PE_264 replaced by PE_448

//PE_263 replaced by PE_448

//PE_262 replaced by PE_448

//PE_261 replaced by PE_448

//PE_260 replaced by PE_448

//PE_259 replaced by PE_448

//PE_258 replaced by PE_448

//PE_257 replaced by PE_448

//PE_256 replaced by PE_448

//PE_383 replaced by PE_448

//PE_382 replaced by PE_448

//PE_381 replaced by PE_448

//PE_380 replaced by PE_448

//PE_379 replaced by PE_448

//PE_378 replaced by PE_448

//PE_377 replaced by PE_448

//PE_376 replaced by PE_448

//PE_375 replaced by PE_448

//PE_374 replaced by PE_448

//PE_373 replaced by PE_448

//PE_372 replaced by PE_448

//PE_371 replaced by PE_448

//PE_370 replaced by PE_448

//PE_369 replaced by PE_448

//PE_368 replaced by PE_448

//PE_367 replaced by PE_448

//PE_366 replaced by PE_448

//PE_365 replaced by PE_448

//PE_364 replaced by PE_448

//PE_363 replaced by PE_448

//PE_362 replaced by PE_448

//PE_361 replaced by PE_448

//PE_360 replaced by PE_448

//PE_359 replaced by PE_448

//PE_358 replaced by PE_448

//PE_357 replaced by PE_448

//PE_356 replaced by PE_448

//PE_355 replaced by PE_448

//PE_354 replaced by PE_448

//PE_353 replaced by PE_448

//PE_352 replaced by PE_448

//PE_351 replaced by PE_448

//PE_350 replaced by PE_448

//PE_349 replaced by PE_448

//PE_348 replaced by PE_448

//PE_347 replaced by PE_448

//PE_346 replaced by PE_448

//PE_345 replaced by PE_448

//PE_344 replaced by PE_448

//PE_343 replaced by PE_448

//PE_342 replaced by PE_448

//PE_341 replaced by PE_448

//PE_340 replaced by PE_448

//PE_339 replaced by PE_448

//PE_338 replaced by PE_448

//PE_337 replaced by PE_448

//PE_336 replaced by PE_448

//PE_335 replaced by PE_448

//PE_334 replaced by PE_448

//PE_333 replaced by PE_448

//PE_332 replaced by PE_448

//PE_331 replaced by PE_448

//PE_330 replaced by PE_448

//PE_329 replaced by PE_448

//PE_328 replaced by PE_448

//PE_327 replaced by PE_448

//PE_326 replaced by PE_448

//PE_325 replaced by PE_448

//PE_324 replaced by PE_448

//PE_323 replaced by PE_448

//PE_322 replaced by PE_448

//PE_321 replaced by PE_448

//PE_320 replaced by PE_448

//PE_447 replaced by PE_448

//PE_446 replaced by PE_448

//PE_445 replaced by PE_448

//PE_444 replaced by PE_448

//PE_443 replaced by PE_448

//PE_442 replaced by PE_448

//PE_441 replaced by PE_448

//PE_440 replaced by PE_448

//PE_439 replaced by PE_448

//PE_438 replaced by PE_448

//PE_437 replaced by PE_448

//PE_436 replaced by PE_448

//PE_435 replaced by PE_448

//PE_434 replaced by PE_448

//PE_433 replaced by PE_448

//PE_432 replaced by PE_448

//PE_431 replaced by PE_448

//PE_430 replaced by PE_448

//PE_429 replaced by PE_448

//PE_428 replaced by PE_448

//PE_427 replaced by PE_448

//PE_426 replaced by PE_448

//PE_425 replaced by PE_448

//PE_424 replaced by PE_448

//PE_423 replaced by PE_448

//PE_422 replaced by PE_448

//PE_421 replaced by PE_448

//PE_420 replaced by PE_448

//PE_419 replaced by PE_448

//PE_418 replaced by PE_448

//PE_417 replaced by PE_448

//PE_416 replaced by PE_448

//PE_415 replaced by PE_448

//PE_414 replaced by PE_448

//PE_413 replaced by PE_448

//PE_412 replaced by PE_448

//PE_411 replaced by PE_448

//PE_410 replaced by PE_448

//PE_409 replaced by PE_448

//PE_408 replaced by PE_448

//PE_407 replaced by PE_448

//PE_406 replaced by PE_448

//PE_405 replaced by PE_448

//PE_404 replaced by PE_448

//PE_403 replaced by PE_448

//PE_402 replaced by PE_448

//PE_401 replaced by PE_448

//PE_400 replaced by PE_448

//PE_399 replaced by PE_448

//PE_398 replaced by PE_448

//PE_397 replaced by PE_448

//PE_396 replaced by PE_448

//PE_395 replaced by PE_448

//PE_394 replaced by PE_448

//PE_393 replaced by PE_448

//PE_392 replaced by PE_448

//PE_391 replaced by PE_448

//PE_390 replaced by PE_448

//PE_389 replaced by PE_448

//PE_388 replaced by PE_448

//PE_387 replaced by PE_448

//PE_386 replaced by PE_448

//PE_385 replaced by PE_448

//PE_384 replaced by PE_448

//PE_511 replaced by PE_448

//PE_510 replaced by PE_448

//PE_509 replaced by PE_448

//PE_508 replaced by PE_448

//PE_507 replaced by PE_448

//PE_506 replaced by PE_448

//PE_505 replaced by PE_448

//PE_504 replaced by PE_448

//PE_503 replaced by PE_448

//PE_502 replaced by PE_448

//PE_501 replaced by PE_448

//PE_500 replaced by PE_448

//PE_499 replaced by PE_448

//PE_498 replaced by PE_448

//PE_497 replaced by PE_448

//PE_496 replaced by PE_448

//PE_495 replaced by PE_448

//PE_494 replaced by PE_448

//PE_493 replaced by PE_448

//PE_492 replaced by PE_448

//PE_491 replaced by PE_448

//PE_490 replaced by PE_448

//PE_489 replaced by PE_448

//PE_488 replaced by PE_448

//PE_487 replaced by PE_448

//PE_486 replaced by PE_448

//PE_485 replaced by PE_448

//PE_484 replaced by PE_448

//PE_483 replaced by PE_448

//PE_482 replaced by PE_448

//PE_481 replaced by PE_448

//PE_480 replaced by PE_448

//PE_479 replaced by PE_448

//PE_478 replaced by PE_448

//PE_477 replaced by PE_448

//PE_476 replaced by PE_448

//PE_475 replaced by PE_448

//PE_474 replaced by PE_448

//PE_473 replaced by PE_448

//PE_472 replaced by PE_448

//PE_471 replaced by PE_448

//PE_470 replaced by PE_448

//PE_469 replaced by PE_448

//PE_468 replaced by PE_448

//PE_467 replaced by PE_448

//PE_466 replaced by PE_448

//PE_465 replaced by PE_448

//PE_464 replaced by PE_448

//PE_463 replaced by PE_448

//PE_462 replaced by PE_448

//PE_461 replaced by PE_448

//PE_460 replaced by PE_448

//PE_459 replaced by PE_448

//PE_458 replaced by PE_448

//PE_457 replaced by PE_448

//PE_456 replaced by PE_448

//PE_455 replaced by PE_448

//PE_454 replaced by PE_448

//PE_453 replaced by PE_448

//PE_452 replaced by PE_448

//PE_451 replaced by PE_448

//PE_450 replaced by PE_448

//PE_449 replaced by PE_448

module PE_448 (
  input      [7:0]    activate,
  input      [7:0]    weight,
  input               valid,
  input      [15:0]   signCount,
  output     [7:0]    acount,
  output     [7:0]    bcount,
  output reg [31:0]   PE_OUT,
  output              finish,
  input               clk,
  input               reset
);

  wire       [15:0]   dsp_P;
  wire       [31:0]   _zz_reg1;
  wire       [31:0]   _zz_reg1_1;
  wire       [31:0]   _zz_reg1_2;
  reg        [31:0]   reg1;
  reg                 valid_regNext;
  reg                 valid_regNext_regNext;
  reg        [15:0]   finishCnt_count;
  wire                finishCnt_valid;
  reg                 valid_regNext_1;
  reg        [7:0]    activate_regNext;
  reg        [7:0]    weight_regNext;

  assign _zz_reg1 = {{16{dsp_P[15]}}, dsp_P};
  assign _zz_reg1_1 = 32'h0;
  assign _zz_reg1_2 = {{16{dsp_P[15]}}, dsp_P};
  dsp_marco dsp (
    .CLK (clk          ), //i
    .A   (activate[7:0]), //i
    .B   (weight[7:0]  ), //i
    .P   (dsp_P[15:0]  )  //o
  );
  assign finishCnt_valid = ((finishCnt_count == signCount) && valid_regNext_regNext);
  assign finish = finishCnt_valid;
  always @(*) begin
    PE_OUT = 32'h0;
    if(finishCnt_valid) begin
      PE_OUT = reg1;
    end
  end

  assign acount = activate_regNext;
  assign bcount = weight_regNext;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      reg1 <= 32'h0;
      finishCnt_count <= 16'h0;
    end else begin
      if(valid_regNext_regNext) begin
        if(finishCnt_valid) begin
          finishCnt_count <= 16'h0;
        end else begin
          finishCnt_count <= (finishCnt_count + 16'h0001);
        end
      end
      if(finishCnt_valid) begin
        reg1 <= (valid ? _zz_reg1 : _zz_reg1_1);
      end else begin
        if(valid_regNext_1) begin
          reg1 <= ($signed(_zz_reg1_2) + $signed(reg1));
        end
      end
    end
  end

  always @(posedge clk) begin
    valid_regNext <= valid;
    valid_regNext_regNext <= valid_regNext;
    valid_regNext_1 <= valid;
    activate_regNext <= activate;
    weight_regNext <= weight;
  end


endmodule

module Img2Col_OutPut (
  input               start,
  input               NewAddrIn_valid,
  output              NewAddrIn_ready,
  input      [15:0]   NewAddrIn_payload,
  output              SA_Idle,
  output     [15:0]   Raddr,
  output              Raddr_Valid,
  output              SA_End,
  input      [4:0]    Stride,
  input      [4:0]    Kernel_Size,
  input      [15:0]   Window_Size,
  input      [15:0]   InFeature_Size,
  input      [15:0]   InFeature_Channel,
  input      [15:0]   OutFeature_Channel,
  input      [15:0]   OutFeature_Size,
  input      [15:0]   OutCol_Count_Times,
  input      [15:0]   InCol_Count_Times,
  input      [15:0]   OutFeature_Channel_Count_Times,
  input      [12:0]   Sliding_Size,
  input               mReady,
  input               Fifo_Clear,
  output reg          AddrReceived,
  input               LayerEnd,
  output              SA_Row_Cnt_Valid,
  input               clk,
  input               reset
);
  localparam IMG2COL_OUTPUT_ENUM_IDLE = 7'd1;
  localparam IMG2COL_OUTPUT_ENUM_INIT = 7'd2;
  localparam IMG2COL_OUTPUT_ENUM_INIT_ADDR = 7'd4;
  localparam IMG2COL_OUTPUT_ENUM_SA_COMPUTE = 7'd8;
  localparam IMG2COL_OUTPUT_ENUM_UPDATE_ADDR = 7'd16;
  localparam IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY = 7'd32;
  localparam IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR = 7'd64;

  reg                 RaddrFifo1_io_push_valid;
  reg        [15:0]   RaddrFifo1_io_push_payload;
  reg                 RaddrFifo1_io_pop_ready;
  wire                RaddrFifo1_io_flush;
  wire                RaddrFifo1_io_push_ready;
  wire                RaddrFifo1_io_pop_valid;
  wire       [15:0]   RaddrFifo1_io_pop_payload;
  wire       [5:0]    RaddrFifo1_io_occupancy;
  wire       [5:0]    RaddrFifo1_io_availability;
  wire       [4:0]    _zz_Raddr_Init_Cnt_valid;
  wire       [4:0]    _zz_Raddr_Update_Cnt_valid;
  wire       [12:0]   _zz_In_Channel_Process_Cnt_valid;
  wire       [12:0]   _zz_In_Channel_Process_Cnt_valid_1;
  wire       [15:0]   _zz_Window_Col_Cnt_valid;
  wire       [4:0]    _zz_Window_Col_Cnt_valid_1;
  wire       [15:0]   _zz_Window_Row_Cnt_valid;
  wire       [4:0]    _zz_Window_Row_Cnt_valid_1;
  wire       [15:0]   _zz_Out_Channel_Cnt_valid;
  wire       [15:0]   _zz_Out_Col_Cnt_valid;
  wire       [15:0]   _zz_when_Data_Generate_V2_l498;
  wire       [15:0]   _zz_when_Data_Generate_V2_l498_1;
  wire       [15:0]   _zz_WindowSize_Cnt_valid;
  wire       [15:0]   _zz_WindowSize_Cnt_valid_1;
  wire       [31:0]   _zz_Kernel_Base_Addr;
  wire       [15:0]   _zz_Kernel_Base_Addr_1;
  wire       [31:0]   _zz_Kernel_Addr;
  wire       [15:0]   _zz_Kernel_Addr_1;
  wire       [31:0]   _zz_Kernel_Addr_2;
  wire       [31:0]   _zz_Kernel_Addr_3;
  wire       [31:0]   _zz_Kernel_Addr_4;
  wire       [31:0]   _zz_Raddr;
  wire       [31:0]   _zz_Raddr_1;
  reg                 start_regNext;
  wire                when_Data_Generate_V2_l344;
  reg        [6:0]    Fsm_currentState;
  reg        [6:0]    Fsm_nextState;
  wire                Fsm_Init_End;
  wire                Fsm_Addr_Inited;
  wire                Fsm_SA_Computed;
  wire                Fsm_Addr_Updated;
  wire                Fsm_LayerEnd;
  wire                Fsm_NextReady;
  wire                Fsm_Fifo_Clear;
  wire                when_Data_Generate_V2_l376;
  wire                when_WaCounter_l19;
  reg        [2:0]    Init_Count_count;
  reg                 Init_Count_valid;
  wire                when_WaCounter_l14;
  reg        [15:0]   Row_Base_Addr;
  wire                Img2Col_SubModule_RaddrFifo1_io_pop_fire;
  wire                Img2Col_SubModule_RaddrFifo1_io_push_fire;
  wire                when_WaCounter_l40;
  reg        [4:0]    Raddr_Init_Cnt_count;
  wire                Raddr_Init_Cnt_valid;
  wire                Img2Col_SubModule_RaddrFifo1_io_push_fire_1;
  wire                when_WaCounter_l40_1;
  reg        [4:0]    Raddr_Update_Cnt_count;
  wire                Raddr_Update_Cnt_valid;
  wire                when_Data_Generate_V2_l463;
  wire                when_WaCounter_l40_2;
  reg        [2:0]    SA_Row_Cnt_count;
  reg                 SA_Row_Cnt_valid_1;
  reg        [12:0]   In_Channel_Process_Cnt_count;
  wire                In_Channel_Process_Cnt_valid;
  reg        [15:0]   Window_Col_Cnt_count;
  wire                Window_Col_Cnt_valid;
  reg        [15:0]   Window_Row_Cnt_count;
  wire                Window_Row_Cnt_valid;
  reg        [15:0]   Out_Channel_Cnt_count;
  wire                Out_Channel_Cnt_valid;
  reg        [15:0]   Out_Col_Cnt_count;
  wire                Out_Col_Cnt_valid;
  reg        [15:0]   OutFeature_Col_Lefted;
  wire                when_Data_Generate_V2_l495;
  wire                when_Data_Generate_V2_l498;
  reg        [12:0]   WindowSize_Cnt_count;
  wire                WindowSize_Cnt_valid;
  reg        [31:0]   Kernel_Addr;
  reg        [31:0]   Kernel_Base_Addr;
  wire                when_Data_Generate_V2_l523;
  wire                when_Data_Generate_V2_l533;
  wire                Img2Col_SubModule_RaddrFifo1_io_push_fire_2;
  wire                when_Data_Generate_V2_l537;
  `ifndef SYNTHESIS
  reg [119:0] Fsm_currentState_string;
  reg [119:0] Fsm_nextState_string;
  `endif


  assign _zz_Raddr_Init_Cnt_valid = (Kernel_Size - 5'h01);
  assign _zz_Raddr_Update_Cnt_valid = (Stride - 5'h01);
  assign _zz_In_Channel_Process_Cnt_valid = (_zz_In_Channel_Process_Cnt_valid_1 - 13'h0001);
  assign _zz_In_Channel_Process_Cnt_valid_1 = (InFeature_Channel >>> 3);
  assign _zz_Window_Col_Cnt_valid_1 = (Kernel_Size - 5'h01);
  assign _zz_Window_Col_Cnt_valid = {11'd0, _zz_Window_Col_Cnt_valid_1};
  assign _zz_Window_Row_Cnt_valid_1 = (Kernel_Size - 5'h01);
  assign _zz_Window_Row_Cnt_valid = {11'd0, _zz_Window_Row_Cnt_valid_1};
  assign _zz_Out_Channel_Cnt_valid = (OutFeature_Channel_Count_Times - 16'h0001);
  assign _zz_Out_Col_Cnt_valid = (OutCol_Count_Times - 16'h0001);
  assign _zz_when_Data_Generate_V2_l498 = {13'd0, SA_Row_Cnt_count};
  assign _zz_when_Data_Generate_V2_l498_1 = (OutFeature_Col_Lefted - 16'h0001);
  assign _zz_WindowSize_Cnt_valid = {3'd0, WindowSize_Cnt_count};
  assign _zz_WindowSize_Cnt_valid_1 = (Window_Size - 16'h0001);
  assign _zz_Kernel_Base_Addr_1 = ({3'd0,Sliding_Size} <<< 3);
  assign _zz_Kernel_Base_Addr = {16'd0, _zz_Kernel_Base_Addr_1};
  assign _zz_Kernel_Addr_1 = ({3'd0,Sliding_Size} <<< 3);
  assign _zz_Kernel_Addr = {16'd0, _zz_Kernel_Addr_1};
  assign _zz_Kernel_Addr_2 = (Kernel_Base_Addr + _zz_Kernel_Addr_3);
  assign _zz_Kernel_Addr_3 = {19'd0, WindowSize_Cnt_count};
  assign _zz_Kernel_Addr_4 = {19'd0, Sliding_Size};
  assign _zz_Raddr = (Kernel_Addr + _zz_Raddr_1);
  assign _zz_Raddr_1 = {16'd0, Row_Base_Addr};
  WaddrOffset_Fifo_2 RaddrFifo1 (
    .io_push_valid   (RaddrFifo1_io_push_valid        ), //i
    .io_push_ready   (RaddrFifo1_io_push_ready        ), //o
    .io_push_payload (RaddrFifo1_io_push_payload[15:0]), //i
    .io_pop_valid    (RaddrFifo1_io_pop_valid         ), //o
    .io_pop_ready    (RaddrFifo1_io_pop_ready         ), //i
    .io_pop_payload  (RaddrFifo1_io_pop_payload[15:0] ), //o
    .io_flush        (RaddrFifo1_io_flush             ), //i
    .io_occupancy    (RaddrFifo1_io_occupancy[5:0]    ), //o
    .io_availability (RaddrFifo1_io_availability[5:0] ), //o
    .clk             (clk                             ), //i
    .reset           (reset                           )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      IMG2COL_OUTPUT_ENUM_IDLE : Fsm_currentState_string = "IDLE           ";
      IMG2COL_OUTPUT_ENUM_INIT : Fsm_currentState_string = "INIT           ";
      IMG2COL_OUTPUT_ENUM_INIT_ADDR : Fsm_currentState_string = "INIT_ADDR      ";
      IMG2COL_OUTPUT_ENUM_SA_COMPUTE : Fsm_currentState_string = "SA_COMPUTE     ";
      IMG2COL_OUTPUT_ENUM_UPDATE_ADDR : Fsm_currentState_string = "UPDATE_ADDR    ";
      IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY : Fsm_currentState_string = "WAIT_NEXT_READY";
      IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR : Fsm_currentState_string = "WAIT_FIFO_CLEAR";
      default : Fsm_currentState_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      IMG2COL_OUTPUT_ENUM_IDLE : Fsm_nextState_string = "IDLE           ";
      IMG2COL_OUTPUT_ENUM_INIT : Fsm_nextState_string = "INIT           ";
      IMG2COL_OUTPUT_ENUM_INIT_ADDR : Fsm_nextState_string = "INIT_ADDR      ";
      IMG2COL_OUTPUT_ENUM_SA_COMPUTE : Fsm_nextState_string = "SA_COMPUTE     ";
      IMG2COL_OUTPUT_ENUM_UPDATE_ADDR : Fsm_nextState_string = "UPDATE_ADDR    ";
      IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY : Fsm_nextState_string = "WAIT_NEXT_READY";
      IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR : Fsm_nextState_string = "WAIT_FIFO_CLEAR";
      default : Fsm_nextState_string = "???????????????";
    endcase
  end
  `endif

  assign when_Data_Generate_V2_l344 = (start && (! start_regNext));
  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_IDLE) == IMG2COL_OUTPUT_ENUM_IDLE) : begin
        if(when_Data_Generate_V2_l344) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_INIT;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_IDLE;
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_INIT) == IMG2COL_OUTPUT_ENUM_INIT) : begin
        if(Fsm_Init_End) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_INIT_ADDR;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_INIT;
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_INIT_ADDR) == IMG2COL_OUTPUT_ENUM_INIT_ADDR) : begin
        if(Fsm_Addr_Inited) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_INIT_ADDR;
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY) == IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY) : begin
        if(Fsm_NextReady) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_SA_COMPUTE;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY;
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) == IMG2COL_OUTPUT_ENUM_SA_COMPUTE) : begin
        if(Fsm_LayerEnd) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_IDLE;
        end else begin
          if(Fsm_SA_Computed) begin
            Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR;
          end else begin
            if(when_Data_Generate_V2_l376) begin
              Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY;
            end else begin
              Fsm_nextState = IMG2COL_OUTPUT_ENUM_SA_COMPUTE;
            end
          end
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR) == IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR) : begin
        if(Fsm_Fifo_Clear) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_UPDATE_ADDR;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR;
        end
      end
      default : begin
        if(Fsm_Addr_Updated) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_UPDATE_ADDR;
        end
      end
    endcase
  end

  assign when_Data_Generate_V2_l376 = (! Fsm_NextReady);
  assign when_WaCounter_l19 = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT) != 7'b0000000);
  assign when_WaCounter_l14 = (Init_Count_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l14) begin
      Init_Count_valid = 1'b1;
    end else begin
      Init_Count_valid = 1'b0;
    end
  end

  assign Fsm_Init_End = Init_Count_valid;
  assign Fsm_Fifo_Clear = Fifo_Clear;
  assign NewAddrIn_ready = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT_ADDR) != 7'b0000000) || ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 7'b0000000));
  always @(*) begin
    RaddrFifo1_io_push_valid = 1'b0;
    if(when_Data_Generate_V2_l533) begin
      RaddrFifo1_io_push_valid = NewAddrIn_valid;
    end else begin
      if(when_Data_Generate_V2_l537) begin
        RaddrFifo1_io_push_valid = NewAddrIn_valid;
      end else begin
        RaddrFifo1_io_push_valid = Window_Col_Cnt_valid;
      end
    end
  end

  always @(*) begin
    RaddrFifo1_io_pop_ready = 1'b0;
    if(when_Data_Generate_V2_l463) begin
      RaddrFifo1_io_pop_ready = 1'b1;
    end
    if(!when_Data_Generate_V2_l533) begin
      if(when_Data_Generate_V2_l537) begin
        RaddrFifo1_io_pop_ready = Img2Col_SubModule_RaddrFifo1_io_push_fire_2;
      end
    end
    if(Window_Col_Cnt_valid) begin
      RaddrFifo1_io_pop_ready = 1'b1;
    end
  end

  assign Img2Col_SubModule_RaddrFifo1_io_pop_fire = (RaddrFifo1_io_pop_valid && RaddrFifo1_io_pop_ready);
  assign Img2Col_SubModule_RaddrFifo1_io_push_fire = (RaddrFifo1_io_push_valid && RaddrFifo1_io_push_ready);
  assign when_WaCounter_l40 = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT_ADDR) != 7'b0000000) && Img2Col_SubModule_RaddrFifo1_io_push_fire);
  assign Raddr_Init_Cnt_valid = ((Raddr_Init_Cnt_count == _zz_Raddr_Init_Cnt_valid) && when_WaCounter_l40);
  assign Fsm_Addr_Inited = Raddr_Init_Cnt_valid;
  assign Img2Col_SubModule_RaddrFifo1_io_push_fire_1 = (RaddrFifo1_io_push_valid && RaddrFifo1_io_push_ready);
  assign when_WaCounter_l40_1 = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 7'b0000000) && Img2Col_SubModule_RaddrFifo1_io_push_fire_1);
  assign Raddr_Update_Cnt_valid = ((Raddr_Update_Cnt_count == _zz_Raddr_Update_Cnt_valid) && when_WaCounter_l40_1);
  assign Fsm_Addr_Updated = Raddr_Update_Cnt_valid;
  assign Fsm_NextReady = mReady;
  always @(*) begin
    AddrReceived = 1'b0;
    if(when_Data_Generate_V2_l463) begin
      AddrReceived = 1'b1;
    end
  end

  assign when_Data_Generate_V2_l463 = ((((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT_ADDR) != 7'b0000000) && ((Fsm_nextState & IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY) != 7'b0000000)) || (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 7'b0000000) && ((Fsm_nextState & IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY) != 7'b0000000)));
  assign when_WaCounter_l40_2 = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) != 7'b0000000) && mReady);
  always @(*) begin
    SA_Row_Cnt_valid_1 = ((SA_Row_Cnt_count == 3'b111) && when_WaCounter_l40_2);
    if(when_Data_Generate_V2_l498) begin
      SA_Row_Cnt_valid_1 = 1'b1;
    end
  end

  assign SA_Row_Cnt_Valid = SA_Row_Cnt_valid_1;
  assign In_Channel_Process_Cnt_valid = ((In_Channel_Process_Cnt_count == _zz_In_Channel_Process_Cnt_valid) && SA_Row_Cnt_valid_1);
  assign Window_Col_Cnt_valid = ((Window_Col_Cnt_count == _zz_Window_Col_Cnt_valid) && In_Channel_Process_Cnt_valid);
  assign Window_Row_Cnt_valid = ((Window_Row_Cnt_count == _zz_Window_Row_Cnt_valid) && Window_Col_Cnt_valid);
  assign Out_Channel_Cnt_valid = ((Out_Channel_Cnt_count == _zz_Out_Channel_Cnt_valid) && Window_Row_Cnt_valid);
  assign Out_Col_Cnt_valid = ((Out_Col_Cnt_count == _zz_Out_Col_Cnt_valid) && Out_Channel_Cnt_valid);
  assign SA_End = Out_Col_Cnt_valid;
  assign when_Data_Generate_V2_l495 = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT) != 7'b0000000);
  assign when_Data_Generate_V2_l498 = (((_zz_when_Data_Generate_V2_l498 == _zz_when_Data_Generate_V2_l498_1) && mReady) && ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) != 7'b0000000));
  assign WindowSize_Cnt_valid = ((_zz_WindowSize_Cnt_valid == _zz_WindowSize_Cnt_valid_1) && SA_Row_Cnt_valid_1);
  assign when_Data_Generate_V2_l523 = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) != 7'b0000000) && mReady);
  assign Raddr = _zz_Raddr[15:0];
  assign Fsm_SA_Computed = Out_Col_Cnt_valid;
  assign SA_Idle = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_IDLE) != 7'b0000000) || ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 7'b0000000));
  assign when_Data_Generate_V2_l533 = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT_ADDR) != 7'b0000000);
  always @(*) begin
    if(when_Data_Generate_V2_l533) begin
      RaddrFifo1_io_push_payload = NewAddrIn_payload;
    end else begin
      if(when_Data_Generate_V2_l537) begin
        RaddrFifo1_io_push_payload = NewAddrIn_payload;
      end else begin
        RaddrFifo1_io_push_payload = Row_Base_Addr;
      end
    end
  end

  assign Img2Col_SubModule_RaddrFifo1_io_push_fire_2 = (RaddrFifo1_io_push_valid && RaddrFifo1_io_push_ready);
  assign when_Data_Generate_V2_l537 = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 7'b0000000);
  assign Raddr_Valid = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) != 7'b0000000) && mReady);
  assign Fsm_LayerEnd = LayerEnd;
  assign RaddrFifo1_io_flush = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_IDLE) != 7'b0000000);
  always @(posedge clk) begin
    start_regNext <= start;
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= IMG2COL_OUTPUT_ENUM_IDLE;
      Init_Count_count <= 3'b000;
      Row_Base_Addr <= 16'h0;
      Raddr_Init_Cnt_count <= 5'h0;
      Raddr_Update_Cnt_count <= 5'h0;
      SA_Row_Cnt_count <= 3'b000;
      In_Channel_Process_Cnt_count <= 13'h0;
      Window_Col_Cnt_count <= 16'h0;
      Window_Row_Cnt_count <= 16'h0;
      Out_Channel_Cnt_count <= 16'h0;
      Out_Col_Cnt_count <= 16'h0;
      OutFeature_Col_Lefted <= 16'h0;
      WindowSize_Cnt_count <= 13'h0;
      Kernel_Addr <= 32'h0;
      Kernel_Base_Addr <= 32'h0;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l19) begin
        Init_Count_count <= (Init_Count_count + 3'b001);
        if(Init_Count_valid) begin
          Init_Count_count <= 3'b000;
        end
      end
      if(Img2Col_SubModule_RaddrFifo1_io_pop_fire) begin
        Row_Base_Addr <= RaddrFifo1_io_pop_payload;
      end
      if(when_WaCounter_l40) begin
        if(Raddr_Init_Cnt_valid) begin
          Raddr_Init_Cnt_count <= 5'h0;
        end else begin
          Raddr_Init_Cnt_count <= (Raddr_Init_Cnt_count + 5'h01);
        end
      end
      if(when_WaCounter_l40_1) begin
        if(Raddr_Update_Cnt_valid) begin
          Raddr_Update_Cnt_count <= 5'h0;
        end else begin
          Raddr_Update_Cnt_count <= (Raddr_Update_Cnt_count + 5'h01);
        end
      end
      if(when_WaCounter_l40_2) begin
        if(SA_Row_Cnt_valid_1) begin
          SA_Row_Cnt_count <= 3'b000;
        end else begin
          SA_Row_Cnt_count <= (SA_Row_Cnt_count + 3'b001);
        end
      end
      if(SA_Row_Cnt_valid_1) begin
        if(In_Channel_Process_Cnt_valid) begin
          In_Channel_Process_Cnt_count <= 13'h0;
        end else begin
          In_Channel_Process_Cnt_count <= (In_Channel_Process_Cnt_count + 13'h0001);
        end
      end
      if(In_Channel_Process_Cnt_valid) begin
        if(Window_Col_Cnt_valid) begin
          Window_Col_Cnt_count <= 16'h0;
        end else begin
          Window_Col_Cnt_count <= (Window_Col_Cnt_count + 16'h0001);
        end
      end
      if(Window_Col_Cnt_valid) begin
        if(Window_Row_Cnt_valid) begin
          Window_Row_Cnt_count <= 16'h0;
        end else begin
          Window_Row_Cnt_count <= (Window_Row_Cnt_count + 16'h0001);
        end
      end
      if(Window_Row_Cnt_valid) begin
        if(Out_Channel_Cnt_valid) begin
          Out_Channel_Cnt_count <= 16'h0;
        end else begin
          Out_Channel_Cnt_count <= (Out_Channel_Cnt_count + 16'h0001);
        end
      end
      if(Out_Channel_Cnt_valid) begin
        if(Out_Col_Cnt_valid) begin
          Out_Col_Cnt_count <= 16'h0;
        end else begin
          Out_Col_Cnt_count <= (Out_Col_Cnt_count + 16'h0001);
        end
      end
      if(Out_Col_Cnt_valid) begin
        OutFeature_Col_Lefted <= OutFeature_Size;
      end else begin
        if(Out_Channel_Cnt_valid) begin
          OutFeature_Col_Lefted <= (OutFeature_Col_Lefted - 16'h0008);
        end else begin
          if(when_Data_Generate_V2_l495) begin
            OutFeature_Col_Lefted <= OutFeature_Size;
          end
        end
      end
      if(when_Data_Generate_V2_l498) begin
        SA_Row_Cnt_count <= 3'b000;
      end
      if(SA_Row_Cnt_valid_1) begin
        if(WindowSize_Cnt_valid) begin
          WindowSize_Cnt_count <= 13'h0;
        end else begin
          WindowSize_Cnt_count <= (WindowSize_Cnt_count + 13'h0001);
        end
      end
      if(Out_Col_Cnt_valid) begin
        Kernel_Base_Addr <= 32'h0;
      end else begin
        if(Out_Channel_Cnt_valid) begin
          Kernel_Base_Addr <= (Kernel_Base_Addr + _zz_Kernel_Base_Addr);
        end
      end
      if(Out_Col_Cnt_valid) begin
        Kernel_Addr <= 32'h0;
      end else begin
        if(Out_Channel_Cnt_valid) begin
          Kernel_Addr <= (Kernel_Base_Addr + _zz_Kernel_Addr);
        end else begin
          if(Window_Row_Cnt_valid) begin
            Kernel_Addr <= Kernel_Base_Addr;
          end else begin
            if(WindowSize_Cnt_valid) begin
              Kernel_Addr <= Kernel_Base_Addr;
            end else begin
              if(SA_Row_Cnt_valid_1) begin
                Kernel_Addr <= (_zz_Kernel_Addr_2 + 32'h00000001);
              end else begin
                if(when_Data_Generate_V2_l523) begin
                  Kernel_Addr <= (Kernel_Addr + _zz_Kernel_Addr_4);
                end
              end
            end
          end
        end
      end
    end
  end


endmodule

//WaddrOffset_Fifo_1 replaced by WaddrOffset_Fifo_2

//WaddrOffset_Fifo replaced by WaddrOffset_Fifo_2

module WaddrOffset_Fifo_2 (
  input               io_push_valid,
  output              io_push_ready,
  input      [15:0]   io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [15:0]   io_pop_payload,
  input               io_flush,
  output reg [5:0]    io_occupancy,
  output reg [5:0]    io_availability,
  input               clk,
  input               reset
);

  reg        [15:0]   _zz_logic_ram_port0;
  wire       [5:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [5:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [15:0]   _zz_logic_ram_port_1;
  wire       [5:0]    _zz_io_occupancy;
  wire       [5:0]    _zz_io_availability;
  wire       [5:0]    _zz_io_availability_1;
  wire       [5:0]    _zz_io_availability_2;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [5:0]    logic_pushPtr_valueNext;
  reg        [5:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [5:0]    logic_popPtr_valueNext;
  reg        [5:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1122;
  wire       [5:0]    logic_ptrDif;
  reg [15:0] logic_ram [0:32];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {5'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {5'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_occupancy = (6'h21 + logic_ptrDif);
  assign _zz_io_availability = (6'h21 + _zz_io_availability_1);
  assign _zz_io_availability_1 = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_availability_2 = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  assign _zz_logic_ram_port_1 = io_push_payload;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 6'h20);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    if(logic_pushPtr_willOverflow) begin
      logic_pushPtr_valueNext = 6'h0;
    end else begin
      logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    end
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 6'h0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 6'h20);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    if(logic_popPtr_willOverflow) begin
      logic_popPtr_valueNext = 6'h0;
    end else begin
      logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    end
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 6'h0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1122 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  always @(*) begin
    if(logic_ptrMatch) begin
      io_occupancy = (logic_risingOccupancy ? 6'h21 : 6'h0);
    end else begin
      io_occupancy = ((logic_popPtr_value < logic_pushPtr_value) ? logic_ptrDif : _zz_io_occupancy);
    end
  end

  always @(*) begin
    if(logic_ptrMatch) begin
      io_availability = (logic_risingOccupancy ? 6'h0 : 6'h21);
    end else begin
      io_availability = ((logic_popPtr_value < logic_pushPtr_value) ? _zz_io_availability : _zz_io_availability_2);
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_pushPtr_value <= 6'h0;
      logic_popPtr_value <= 6'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1122) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule
