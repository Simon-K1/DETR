// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : AA
// Git hash  : 99c8b6a5c98a226ddc61052be1039b9109e1b352

`timescale 1ns/1ps

module AA (
  input      [0:0]    BB
);



endmodule
