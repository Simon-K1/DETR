// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : MyAxi
// Git hash  : 69cdb32185966f761874d999a3de38a7fe9fad42

`timescale 1ns/1ps

module MyAxi (
  input               io_ACLK,
  input               io_rst,
  input               clk,
  input               reset
);

  wire       [31:0]   aa;

  assign aa = 32'h0;

endmodule
