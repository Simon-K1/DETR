// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : SA_3D
// Git hash  : 993282cd44901a5d48c9a83e85082faf9538d012

`timescale 1ns/1ps

module SA_3D (
  input      [7:0]    _zz_io_MatrixA_0,
  input      [7:0]    _zz_io_MatrixA_1,
  input      [7:0]    _zz_io_MatrixA_2,
  input      [7:0]    _zz_io_MatrixA_3,
  input      [7:0]    _zz_io_MatrixA_4,
  input      [7:0]    _zz_io_MatrixA_5,
  input      [7:0]    _zz_io_MatrixA_6,
  input      [7:0]    _zz_io_MatrixA_7,
  input      [7:0]    _zz_io_MatrixB_0,
  input      [7:0]    _zz_io_MatrixB_1,
  input      [7:0]    _zz_io_MatrixB_2,
  input      [7:0]    _zz_io_MatrixB_3,
  input      [7:0]    _zz_io_MatrixB_4,
  input      [7:0]    _zz_io_MatrixB_5,
  input      [7:0]    _zz_io_MatrixB_6,
  input      [7:0]    _zz_io_MatrixB_7,
  input               _zz_io_A_Valid_0,
  input               _zz_io_A_Valid_1,
  input               _zz_io_A_Valid_2,
  input               _zz_io_A_Valid_3,
  input               _zz_io_A_Valid_4,
  input               _zz_io_A_Valid_5,
  input               _zz_io_A_Valid_6,
  input               _zz_io_A_Valid_7,
  input               _zz_io_B_Valid_0,
  input               _zz_io_B_Valid_1,
  input               _zz_io_B_Valid_2,
  input               _zz_io_B_Valid_3,
  input               _zz_io_B_Valid_4,
  input               _zz_io_B_Valid_5,
  input               _zz_io_B_Valid_6,
  input               _zz_io_B_Valid_7,
  input      [15:0]   _zz_io_signCount,
  input               clk,
  input      [7:0]    _zz_io_MatrixA_0_1,
  input      [7:0]    _zz_io_MatrixA_1_1,
  input      [7:0]    _zz_io_MatrixA_2_1,
  input      [7:0]    _zz_io_MatrixA_3_1,
  input      [7:0]    _zz_io_MatrixA_4_1,
  input      [7:0]    _zz_io_MatrixA_5_1,
  input      [7:0]    _zz_io_MatrixA_6_1,
  input      [7:0]    _zz_io_MatrixA_7_1,
  input      [7:0]    _zz_io_MatrixB_0_1,
  input      [7:0]    _zz_io_MatrixB_1_1,
  input      [7:0]    _zz_io_MatrixB_2_1,
  input      [7:0]    _zz_io_MatrixB_3_1,
  input      [7:0]    _zz_io_MatrixB_4_1,
  input      [7:0]    _zz_io_MatrixB_5_1,
  input      [7:0]    _zz_io_MatrixB_6_1,
  input      [7:0]    _zz_io_MatrixB_7_1,
  input               _zz_io_A_Valid_0_1,
  input               _zz_io_A_Valid_1_1,
  input               _zz_io_A_Valid_2_1,
  input               _zz_io_A_Valid_3_1,
  input               _zz_io_A_Valid_4_1,
  input               _zz_io_A_Valid_5_1,
  input               _zz_io_A_Valid_6_1,
  input               _zz_io_A_Valid_7_1,
  input               _zz_io_B_Valid_0_1,
  input               _zz_io_B_Valid_1_1,
  input               _zz_io_B_Valid_2_1,
  input               _zz_io_B_Valid_3_1,
  input               _zz_io_B_Valid_4_1,
  input               _zz_io_B_Valid_5_1,
  input               _zz_io_B_Valid_6_1,
  input               _zz_io_B_Valid_7_1,
  input      [15:0]   _zz_io_signCount_1,
  input      [7:0]    _zz_io_MatrixA_0_2,
  input      [7:0]    _zz_io_MatrixA_1_2,
  input      [7:0]    _zz_io_MatrixA_2_2,
  input      [7:0]    _zz_io_MatrixA_3_2,
  input      [7:0]    _zz_io_MatrixA_4_2,
  input      [7:0]    _zz_io_MatrixA_5_2,
  input      [7:0]    _zz_io_MatrixA_6_2,
  input      [7:0]    _zz_io_MatrixA_7_2,
  input      [7:0]    _zz_io_MatrixB_0_2,
  input      [7:0]    _zz_io_MatrixB_1_2,
  input      [7:0]    _zz_io_MatrixB_2_2,
  input      [7:0]    _zz_io_MatrixB_3_2,
  input      [7:0]    _zz_io_MatrixB_4_2,
  input      [7:0]    _zz_io_MatrixB_5_2,
  input      [7:0]    _zz_io_MatrixB_6_2,
  input      [7:0]    _zz_io_MatrixB_7_2,
  input               _zz_io_A_Valid_0_2,
  input               _zz_io_A_Valid_1_2,
  input               _zz_io_A_Valid_2_2,
  input               _zz_io_A_Valid_3_2,
  input               _zz_io_A_Valid_4_2,
  input               _zz_io_A_Valid_5_2,
  input               _zz_io_A_Valid_6_2,
  input               _zz_io_A_Valid_7_2,
  input               _zz_io_B_Valid_0_2,
  input               _zz_io_B_Valid_1_2,
  input               _zz_io_B_Valid_2_2,
  input               _zz_io_B_Valid_3_2,
  input               _zz_io_B_Valid_4_2,
  input               _zz_io_B_Valid_5_2,
  input               _zz_io_B_Valid_6_2,
  input               _zz_io_B_Valid_7_2,
  input      [15:0]   _zz_io_signCount_2,
  input      [7:0]    _zz_io_MatrixA_0_3,
  input      [7:0]    _zz_io_MatrixA_1_3,
  input      [7:0]    _zz_io_MatrixA_2_3,
  input      [7:0]    _zz_io_MatrixA_3_3,
  input      [7:0]    _zz_io_MatrixA_4_3,
  input      [7:0]    _zz_io_MatrixA_5_3,
  input      [7:0]    _zz_io_MatrixA_6_3,
  input      [7:0]    _zz_io_MatrixA_7_3,
  input      [7:0]    _zz_io_MatrixB_0_3,
  input      [7:0]    _zz_io_MatrixB_1_3,
  input      [7:0]    _zz_io_MatrixB_2_3,
  input      [7:0]    _zz_io_MatrixB_3_3,
  input      [7:0]    _zz_io_MatrixB_4_3,
  input      [7:0]    _zz_io_MatrixB_5_3,
  input      [7:0]    _zz_io_MatrixB_6_3,
  input      [7:0]    _zz_io_MatrixB_7_3,
  input               _zz_io_A_Valid_0_3,
  input               _zz_io_A_Valid_1_3,
  input               _zz_io_A_Valid_2_3,
  input               _zz_io_A_Valid_3_3,
  input               _zz_io_A_Valid_4_3,
  input               _zz_io_A_Valid_5_3,
  input               _zz_io_A_Valid_6_3,
  input               _zz_io_A_Valid_7_3,
  input               _zz_io_B_Valid_0_3,
  input               _zz_io_B_Valid_1_3,
  input               _zz_io_B_Valid_2_3,
  input               _zz_io_B_Valid_3_3,
  input               _zz_io_B_Valid_4_3,
  input               _zz_io_B_Valid_5_3,
  input               _zz_io_B_Valid_6_3,
  input               _zz_io_B_Valid_7_3,
  input      [15:0]   _zz_io_signCount_3,
  input      [7:0]    _zz_io_MatrixA_0_4,
  input      [7:0]    _zz_io_MatrixA_1_4,
  input      [7:0]    _zz_io_MatrixA_2_4,
  input      [7:0]    _zz_io_MatrixA_3_4,
  input      [7:0]    _zz_io_MatrixA_4_4,
  input      [7:0]    _zz_io_MatrixA_5_4,
  input      [7:0]    _zz_io_MatrixA_6_4,
  input      [7:0]    _zz_io_MatrixA_7_4,
  input      [7:0]    _zz_io_MatrixB_0_4,
  input      [7:0]    _zz_io_MatrixB_1_4,
  input      [7:0]    _zz_io_MatrixB_2_4,
  input      [7:0]    _zz_io_MatrixB_3_4,
  input      [7:0]    _zz_io_MatrixB_4_4,
  input      [7:0]    _zz_io_MatrixB_5_4,
  input      [7:0]    _zz_io_MatrixB_6_4,
  input      [7:0]    _zz_io_MatrixB_7_4,
  input               _zz_io_A_Valid_0_4,
  input               _zz_io_A_Valid_1_4,
  input               _zz_io_A_Valid_2_4,
  input               _zz_io_A_Valid_3_4,
  input               _zz_io_A_Valid_4_4,
  input               _zz_io_A_Valid_5_4,
  input               _zz_io_A_Valid_6_4,
  input               _zz_io_A_Valid_7_4,
  input               _zz_io_B_Valid_0_4,
  input               _zz_io_B_Valid_1_4,
  input               _zz_io_B_Valid_2_4,
  input               _zz_io_B_Valid_3_4,
  input               _zz_io_B_Valid_4_4,
  input               _zz_io_B_Valid_5_4,
  input               _zz_io_B_Valid_6_4,
  input               _zz_io_B_Valid_7_4,
  input      [15:0]   _zz_io_signCount_4,
  input      [7:0]    _zz_io_MatrixA_0_5,
  input      [7:0]    _zz_io_MatrixA_1_5,
  input      [7:0]    _zz_io_MatrixA_2_5,
  input      [7:0]    _zz_io_MatrixA_3_5,
  input      [7:0]    _zz_io_MatrixA_4_5,
  input      [7:0]    _zz_io_MatrixA_5_5,
  input      [7:0]    _zz_io_MatrixA_6_5,
  input      [7:0]    _zz_io_MatrixA_7_5,
  input      [7:0]    _zz_io_MatrixB_0_5,
  input      [7:0]    _zz_io_MatrixB_1_5,
  input      [7:0]    _zz_io_MatrixB_2_5,
  input      [7:0]    _zz_io_MatrixB_3_5,
  input      [7:0]    _zz_io_MatrixB_4_5,
  input      [7:0]    _zz_io_MatrixB_5_5,
  input      [7:0]    _zz_io_MatrixB_6_5,
  input      [7:0]    _zz_io_MatrixB_7_5,
  input               _zz_io_A_Valid_0_5,
  input               _zz_io_A_Valid_1_5,
  input               _zz_io_A_Valid_2_5,
  input               _zz_io_A_Valid_3_5,
  input               _zz_io_A_Valid_4_5,
  input               _zz_io_A_Valid_5_5,
  input               _zz_io_A_Valid_6_5,
  input               _zz_io_A_Valid_7_5,
  input               _zz_io_B_Valid_0_5,
  input               _zz_io_B_Valid_1_5,
  input               _zz_io_B_Valid_2_5,
  input               _zz_io_B_Valid_3_5,
  input               _zz_io_B_Valid_4_5,
  input               _zz_io_B_Valid_5_5,
  input               _zz_io_B_Valid_6_5,
  input               _zz_io_B_Valid_7_5,
  input      [15:0]   _zz_io_signCount_5,
  input      [7:0]    _zz_io_MatrixA_0_6,
  input      [7:0]    _zz_io_MatrixA_1_6,
  input      [7:0]    _zz_io_MatrixA_2_6,
  input      [7:0]    _zz_io_MatrixA_3_6,
  input      [7:0]    _zz_io_MatrixA_4_6,
  input      [7:0]    _zz_io_MatrixA_5_6,
  input      [7:0]    _zz_io_MatrixA_6_6,
  input      [7:0]    _zz_io_MatrixA_7_6,
  input      [7:0]    _zz_io_MatrixB_0_6,
  input      [7:0]    _zz_io_MatrixB_1_6,
  input      [7:0]    _zz_io_MatrixB_2_6,
  input      [7:0]    _zz_io_MatrixB_3_6,
  input      [7:0]    _zz_io_MatrixB_4_6,
  input      [7:0]    _zz_io_MatrixB_5_6,
  input      [7:0]    _zz_io_MatrixB_6_6,
  input      [7:0]    _zz_io_MatrixB_7_6,
  input               _zz_io_A_Valid_0_6,
  input               _zz_io_A_Valid_1_6,
  input               _zz_io_A_Valid_2_6,
  input               _zz_io_A_Valid_3_6,
  input               _zz_io_A_Valid_4_6,
  input               _zz_io_A_Valid_5_6,
  input               _zz_io_A_Valid_6_6,
  input               _zz_io_A_Valid_7_6,
  input               _zz_io_B_Valid_0_6,
  input               _zz_io_B_Valid_1_6,
  input               _zz_io_B_Valid_2_6,
  input               _zz_io_B_Valid_3_6,
  input               _zz_io_B_Valid_4_6,
  input               _zz_io_B_Valid_5_6,
  input               _zz_io_B_Valid_6_6,
  input               _zz_io_B_Valid_7_6,
  input      [15:0]   _zz_io_signCount_6,
  input      [7:0]    _zz_io_MatrixA_0_7,
  input      [7:0]    _zz_io_MatrixA_1_7,
  input      [7:0]    _zz_io_MatrixA_2_7,
  input      [7:0]    _zz_io_MatrixA_3_7,
  input      [7:0]    _zz_io_MatrixA_4_7,
  input      [7:0]    _zz_io_MatrixA_5_7,
  input      [7:0]    _zz_io_MatrixA_6_7,
  input      [7:0]    _zz_io_MatrixA_7_7,
  input      [7:0]    _zz_io_MatrixB_0_7,
  input      [7:0]    _zz_io_MatrixB_1_7,
  input      [7:0]    _zz_io_MatrixB_2_7,
  input      [7:0]    _zz_io_MatrixB_3_7,
  input      [7:0]    _zz_io_MatrixB_4_7,
  input      [7:0]    _zz_io_MatrixB_5_7,
  input      [7:0]    _zz_io_MatrixB_6_7,
  input      [7:0]    _zz_io_MatrixB_7_7,
  input               _zz_io_A_Valid_0_7,
  input               _zz_io_A_Valid_1_7,
  input               _zz_io_A_Valid_2_7,
  input               _zz_io_A_Valid_3_7,
  input               _zz_io_A_Valid_4_7,
  input               _zz_io_A_Valid_5_7,
  input               _zz_io_A_Valid_6_7,
  input               _zz_io_A_Valid_7_7,
  input               _zz_io_B_Valid_0_7,
  input               _zz_io_B_Valid_1_7,
  input               _zz_io_B_Valid_2_7,
  input               _zz_io_B_Valid_3_7,
  input               _zz_io_B_Valid_4_7,
  input               _zz_io_B_Valid_5_7,
  input               _zz_io_B_Valid_6_7,
  input               _zz_io_B_Valid_7_7,
  input      [15:0]   _zz_io_signCount_7,
  input               reset
);

  wire                sA_2D_8_start;
  wire                sA_2D_9_start;
  wire                sA_2D_10_start;
  wire                sA_2D_11_start;
  wire                sA_2D_12_start;
  wire                sA_2D_13_start;
  wire                sA_2D_14_start;
  wire                sA_2D_15_start;
  wire       [31:0]   sA_2D_8_MatrixC_0;
  wire       [31:0]   sA_2D_8_MatrixC_1;
  wire       [31:0]   sA_2D_8_MatrixC_2;
  wire       [31:0]   sA_2D_8_MatrixC_3;
  wire       [31:0]   sA_2D_8_MatrixC_4;
  wire       [31:0]   sA_2D_8_MatrixC_5;
  wire       [31:0]   sA_2D_8_MatrixC_6;
  wire       [31:0]   sA_2D_8_MatrixC_7;
  wire                sA_2D_8_C_Valid_0;
  wire                sA_2D_8_C_Valid_1;
  wire                sA_2D_8_C_Valid_2;
  wire                sA_2D_8_C_Valid_3;
  wire                sA_2D_8_C_Valid_4;
  wire                sA_2D_8_C_Valid_5;
  wire                sA_2D_8_C_Valid_6;
  wire                sA_2D_8_C_Valid_7;
  wire       [31:0]   sA_2D_9_MatrixC_0;
  wire       [31:0]   sA_2D_9_MatrixC_1;
  wire       [31:0]   sA_2D_9_MatrixC_2;
  wire       [31:0]   sA_2D_9_MatrixC_3;
  wire       [31:0]   sA_2D_9_MatrixC_4;
  wire       [31:0]   sA_2D_9_MatrixC_5;
  wire       [31:0]   sA_2D_9_MatrixC_6;
  wire       [31:0]   sA_2D_9_MatrixC_7;
  wire                sA_2D_9_C_Valid_0;
  wire                sA_2D_9_C_Valid_1;
  wire                sA_2D_9_C_Valid_2;
  wire                sA_2D_9_C_Valid_3;
  wire                sA_2D_9_C_Valid_4;
  wire                sA_2D_9_C_Valid_5;
  wire                sA_2D_9_C_Valid_6;
  wire                sA_2D_9_C_Valid_7;
  wire       [31:0]   sA_2D_10_MatrixC_0;
  wire       [31:0]   sA_2D_10_MatrixC_1;
  wire       [31:0]   sA_2D_10_MatrixC_2;
  wire       [31:0]   sA_2D_10_MatrixC_3;
  wire       [31:0]   sA_2D_10_MatrixC_4;
  wire       [31:0]   sA_2D_10_MatrixC_5;
  wire       [31:0]   sA_2D_10_MatrixC_6;
  wire       [31:0]   sA_2D_10_MatrixC_7;
  wire                sA_2D_10_C_Valid_0;
  wire                sA_2D_10_C_Valid_1;
  wire                sA_2D_10_C_Valid_2;
  wire                sA_2D_10_C_Valid_3;
  wire                sA_2D_10_C_Valid_4;
  wire                sA_2D_10_C_Valid_5;
  wire                sA_2D_10_C_Valid_6;
  wire                sA_2D_10_C_Valid_7;
  wire       [31:0]   sA_2D_11_MatrixC_0;
  wire       [31:0]   sA_2D_11_MatrixC_1;
  wire       [31:0]   sA_2D_11_MatrixC_2;
  wire       [31:0]   sA_2D_11_MatrixC_3;
  wire       [31:0]   sA_2D_11_MatrixC_4;
  wire       [31:0]   sA_2D_11_MatrixC_5;
  wire       [31:0]   sA_2D_11_MatrixC_6;
  wire       [31:0]   sA_2D_11_MatrixC_7;
  wire                sA_2D_11_C_Valid_0;
  wire                sA_2D_11_C_Valid_1;
  wire                sA_2D_11_C_Valid_2;
  wire                sA_2D_11_C_Valid_3;
  wire                sA_2D_11_C_Valid_4;
  wire                sA_2D_11_C_Valid_5;
  wire                sA_2D_11_C_Valid_6;
  wire                sA_2D_11_C_Valid_7;
  wire       [31:0]   sA_2D_12_MatrixC_0;
  wire       [31:0]   sA_2D_12_MatrixC_1;
  wire       [31:0]   sA_2D_12_MatrixC_2;
  wire       [31:0]   sA_2D_12_MatrixC_3;
  wire       [31:0]   sA_2D_12_MatrixC_4;
  wire       [31:0]   sA_2D_12_MatrixC_5;
  wire       [31:0]   sA_2D_12_MatrixC_6;
  wire       [31:0]   sA_2D_12_MatrixC_7;
  wire                sA_2D_12_C_Valid_0;
  wire                sA_2D_12_C_Valid_1;
  wire                sA_2D_12_C_Valid_2;
  wire                sA_2D_12_C_Valid_3;
  wire                sA_2D_12_C_Valid_4;
  wire                sA_2D_12_C_Valid_5;
  wire                sA_2D_12_C_Valid_6;
  wire                sA_2D_12_C_Valid_7;
  wire       [31:0]   sA_2D_13_MatrixC_0;
  wire       [31:0]   sA_2D_13_MatrixC_1;
  wire       [31:0]   sA_2D_13_MatrixC_2;
  wire       [31:0]   sA_2D_13_MatrixC_3;
  wire       [31:0]   sA_2D_13_MatrixC_4;
  wire       [31:0]   sA_2D_13_MatrixC_5;
  wire       [31:0]   sA_2D_13_MatrixC_6;
  wire       [31:0]   sA_2D_13_MatrixC_7;
  wire                sA_2D_13_C_Valid_0;
  wire                sA_2D_13_C_Valid_1;
  wire                sA_2D_13_C_Valid_2;
  wire                sA_2D_13_C_Valid_3;
  wire                sA_2D_13_C_Valid_4;
  wire                sA_2D_13_C_Valid_5;
  wire                sA_2D_13_C_Valid_6;
  wire                sA_2D_13_C_Valid_7;
  wire       [31:0]   sA_2D_14_MatrixC_0;
  wire       [31:0]   sA_2D_14_MatrixC_1;
  wire       [31:0]   sA_2D_14_MatrixC_2;
  wire       [31:0]   sA_2D_14_MatrixC_3;
  wire       [31:0]   sA_2D_14_MatrixC_4;
  wire       [31:0]   sA_2D_14_MatrixC_5;
  wire       [31:0]   sA_2D_14_MatrixC_6;
  wire       [31:0]   sA_2D_14_MatrixC_7;
  wire                sA_2D_14_C_Valid_0;
  wire                sA_2D_14_C_Valid_1;
  wire                sA_2D_14_C_Valid_2;
  wire                sA_2D_14_C_Valid_3;
  wire                sA_2D_14_C_Valid_4;
  wire                sA_2D_14_C_Valid_5;
  wire                sA_2D_14_C_Valid_6;
  wire                sA_2D_14_C_Valid_7;
  wire       [31:0]   sA_2D_15_MatrixC_0;
  wire       [31:0]   sA_2D_15_MatrixC_1;
  wire       [31:0]   sA_2D_15_MatrixC_2;
  wire       [31:0]   sA_2D_15_MatrixC_3;
  wire       [31:0]   sA_2D_15_MatrixC_4;
  wire       [31:0]   sA_2D_15_MatrixC_5;
  wire       [31:0]   sA_2D_15_MatrixC_6;
  wire       [31:0]   sA_2D_15_MatrixC_7;
  wire                sA_2D_15_C_Valid_0;
  wire                sA_2D_15_C_Valid_1;
  wire                sA_2D_15_C_Valid_2;
  wire                sA_2D_15_C_Valid_3;
  wire                sA_2D_15_C_Valid_4;
  wire                sA_2D_15_C_Valid_5;
  wire                sA_2D_15_C_Valid_6;
  wire                sA_2D_15_C_Valid_7;

  SA_2D sA_2D_8 (
    .io_MatrixA_0 (_zz_io_MatrixA_0[7:0]  ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1[7:0]  ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2[7:0]  ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3[7:0]  ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4[7:0]  ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5[7:0]  ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6[7:0]  ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7[7:0]  ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0[7:0]  ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1[7:0]  ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2[7:0]  ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3[7:0]  ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4[7:0]  ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5[7:0]  ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6[7:0]  ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7[7:0]  ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0       ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1       ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2       ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3       ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4       ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5       ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6       ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7       ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0       ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1       ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2       ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3       ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4       ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5       ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6       ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7       ), //i
    .io_signCount (_zz_io_signCount[15:0] ), //i
    .MatrixC_0    (sA_2D_8_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_8_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_8_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_8_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_8_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_8_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_8_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_8_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_8_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_8_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_8_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_8_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_8_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_8_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_8_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_8_C_Valid_7      ), //o
    .start        (sA_2D_8_start          ), //i
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  SA_2D sA_2D_9 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_1[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_1[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_1[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_1[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_1[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_1[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_1[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_1[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_1[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_1[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_1[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_1[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_1[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_1[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_1[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_1[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_1      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_1      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_1      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_1      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_1      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_1      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_1      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_1      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_1      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_1      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_1      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_1      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_1      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_1      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_1      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_1      ), //i
    .io_signCount (_zz_io_signCount_1[15:0]), //i
    .MatrixC_0    (sA_2D_9_MatrixC_0[31:0] ), //o
    .MatrixC_1    (sA_2D_9_MatrixC_1[31:0] ), //o
    .MatrixC_2    (sA_2D_9_MatrixC_2[31:0] ), //o
    .MatrixC_3    (sA_2D_9_MatrixC_3[31:0] ), //o
    .MatrixC_4    (sA_2D_9_MatrixC_4[31:0] ), //o
    .MatrixC_5    (sA_2D_9_MatrixC_5[31:0] ), //o
    .MatrixC_6    (sA_2D_9_MatrixC_6[31:0] ), //o
    .MatrixC_7    (sA_2D_9_MatrixC_7[31:0] ), //o
    .C_Valid_0    (sA_2D_9_C_Valid_0       ), //o
    .C_Valid_1    (sA_2D_9_C_Valid_1       ), //o
    .C_Valid_2    (sA_2D_9_C_Valid_2       ), //o
    .C_Valid_3    (sA_2D_9_C_Valid_3       ), //o
    .C_Valid_4    (sA_2D_9_C_Valid_4       ), //o
    .C_Valid_5    (sA_2D_9_C_Valid_5       ), //o
    .C_Valid_6    (sA_2D_9_C_Valid_6       ), //o
    .C_Valid_7    (sA_2D_9_C_Valid_7       ), //o
    .start        (sA_2D_9_start           ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );
  SA_2D sA_2D_10 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_2[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_2[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_2[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_2[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_2[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_2[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_2[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_2[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_2[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_2[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_2[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_2[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_2[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_2[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_2[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_2[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_2      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_2      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_2      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_2      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_2      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_2      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_2      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_2      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_2      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_2      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_2      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_2      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_2      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_2      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_2      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_2      ), //i
    .io_signCount (_zz_io_signCount_2[15:0]), //i
    .MatrixC_0    (sA_2D_10_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_10_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_10_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_10_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_10_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_10_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_10_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_10_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_10_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_10_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_10_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_10_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_10_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_10_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_10_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_10_C_Valid_7      ), //o
    .start        (sA_2D_10_start          ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );
  SA_2D sA_2D_11 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_3[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_3[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_3[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_3[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_3[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_3[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_3[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_3[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_3[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_3[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_3[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_3[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_3[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_3[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_3[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_3[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_3      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_3      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_3      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_3      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_3      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_3      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_3      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_3      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_3      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_3      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_3      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_3      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_3      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_3      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_3      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_3      ), //i
    .io_signCount (_zz_io_signCount_3[15:0]), //i
    .MatrixC_0    (sA_2D_11_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_11_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_11_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_11_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_11_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_11_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_11_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_11_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_11_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_11_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_11_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_11_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_11_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_11_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_11_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_11_C_Valid_7      ), //o
    .start        (sA_2D_11_start          ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );
  SA_2D sA_2D_12 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_4[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_4[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_4[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_4[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_4[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_4[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_4[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_4[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_4[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_4[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_4[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_4[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_4[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_4[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_4[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_4[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_4      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_4      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_4      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_4      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_4      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_4      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_4      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_4      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_4      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_4      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_4      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_4      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_4      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_4      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_4      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_4      ), //i
    .io_signCount (_zz_io_signCount_4[15:0]), //i
    .MatrixC_0    (sA_2D_12_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_12_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_12_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_12_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_12_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_12_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_12_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_12_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_12_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_12_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_12_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_12_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_12_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_12_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_12_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_12_C_Valid_7      ), //o
    .start        (sA_2D_12_start          ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );
  SA_2D sA_2D_13 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_5[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_5[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_5[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_5[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_5[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_5[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_5[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_5[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_5[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_5[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_5[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_5[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_5[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_5[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_5[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_5[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_5      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_5      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_5      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_5      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_5      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_5      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_5      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_5      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_5      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_5      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_5      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_5      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_5      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_5      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_5      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_5      ), //i
    .io_signCount (_zz_io_signCount_5[15:0]), //i
    .MatrixC_0    (sA_2D_13_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_13_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_13_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_13_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_13_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_13_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_13_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_13_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_13_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_13_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_13_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_13_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_13_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_13_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_13_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_13_C_Valid_7      ), //o
    .start        (sA_2D_13_start          ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );
  SA_2D sA_2D_14 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_6[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_6[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_6[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_6[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_6[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_6[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_6[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_6[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_6[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_6[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_6[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_6[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_6[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_6[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_6[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_6[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_6      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_6      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_6      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_6      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_6      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_6      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_6      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_6      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_6      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_6      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_6      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_6      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_6      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_6      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_6      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_6      ), //i
    .io_signCount (_zz_io_signCount_6[15:0]), //i
    .MatrixC_0    (sA_2D_14_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_14_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_14_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_14_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_14_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_14_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_14_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_14_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_14_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_14_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_14_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_14_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_14_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_14_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_14_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_14_C_Valid_7      ), //o
    .start        (sA_2D_14_start          ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );
  SA_2D sA_2D_15 (
    .io_MatrixA_0 (_zz_io_MatrixA_0_7[7:0] ), //i
    .io_MatrixA_1 (_zz_io_MatrixA_1_7[7:0] ), //i
    .io_MatrixA_2 (_zz_io_MatrixA_2_7[7:0] ), //i
    .io_MatrixA_3 (_zz_io_MatrixA_3_7[7:0] ), //i
    .io_MatrixA_4 (_zz_io_MatrixA_4_7[7:0] ), //i
    .io_MatrixA_5 (_zz_io_MatrixA_5_7[7:0] ), //i
    .io_MatrixA_6 (_zz_io_MatrixA_6_7[7:0] ), //i
    .io_MatrixA_7 (_zz_io_MatrixA_7_7[7:0] ), //i
    .io_MatrixB_0 (_zz_io_MatrixB_0_7[7:0] ), //i
    .io_MatrixB_1 (_zz_io_MatrixB_1_7[7:0] ), //i
    .io_MatrixB_2 (_zz_io_MatrixB_2_7[7:0] ), //i
    .io_MatrixB_3 (_zz_io_MatrixB_3_7[7:0] ), //i
    .io_MatrixB_4 (_zz_io_MatrixB_4_7[7:0] ), //i
    .io_MatrixB_5 (_zz_io_MatrixB_5_7[7:0] ), //i
    .io_MatrixB_6 (_zz_io_MatrixB_6_7[7:0] ), //i
    .io_MatrixB_7 (_zz_io_MatrixB_7_7[7:0] ), //i
    .io_A_Valid_0 (_zz_io_A_Valid_0_7      ), //i
    .io_A_Valid_1 (_zz_io_A_Valid_1_7      ), //i
    .io_A_Valid_2 (_zz_io_A_Valid_2_7      ), //i
    .io_A_Valid_3 (_zz_io_A_Valid_3_7      ), //i
    .io_A_Valid_4 (_zz_io_A_Valid_4_7      ), //i
    .io_A_Valid_5 (_zz_io_A_Valid_5_7      ), //i
    .io_A_Valid_6 (_zz_io_A_Valid_6_7      ), //i
    .io_A_Valid_7 (_zz_io_A_Valid_7_7      ), //i
    .io_B_Valid_0 (_zz_io_B_Valid_0_7      ), //i
    .io_B_Valid_1 (_zz_io_B_Valid_1_7      ), //i
    .io_B_Valid_2 (_zz_io_B_Valid_2_7      ), //i
    .io_B_Valid_3 (_zz_io_B_Valid_3_7      ), //i
    .io_B_Valid_4 (_zz_io_B_Valid_4_7      ), //i
    .io_B_Valid_5 (_zz_io_B_Valid_5_7      ), //i
    .io_B_Valid_6 (_zz_io_B_Valid_6_7      ), //i
    .io_B_Valid_7 (_zz_io_B_Valid_7_7      ), //i
    .io_signCount (_zz_io_signCount_7[15:0]), //i
    .MatrixC_0    (sA_2D_15_MatrixC_0[31:0]), //o
    .MatrixC_1    (sA_2D_15_MatrixC_1[31:0]), //o
    .MatrixC_2    (sA_2D_15_MatrixC_2[31:0]), //o
    .MatrixC_3    (sA_2D_15_MatrixC_3[31:0]), //o
    .MatrixC_4    (sA_2D_15_MatrixC_4[31:0]), //o
    .MatrixC_5    (sA_2D_15_MatrixC_5[31:0]), //o
    .MatrixC_6    (sA_2D_15_MatrixC_6[31:0]), //o
    .MatrixC_7    (sA_2D_15_MatrixC_7[31:0]), //o
    .C_Valid_0    (sA_2D_15_C_Valid_0      ), //o
    .C_Valid_1    (sA_2D_15_C_Valid_1      ), //o
    .C_Valid_2    (sA_2D_15_C_Valid_2      ), //o
    .C_Valid_3    (sA_2D_15_C_Valid_3      ), //o
    .C_Valid_4    (sA_2D_15_C_Valid_4      ), //o
    .C_Valid_5    (sA_2D_15_C_Valid_5      ), //o
    .C_Valid_6    (sA_2D_15_C_Valid_6      ), //o
    .C_Valid_7    (sA_2D_15_C_Valid_7      ), //o
    .start        (sA_2D_15_start          ), //i
    .clk          (clk                     ), //i
    .reset        (reset                   )  //i
  );

endmodule

//SA_2D_7 replaced by SA_2D

//SA_2D_6 replaced by SA_2D

//SA_2D_5 replaced by SA_2D

//SA_2D_4 replaced by SA_2D

//SA_2D_3 replaced by SA_2D

//SA_2D_2 replaced by SA_2D

//SA_2D_1 replaced by SA_2D

module SA_2D (
  input      [7:0]    io_MatrixA_0,
  input      [7:0]    io_MatrixA_1,
  input      [7:0]    io_MatrixA_2,
  input      [7:0]    io_MatrixA_3,
  input      [7:0]    io_MatrixA_4,
  input      [7:0]    io_MatrixA_5,
  input      [7:0]    io_MatrixA_6,
  input      [7:0]    io_MatrixA_7,
  input      [7:0]    io_MatrixB_0,
  input      [7:0]    io_MatrixB_1,
  input      [7:0]    io_MatrixB_2,
  input      [7:0]    io_MatrixB_3,
  input      [7:0]    io_MatrixB_4,
  input      [7:0]    io_MatrixB_5,
  input      [7:0]    io_MatrixB_6,
  input      [7:0]    io_MatrixB_7,
  input               io_A_Valid_0,
  input               io_A_Valid_1,
  input               io_A_Valid_2,
  input               io_A_Valid_3,
  input               io_A_Valid_4,
  input               io_A_Valid_5,
  input               io_A_Valid_6,
  input               io_A_Valid_7,
  input               io_B_Valid_0,
  input               io_B_Valid_1,
  input               io_B_Valid_2,
  input               io_B_Valid_3,
  input               io_B_Valid_4,
  input               io_B_Valid_5,
  input               io_B_Valid_6,
  input               io_B_Valid_7,
  input      [15:0]   io_signCount,
  output reg [31:0]   MatrixC_0,
  output reg [31:0]   MatrixC_1,
  output reg [31:0]   MatrixC_2,
  output reg [31:0]   MatrixC_3,
  output reg [31:0]   MatrixC_4,
  output reg [31:0]   MatrixC_5,
  output reg [31:0]   MatrixC_6,
  output reg [31:0]   MatrixC_7,
  output              C_Valid_0,
  output              C_Valid_1,
  output              C_Valid_2,
  output              C_Valid_3,
  output              C_Valid_4,
  output              C_Valid_5,
  output              C_Valid_6,
  output              C_Valid_7,
  input               start,
  input               clk,
  input               reset
);

  wire                pE_512_valid;
  wire                pE_513_valid;
  wire                pE_514_valid;
  wire                pE_515_valid;
  wire                pE_516_valid;
  wire                pE_517_valid;
  wire                pE_518_valid;
  wire                pE_519_valid;
  wire                pE_520_valid;
  wire                pE_521_valid;
  wire                pE_522_valid;
  wire                pE_523_valid;
  wire                pE_524_valid;
  wire                pE_525_valid;
  wire                pE_526_valid;
  wire                pE_527_valid;
  wire                pE_528_valid;
  wire                pE_529_valid;
  wire                pE_530_valid;
  wire                pE_531_valid;
  wire                pE_532_valid;
  wire                pE_533_valid;
  wire                pE_534_valid;
  wire                pE_535_valid;
  wire                pE_536_valid;
  wire                pE_537_valid;
  wire                pE_538_valid;
  wire                pE_539_valid;
  wire                pE_540_valid;
  wire                pE_541_valid;
  wire                pE_542_valid;
  wire                pE_543_valid;
  wire                pE_544_valid;
  wire                pE_545_valid;
  wire                pE_546_valid;
  wire                pE_547_valid;
  wire                pE_548_valid;
  wire                pE_549_valid;
  wire                pE_550_valid;
  wire                pE_551_valid;
  wire                pE_552_valid;
  wire                pE_553_valid;
  wire                pE_554_valid;
  wire                pE_555_valid;
  wire                pE_556_valid;
  wire                pE_557_valid;
  wire                pE_558_valid;
  wire                pE_559_valid;
  wire                pE_560_valid;
  wire                pE_561_valid;
  wire                pE_562_valid;
  wire                pE_563_valid;
  wire                pE_564_valid;
  wire                pE_565_valid;
  wire                pE_566_valid;
  wire                pE_567_valid;
  wire                pE_568_valid;
  wire                pE_569_valid;
  wire                pE_570_valid;
  wire                pE_571_valid;
  wire                pE_572_valid;
  wire                pE_573_valid;
  wire                pE_574_valid;
  wire                pE_575_valid;
  wire       [7:0]    pE_512_acount;
  wire       [7:0]    pE_512_bcount;
  wire       [31:0]   pE_512_PE_OUT;
  wire                pE_512_finish;
  wire       [7:0]    pE_513_acount;
  wire       [7:0]    pE_513_bcount;
  wire       [31:0]   pE_513_PE_OUT;
  wire                pE_513_finish;
  wire       [7:0]    pE_514_acount;
  wire       [7:0]    pE_514_bcount;
  wire       [31:0]   pE_514_PE_OUT;
  wire                pE_514_finish;
  wire       [7:0]    pE_515_acount;
  wire       [7:0]    pE_515_bcount;
  wire       [31:0]   pE_515_PE_OUT;
  wire                pE_515_finish;
  wire       [7:0]    pE_516_acount;
  wire       [7:0]    pE_516_bcount;
  wire       [31:0]   pE_516_PE_OUT;
  wire                pE_516_finish;
  wire       [7:0]    pE_517_acount;
  wire       [7:0]    pE_517_bcount;
  wire       [31:0]   pE_517_PE_OUT;
  wire                pE_517_finish;
  wire       [7:0]    pE_518_acount;
  wire       [7:0]    pE_518_bcount;
  wire       [31:0]   pE_518_PE_OUT;
  wire                pE_518_finish;
  wire       [7:0]    pE_519_acount;
  wire       [7:0]    pE_519_bcount;
  wire       [31:0]   pE_519_PE_OUT;
  wire                pE_519_finish;
  wire       [7:0]    pE_520_acount;
  wire       [7:0]    pE_520_bcount;
  wire       [31:0]   pE_520_PE_OUT;
  wire                pE_520_finish;
  wire       [7:0]    pE_521_acount;
  wire       [7:0]    pE_521_bcount;
  wire       [31:0]   pE_521_PE_OUT;
  wire                pE_521_finish;
  wire       [7:0]    pE_522_acount;
  wire       [7:0]    pE_522_bcount;
  wire       [31:0]   pE_522_PE_OUT;
  wire                pE_522_finish;
  wire       [7:0]    pE_523_acount;
  wire       [7:0]    pE_523_bcount;
  wire       [31:0]   pE_523_PE_OUT;
  wire                pE_523_finish;
  wire       [7:0]    pE_524_acount;
  wire       [7:0]    pE_524_bcount;
  wire       [31:0]   pE_524_PE_OUT;
  wire                pE_524_finish;
  wire       [7:0]    pE_525_acount;
  wire       [7:0]    pE_525_bcount;
  wire       [31:0]   pE_525_PE_OUT;
  wire                pE_525_finish;
  wire       [7:0]    pE_526_acount;
  wire       [7:0]    pE_526_bcount;
  wire       [31:0]   pE_526_PE_OUT;
  wire                pE_526_finish;
  wire       [7:0]    pE_527_acount;
  wire       [7:0]    pE_527_bcount;
  wire       [31:0]   pE_527_PE_OUT;
  wire                pE_527_finish;
  wire       [7:0]    pE_528_acount;
  wire       [7:0]    pE_528_bcount;
  wire       [31:0]   pE_528_PE_OUT;
  wire                pE_528_finish;
  wire       [7:0]    pE_529_acount;
  wire       [7:0]    pE_529_bcount;
  wire       [31:0]   pE_529_PE_OUT;
  wire                pE_529_finish;
  wire       [7:0]    pE_530_acount;
  wire       [7:0]    pE_530_bcount;
  wire       [31:0]   pE_530_PE_OUT;
  wire                pE_530_finish;
  wire       [7:0]    pE_531_acount;
  wire       [7:0]    pE_531_bcount;
  wire       [31:0]   pE_531_PE_OUT;
  wire                pE_531_finish;
  wire       [7:0]    pE_532_acount;
  wire       [7:0]    pE_532_bcount;
  wire       [31:0]   pE_532_PE_OUT;
  wire                pE_532_finish;
  wire       [7:0]    pE_533_acount;
  wire       [7:0]    pE_533_bcount;
  wire       [31:0]   pE_533_PE_OUT;
  wire                pE_533_finish;
  wire       [7:0]    pE_534_acount;
  wire       [7:0]    pE_534_bcount;
  wire       [31:0]   pE_534_PE_OUT;
  wire                pE_534_finish;
  wire       [7:0]    pE_535_acount;
  wire       [7:0]    pE_535_bcount;
  wire       [31:0]   pE_535_PE_OUT;
  wire                pE_535_finish;
  wire       [7:0]    pE_536_acount;
  wire       [7:0]    pE_536_bcount;
  wire       [31:0]   pE_536_PE_OUT;
  wire                pE_536_finish;
  wire       [7:0]    pE_537_acount;
  wire       [7:0]    pE_537_bcount;
  wire       [31:0]   pE_537_PE_OUT;
  wire                pE_537_finish;
  wire       [7:0]    pE_538_acount;
  wire       [7:0]    pE_538_bcount;
  wire       [31:0]   pE_538_PE_OUT;
  wire                pE_538_finish;
  wire       [7:0]    pE_539_acount;
  wire       [7:0]    pE_539_bcount;
  wire       [31:0]   pE_539_PE_OUT;
  wire                pE_539_finish;
  wire       [7:0]    pE_540_acount;
  wire       [7:0]    pE_540_bcount;
  wire       [31:0]   pE_540_PE_OUT;
  wire                pE_540_finish;
  wire       [7:0]    pE_541_acount;
  wire       [7:0]    pE_541_bcount;
  wire       [31:0]   pE_541_PE_OUT;
  wire                pE_541_finish;
  wire       [7:0]    pE_542_acount;
  wire       [7:0]    pE_542_bcount;
  wire       [31:0]   pE_542_PE_OUT;
  wire                pE_542_finish;
  wire       [7:0]    pE_543_acount;
  wire       [7:0]    pE_543_bcount;
  wire       [31:0]   pE_543_PE_OUT;
  wire                pE_543_finish;
  wire       [7:0]    pE_544_acount;
  wire       [7:0]    pE_544_bcount;
  wire       [31:0]   pE_544_PE_OUT;
  wire                pE_544_finish;
  wire       [7:0]    pE_545_acount;
  wire       [7:0]    pE_545_bcount;
  wire       [31:0]   pE_545_PE_OUT;
  wire                pE_545_finish;
  wire       [7:0]    pE_546_acount;
  wire       [7:0]    pE_546_bcount;
  wire       [31:0]   pE_546_PE_OUT;
  wire                pE_546_finish;
  wire       [7:0]    pE_547_acount;
  wire       [7:0]    pE_547_bcount;
  wire       [31:0]   pE_547_PE_OUT;
  wire                pE_547_finish;
  wire       [7:0]    pE_548_acount;
  wire       [7:0]    pE_548_bcount;
  wire       [31:0]   pE_548_PE_OUT;
  wire                pE_548_finish;
  wire       [7:0]    pE_549_acount;
  wire       [7:0]    pE_549_bcount;
  wire       [31:0]   pE_549_PE_OUT;
  wire                pE_549_finish;
  wire       [7:0]    pE_550_acount;
  wire       [7:0]    pE_550_bcount;
  wire       [31:0]   pE_550_PE_OUT;
  wire                pE_550_finish;
  wire       [7:0]    pE_551_acount;
  wire       [7:0]    pE_551_bcount;
  wire       [31:0]   pE_551_PE_OUT;
  wire                pE_551_finish;
  wire       [7:0]    pE_552_acount;
  wire       [7:0]    pE_552_bcount;
  wire       [31:0]   pE_552_PE_OUT;
  wire                pE_552_finish;
  wire       [7:0]    pE_553_acount;
  wire       [7:0]    pE_553_bcount;
  wire       [31:0]   pE_553_PE_OUT;
  wire                pE_553_finish;
  wire       [7:0]    pE_554_acount;
  wire       [7:0]    pE_554_bcount;
  wire       [31:0]   pE_554_PE_OUT;
  wire                pE_554_finish;
  wire       [7:0]    pE_555_acount;
  wire       [7:0]    pE_555_bcount;
  wire       [31:0]   pE_555_PE_OUT;
  wire                pE_555_finish;
  wire       [7:0]    pE_556_acount;
  wire       [7:0]    pE_556_bcount;
  wire       [31:0]   pE_556_PE_OUT;
  wire                pE_556_finish;
  wire       [7:0]    pE_557_acount;
  wire       [7:0]    pE_557_bcount;
  wire       [31:0]   pE_557_PE_OUT;
  wire                pE_557_finish;
  wire       [7:0]    pE_558_acount;
  wire       [7:0]    pE_558_bcount;
  wire       [31:0]   pE_558_PE_OUT;
  wire                pE_558_finish;
  wire       [7:0]    pE_559_acount;
  wire       [7:0]    pE_559_bcount;
  wire       [31:0]   pE_559_PE_OUT;
  wire                pE_559_finish;
  wire       [7:0]    pE_560_acount;
  wire       [7:0]    pE_560_bcount;
  wire       [31:0]   pE_560_PE_OUT;
  wire                pE_560_finish;
  wire       [7:0]    pE_561_acount;
  wire       [7:0]    pE_561_bcount;
  wire       [31:0]   pE_561_PE_OUT;
  wire                pE_561_finish;
  wire       [7:0]    pE_562_acount;
  wire       [7:0]    pE_562_bcount;
  wire       [31:0]   pE_562_PE_OUT;
  wire                pE_562_finish;
  wire       [7:0]    pE_563_acount;
  wire       [7:0]    pE_563_bcount;
  wire       [31:0]   pE_563_PE_OUT;
  wire                pE_563_finish;
  wire       [7:0]    pE_564_acount;
  wire       [7:0]    pE_564_bcount;
  wire       [31:0]   pE_564_PE_OUT;
  wire                pE_564_finish;
  wire       [7:0]    pE_565_acount;
  wire       [7:0]    pE_565_bcount;
  wire       [31:0]   pE_565_PE_OUT;
  wire                pE_565_finish;
  wire       [7:0]    pE_566_acount;
  wire       [7:0]    pE_566_bcount;
  wire       [31:0]   pE_566_PE_OUT;
  wire                pE_566_finish;
  wire       [7:0]    pE_567_acount;
  wire       [7:0]    pE_567_bcount;
  wire       [31:0]   pE_567_PE_OUT;
  wire                pE_567_finish;
  wire       [7:0]    pE_568_acount;
  wire       [7:0]    pE_568_bcount;
  wire       [31:0]   pE_568_PE_OUT;
  wire                pE_568_finish;
  wire       [7:0]    pE_569_acount;
  wire       [7:0]    pE_569_bcount;
  wire       [31:0]   pE_569_PE_OUT;
  wire                pE_569_finish;
  wire       [7:0]    pE_570_acount;
  wire       [7:0]    pE_570_bcount;
  wire       [31:0]   pE_570_PE_OUT;
  wire                pE_570_finish;
  wire       [7:0]    pE_571_acount;
  wire       [7:0]    pE_571_bcount;
  wire       [31:0]   pE_571_PE_OUT;
  wire                pE_571_finish;
  wire       [7:0]    pE_572_acount;
  wire       [7:0]    pE_572_bcount;
  wire       [31:0]   pE_572_PE_OUT;
  wire                pE_572_finish;
  wire       [7:0]    pE_573_acount;
  wire       [7:0]    pE_573_bcount;
  wire       [31:0]   pE_573_PE_OUT;
  wire                pE_573_finish;
  wire       [7:0]    pE_574_acount;
  wire       [7:0]    pE_574_bcount;
  wire       [31:0]   pE_574_PE_OUT;
  wire                pE_574_finish;
  wire       [7:0]    pE_575_acount;
  wire       [7:0]    pE_575_bcount;
  wire       [31:0]   pE_575_PE_OUT;
  wire                pE_575_finish;
  reg        [7:0]    tmp;
  wire                when_SA_3D_l80;
  wire                when_SA_3D_l80_1;
  wire                when_SA_3D_l80_2;
  wire                when_SA_3D_l80_3;
  wire                when_SA_3D_l80_4;
  wire                when_SA_3D_l80_5;
  wire                when_SA_3D_l80_6;
  wire                when_SA_3D_l80_7;
  wire                when_SA_3D_l80_8;
  wire                when_SA_3D_l80_9;
  wire                when_SA_3D_l80_10;
  wire                when_SA_3D_l80_11;
  wire                when_SA_3D_l80_12;
  wire                when_SA_3D_l80_13;
  wire                when_SA_3D_l80_14;
  wire                when_SA_3D_l80_15;
  wire                when_SA_3D_l80_16;
  wire                when_SA_3D_l80_17;
  wire                when_SA_3D_l80_18;
  wire                when_SA_3D_l80_19;
  wire                when_SA_3D_l80_20;
  wire                when_SA_3D_l80_21;
  wire                when_SA_3D_l80_22;
  wire                when_SA_3D_l80_23;
  wire                when_SA_3D_l80_24;
  wire                when_SA_3D_l80_25;
  wire                when_SA_3D_l80_26;
  wire                when_SA_3D_l80_27;
  wire                when_SA_3D_l80_28;
  wire                when_SA_3D_l80_29;
  wire                when_SA_3D_l80_30;
  wire                when_SA_3D_l80_31;
  wire                when_SA_3D_l80_32;
  wire                when_SA_3D_l80_33;
  wire                when_SA_3D_l80_34;
  wire                when_SA_3D_l80_35;
  wire                when_SA_3D_l80_36;
  wire                when_SA_3D_l80_37;
  wire                when_SA_3D_l80_38;
  wire                when_SA_3D_l80_39;
  wire                when_SA_3D_l80_40;
  wire                when_SA_3D_l80_41;
  wire                when_SA_3D_l80_42;
  wire                when_SA_3D_l80_43;
  wire                when_SA_3D_l80_44;
  wire                when_SA_3D_l80_45;
  wire                when_SA_3D_l80_46;
  wire                when_SA_3D_l80_47;
  wire                when_SA_3D_l80_48;
  wire                when_SA_3D_l80_49;
  wire                when_SA_3D_l80_50;
  wire                when_SA_3D_l80_51;
  wire                when_SA_3D_l80_52;
  wire                when_SA_3D_l80_53;
  wire                when_SA_3D_l80_54;
  wire                when_SA_3D_l80_55;
  wire                when_SA_3D_l80_56;
  wire                when_SA_3D_l80_57;
  wire                when_SA_3D_l80_58;
  wire                when_SA_3D_l80_59;
  wire                when_SA_3D_l80_60;
  wire                when_SA_3D_l80_61;
  wire                when_SA_3D_l80_62;
  wire                when_SA_3D_l80_63;
  reg        [15:0]   io_signCount_regNextWhen;
  reg                 io_A_Valid_0_delay_1;
  reg                 io_A_Valid_0_delay_1_1;
  reg                 io_A_Valid_0_delay_2;
  reg                 io_A_Valid_0_delay_1_2;
  reg                 io_A_Valid_0_delay_2_1;
  reg                 io_A_Valid_0_delay_3;
  reg                 io_A_Valid_0_delay_1_3;
  reg                 io_A_Valid_0_delay_2_2;
  reg                 io_A_Valid_0_delay_3_1;
  reg                 io_A_Valid_0_delay_4;
  reg                 io_A_Valid_0_delay_1_4;
  reg                 io_A_Valid_0_delay_2_3;
  reg                 io_A_Valid_0_delay_3_2;
  reg                 io_A_Valid_0_delay_4_1;
  reg                 io_A_Valid_0_delay_5;
  reg                 io_A_Valid_0_delay_1_5;
  reg                 io_A_Valid_0_delay_2_4;
  reg                 io_A_Valid_0_delay_3_3;
  reg                 io_A_Valid_0_delay_4_2;
  reg                 io_A_Valid_0_delay_5_1;
  reg                 io_A_Valid_0_delay_6;
  reg                 io_A_Valid_0_delay_1_6;
  reg                 io_A_Valid_0_delay_2_5;
  reg                 io_A_Valid_0_delay_3_4;
  reg                 io_A_Valid_0_delay_4_3;
  reg                 io_A_Valid_0_delay_5_2;
  reg                 io_A_Valid_0_delay_6_1;
  reg                 io_A_Valid_0_delay_7;
  reg        [15:0]   io_signCount_regNextWhen_1;
  reg                 io_B_Valid_0_delay_1;
  reg                 io_A_Valid_1_delay_1;
  reg                 io_B_Valid_1_delay_1;
  reg                 io_A_Valid_1_delay_1_1;
  reg                 io_A_Valid_1_delay_2;
  reg                 io_B_Valid_2_delay_1;
  reg                 io_A_Valid_1_delay_1_2;
  reg                 io_A_Valid_1_delay_2_1;
  reg                 io_A_Valid_1_delay_3;
  reg                 io_B_Valid_3_delay_1;
  reg                 io_A_Valid_1_delay_1_3;
  reg                 io_A_Valid_1_delay_2_2;
  reg                 io_A_Valid_1_delay_3_1;
  reg                 io_A_Valid_1_delay_4;
  reg                 io_B_Valid_4_delay_1;
  reg                 io_A_Valid_1_delay_1_4;
  reg                 io_A_Valid_1_delay_2_3;
  reg                 io_A_Valid_1_delay_3_2;
  reg                 io_A_Valid_1_delay_4_1;
  reg                 io_A_Valid_1_delay_5;
  reg                 io_B_Valid_5_delay_1;
  reg                 io_A_Valid_1_delay_1_5;
  reg                 io_A_Valid_1_delay_2_4;
  reg                 io_A_Valid_1_delay_3_3;
  reg                 io_A_Valid_1_delay_4_2;
  reg                 io_A_Valid_1_delay_5_1;
  reg                 io_A_Valid_1_delay_6;
  reg                 io_B_Valid_6_delay_1;
  reg                 io_A_Valid_1_delay_1_6;
  reg                 io_A_Valid_1_delay_2_5;
  reg                 io_A_Valid_1_delay_3_4;
  reg                 io_A_Valid_1_delay_4_3;
  reg                 io_A_Valid_1_delay_5_2;
  reg                 io_A_Valid_1_delay_6_1;
  reg                 io_A_Valid_1_delay_7;
  reg                 io_B_Valid_7_delay_1;
  reg        [15:0]   io_signCount_regNextWhen_2;
  reg                 io_B_Valid_0_delay_1_1;
  reg                 io_B_Valid_0_delay_2;
  reg                 io_A_Valid_2_delay_1;
  reg                 io_B_Valid_1_delay_1_1;
  reg                 io_B_Valid_1_delay_2;
  reg                 io_A_Valid_2_delay_1_1;
  reg                 io_A_Valid_2_delay_2;
  reg                 io_B_Valid_2_delay_1_1;
  reg                 io_B_Valid_2_delay_2;
  reg                 io_A_Valid_2_delay_1_2;
  reg                 io_A_Valid_2_delay_2_1;
  reg                 io_A_Valid_2_delay_3;
  reg                 io_B_Valid_3_delay_1_1;
  reg                 io_B_Valid_3_delay_2;
  reg                 io_A_Valid_2_delay_1_3;
  reg                 io_A_Valid_2_delay_2_2;
  reg                 io_A_Valid_2_delay_3_1;
  reg                 io_A_Valid_2_delay_4;
  reg                 io_B_Valid_4_delay_1_1;
  reg                 io_B_Valid_4_delay_2;
  reg                 io_A_Valid_2_delay_1_4;
  reg                 io_A_Valid_2_delay_2_3;
  reg                 io_A_Valid_2_delay_3_2;
  reg                 io_A_Valid_2_delay_4_1;
  reg                 io_A_Valid_2_delay_5;
  reg                 io_B_Valid_5_delay_1_1;
  reg                 io_B_Valid_5_delay_2;
  reg                 io_A_Valid_2_delay_1_5;
  reg                 io_A_Valid_2_delay_2_4;
  reg                 io_A_Valid_2_delay_3_3;
  reg                 io_A_Valid_2_delay_4_2;
  reg                 io_A_Valid_2_delay_5_1;
  reg                 io_A_Valid_2_delay_6;
  reg                 io_B_Valid_6_delay_1_1;
  reg                 io_B_Valid_6_delay_2;
  reg                 io_A_Valid_2_delay_1_6;
  reg                 io_A_Valid_2_delay_2_5;
  reg                 io_A_Valid_2_delay_3_4;
  reg                 io_A_Valid_2_delay_4_3;
  reg                 io_A_Valid_2_delay_5_2;
  reg                 io_A_Valid_2_delay_6_1;
  reg                 io_A_Valid_2_delay_7;
  reg                 io_B_Valid_7_delay_1_1;
  reg                 io_B_Valid_7_delay_2;
  reg        [15:0]   io_signCount_regNextWhen_3;
  reg                 io_B_Valid_0_delay_1_2;
  reg                 io_B_Valid_0_delay_2_1;
  reg                 io_B_Valid_0_delay_3;
  reg                 io_A_Valid_3_delay_1;
  reg                 io_B_Valid_1_delay_1_2;
  reg                 io_B_Valid_1_delay_2_1;
  reg                 io_B_Valid_1_delay_3;
  reg                 io_A_Valid_3_delay_1_1;
  reg                 io_A_Valid_3_delay_2;
  reg                 io_B_Valid_2_delay_1_2;
  reg                 io_B_Valid_2_delay_2_1;
  reg                 io_B_Valid_2_delay_3;
  reg                 io_A_Valid_3_delay_1_2;
  reg                 io_A_Valid_3_delay_2_1;
  reg                 io_A_Valid_3_delay_3;
  reg                 io_B_Valid_3_delay_1_2;
  reg                 io_B_Valid_3_delay_2_1;
  reg                 io_B_Valid_3_delay_3;
  reg                 io_A_Valid_3_delay_1_3;
  reg                 io_A_Valid_3_delay_2_2;
  reg                 io_A_Valid_3_delay_3_1;
  reg                 io_A_Valid_3_delay_4;
  reg                 io_B_Valid_4_delay_1_2;
  reg                 io_B_Valid_4_delay_2_1;
  reg                 io_B_Valid_4_delay_3;
  reg                 io_A_Valid_3_delay_1_4;
  reg                 io_A_Valid_3_delay_2_3;
  reg                 io_A_Valid_3_delay_3_2;
  reg                 io_A_Valid_3_delay_4_1;
  reg                 io_A_Valid_3_delay_5;
  reg                 io_B_Valid_5_delay_1_2;
  reg                 io_B_Valid_5_delay_2_1;
  reg                 io_B_Valid_5_delay_3;
  reg                 io_A_Valid_3_delay_1_5;
  reg                 io_A_Valid_3_delay_2_4;
  reg                 io_A_Valid_3_delay_3_3;
  reg                 io_A_Valid_3_delay_4_2;
  reg                 io_A_Valid_3_delay_5_1;
  reg                 io_A_Valid_3_delay_6;
  reg                 io_B_Valid_6_delay_1_2;
  reg                 io_B_Valid_6_delay_2_1;
  reg                 io_B_Valid_6_delay_3;
  reg                 io_A_Valid_3_delay_1_6;
  reg                 io_A_Valid_3_delay_2_5;
  reg                 io_A_Valid_3_delay_3_4;
  reg                 io_A_Valid_3_delay_4_3;
  reg                 io_A_Valid_3_delay_5_2;
  reg                 io_A_Valid_3_delay_6_1;
  reg                 io_A_Valid_3_delay_7;
  reg                 io_B_Valid_7_delay_1_2;
  reg                 io_B_Valid_7_delay_2_1;
  reg                 io_B_Valid_7_delay_3;
  reg        [15:0]   io_signCount_regNextWhen_4;
  reg                 io_B_Valid_0_delay_1_3;
  reg                 io_B_Valid_0_delay_2_2;
  reg                 io_B_Valid_0_delay_3_1;
  reg                 io_B_Valid_0_delay_4;
  reg                 io_A_Valid_4_delay_1;
  reg                 io_B_Valid_1_delay_1_3;
  reg                 io_B_Valid_1_delay_2_2;
  reg                 io_B_Valid_1_delay_3_1;
  reg                 io_B_Valid_1_delay_4;
  reg                 io_A_Valid_4_delay_1_1;
  reg                 io_A_Valid_4_delay_2;
  reg                 io_B_Valid_2_delay_1_3;
  reg                 io_B_Valid_2_delay_2_2;
  reg                 io_B_Valid_2_delay_3_1;
  reg                 io_B_Valid_2_delay_4;
  reg                 io_A_Valid_4_delay_1_2;
  reg                 io_A_Valid_4_delay_2_1;
  reg                 io_A_Valid_4_delay_3;
  reg                 io_B_Valid_3_delay_1_3;
  reg                 io_B_Valid_3_delay_2_2;
  reg                 io_B_Valid_3_delay_3_1;
  reg                 io_B_Valid_3_delay_4;
  reg                 io_A_Valid_4_delay_1_3;
  reg                 io_A_Valid_4_delay_2_2;
  reg                 io_A_Valid_4_delay_3_1;
  reg                 io_A_Valid_4_delay_4;
  reg                 io_B_Valid_4_delay_1_3;
  reg                 io_B_Valid_4_delay_2_2;
  reg                 io_B_Valid_4_delay_3_1;
  reg                 io_B_Valid_4_delay_4;
  reg                 io_A_Valid_4_delay_1_4;
  reg                 io_A_Valid_4_delay_2_3;
  reg                 io_A_Valid_4_delay_3_2;
  reg                 io_A_Valid_4_delay_4_1;
  reg                 io_A_Valid_4_delay_5;
  reg                 io_B_Valid_5_delay_1_3;
  reg                 io_B_Valid_5_delay_2_2;
  reg                 io_B_Valid_5_delay_3_1;
  reg                 io_B_Valid_5_delay_4;
  reg                 io_A_Valid_4_delay_1_5;
  reg                 io_A_Valid_4_delay_2_4;
  reg                 io_A_Valid_4_delay_3_3;
  reg                 io_A_Valid_4_delay_4_2;
  reg                 io_A_Valid_4_delay_5_1;
  reg                 io_A_Valid_4_delay_6;
  reg                 io_B_Valid_6_delay_1_3;
  reg                 io_B_Valid_6_delay_2_2;
  reg                 io_B_Valid_6_delay_3_1;
  reg                 io_B_Valid_6_delay_4;
  reg                 io_A_Valid_4_delay_1_6;
  reg                 io_A_Valid_4_delay_2_5;
  reg                 io_A_Valid_4_delay_3_4;
  reg                 io_A_Valid_4_delay_4_3;
  reg                 io_A_Valid_4_delay_5_2;
  reg                 io_A_Valid_4_delay_6_1;
  reg                 io_A_Valid_4_delay_7;
  reg                 io_B_Valid_7_delay_1_3;
  reg                 io_B_Valid_7_delay_2_2;
  reg                 io_B_Valid_7_delay_3_1;
  reg                 io_B_Valid_7_delay_4;
  reg        [15:0]   io_signCount_regNextWhen_5;
  reg                 io_B_Valid_0_delay_1_4;
  reg                 io_B_Valid_0_delay_2_3;
  reg                 io_B_Valid_0_delay_3_2;
  reg                 io_B_Valid_0_delay_4_1;
  reg                 io_B_Valid_0_delay_5;
  reg                 io_A_Valid_5_delay_1;
  reg                 io_B_Valid_1_delay_1_4;
  reg                 io_B_Valid_1_delay_2_3;
  reg                 io_B_Valid_1_delay_3_2;
  reg                 io_B_Valid_1_delay_4_1;
  reg                 io_B_Valid_1_delay_5;
  reg                 io_A_Valid_5_delay_1_1;
  reg                 io_A_Valid_5_delay_2;
  reg                 io_B_Valid_2_delay_1_4;
  reg                 io_B_Valid_2_delay_2_3;
  reg                 io_B_Valid_2_delay_3_2;
  reg                 io_B_Valid_2_delay_4_1;
  reg                 io_B_Valid_2_delay_5;
  reg                 io_A_Valid_5_delay_1_2;
  reg                 io_A_Valid_5_delay_2_1;
  reg                 io_A_Valid_5_delay_3;
  reg                 io_B_Valid_3_delay_1_4;
  reg                 io_B_Valid_3_delay_2_3;
  reg                 io_B_Valid_3_delay_3_2;
  reg                 io_B_Valid_3_delay_4_1;
  reg                 io_B_Valid_3_delay_5;
  reg                 io_A_Valid_5_delay_1_3;
  reg                 io_A_Valid_5_delay_2_2;
  reg                 io_A_Valid_5_delay_3_1;
  reg                 io_A_Valid_5_delay_4;
  reg                 io_B_Valid_4_delay_1_4;
  reg                 io_B_Valid_4_delay_2_3;
  reg                 io_B_Valid_4_delay_3_2;
  reg                 io_B_Valid_4_delay_4_1;
  reg                 io_B_Valid_4_delay_5;
  reg                 io_A_Valid_5_delay_1_4;
  reg                 io_A_Valid_5_delay_2_3;
  reg                 io_A_Valid_5_delay_3_2;
  reg                 io_A_Valid_5_delay_4_1;
  reg                 io_A_Valid_5_delay_5;
  reg                 io_B_Valid_5_delay_1_4;
  reg                 io_B_Valid_5_delay_2_3;
  reg                 io_B_Valid_5_delay_3_2;
  reg                 io_B_Valid_5_delay_4_1;
  reg                 io_B_Valid_5_delay_5;
  reg                 io_A_Valid_5_delay_1_5;
  reg                 io_A_Valid_5_delay_2_4;
  reg                 io_A_Valid_5_delay_3_3;
  reg                 io_A_Valid_5_delay_4_2;
  reg                 io_A_Valid_5_delay_5_1;
  reg                 io_A_Valid_5_delay_6;
  reg                 io_B_Valid_6_delay_1_4;
  reg                 io_B_Valid_6_delay_2_3;
  reg                 io_B_Valid_6_delay_3_2;
  reg                 io_B_Valid_6_delay_4_1;
  reg                 io_B_Valid_6_delay_5;
  reg                 io_A_Valid_5_delay_1_6;
  reg                 io_A_Valid_5_delay_2_5;
  reg                 io_A_Valid_5_delay_3_4;
  reg                 io_A_Valid_5_delay_4_3;
  reg                 io_A_Valid_5_delay_5_2;
  reg                 io_A_Valid_5_delay_6_1;
  reg                 io_A_Valid_5_delay_7;
  reg                 io_B_Valid_7_delay_1_4;
  reg                 io_B_Valid_7_delay_2_3;
  reg                 io_B_Valid_7_delay_3_2;
  reg                 io_B_Valid_7_delay_4_1;
  reg                 io_B_Valid_7_delay_5;
  reg        [15:0]   io_signCount_regNextWhen_6;
  reg                 io_B_Valid_0_delay_1_5;
  reg                 io_B_Valid_0_delay_2_4;
  reg                 io_B_Valid_0_delay_3_3;
  reg                 io_B_Valid_0_delay_4_2;
  reg                 io_B_Valid_0_delay_5_1;
  reg                 io_B_Valid_0_delay_6;
  reg                 io_A_Valid_6_delay_1;
  reg                 io_B_Valid_1_delay_1_5;
  reg                 io_B_Valid_1_delay_2_4;
  reg                 io_B_Valid_1_delay_3_3;
  reg                 io_B_Valid_1_delay_4_2;
  reg                 io_B_Valid_1_delay_5_1;
  reg                 io_B_Valid_1_delay_6;
  reg                 io_A_Valid_6_delay_1_1;
  reg                 io_A_Valid_6_delay_2;
  reg                 io_B_Valid_2_delay_1_5;
  reg                 io_B_Valid_2_delay_2_4;
  reg                 io_B_Valid_2_delay_3_3;
  reg                 io_B_Valid_2_delay_4_2;
  reg                 io_B_Valid_2_delay_5_1;
  reg                 io_B_Valid_2_delay_6;
  reg                 io_A_Valid_6_delay_1_2;
  reg                 io_A_Valid_6_delay_2_1;
  reg                 io_A_Valid_6_delay_3;
  reg                 io_B_Valid_3_delay_1_5;
  reg                 io_B_Valid_3_delay_2_4;
  reg                 io_B_Valid_3_delay_3_3;
  reg                 io_B_Valid_3_delay_4_2;
  reg                 io_B_Valid_3_delay_5_1;
  reg                 io_B_Valid_3_delay_6;
  reg                 io_A_Valid_6_delay_1_3;
  reg                 io_A_Valid_6_delay_2_2;
  reg                 io_A_Valid_6_delay_3_1;
  reg                 io_A_Valid_6_delay_4;
  reg                 io_B_Valid_4_delay_1_5;
  reg                 io_B_Valid_4_delay_2_4;
  reg                 io_B_Valid_4_delay_3_3;
  reg                 io_B_Valid_4_delay_4_2;
  reg                 io_B_Valid_4_delay_5_1;
  reg                 io_B_Valid_4_delay_6;
  reg                 io_A_Valid_6_delay_1_4;
  reg                 io_A_Valid_6_delay_2_3;
  reg                 io_A_Valid_6_delay_3_2;
  reg                 io_A_Valid_6_delay_4_1;
  reg                 io_A_Valid_6_delay_5;
  reg                 io_B_Valid_5_delay_1_5;
  reg                 io_B_Valid_5_delay_2_4;
  reg                 io_B_Valid_5_delay_3_3;
  reg                 io_B_Valid_5_delay_4_2;
  reg                 io_B_Valid_5_delay_5_1;
  reg                 io_B_Valid_5_delay_6;
  reg                 io_A_Valid_6_delay_1_5;
  reg                 io_A_Valid_6_delay_2_4;
  reg                 io_A_Valid_6_delay_3_3;
  reg                 io_A_Valid_6_delay_4_2;
  reg                 io_A_Valid_6_delay_5_1;
  reg                 io_A_Valid_6_delay_6;
  reg                 io_B_Valid_6_delay_1_5;
  reg                 io_B_Valid_6_delay_2_4;
  reg                 io_B_Valid_6_delay_3_3;
  reg                 io_B_Valid_6_delay_4_2;
  reg                 io_B_Valid_6_delay_5_1;
  reg                 io_B_Valid_6_delay_6;
  reg                 io_A_Valid_6_delay_1_6;
  reg                 io_A_Valid_6_delay_2_5;
  reg                 io_A_Valid_6_delay_3_4;
  reg                 io_A_Valid_6_delay_4_3;
  reg                 io_A_Valid_6_delay_5_2;
  reg                 io_A_Valid_6_delay_6_1;
  reg                 io_A_Valid_6_delay_7;
  reg                 io_B_Valid_7_delay_1_5;
  reg                 io_B_Valid_7_delay_2_4;
  reg                 io_B_Valid_7_delay_3_3;
  reg                 io_B_Valid_7_delay_4_2;
  reg                 io_B_Valid_7_delay_5_1;
  reg                 io_B_Valid_7_delay_6;
  reg        [15:0]   io_signCount_regNextWhen_7;
  reg                 io_B_Valid_0_delay_1_6;
  reg                 io_B_Valid_0_delay_2_5;
  reg                 io_B_Valid_0_delay_3_4;
  reg                 io_B_Valid_0_delay_4_3;
  reg                 io_B_Valid_0_delay_5_2;
  reg                 io_B_Valid_0_delay_6_1;
  reg                 io_B_Valid_0_delay_7;
  reg                 io_A_Valid_7_delay_1;
  reg                 io_B_Valid_1_delay_1_6;
  reg                 io_B_Valid_1_delay_2_5;
  reg                 io_B_Valid_1_delay_3_4;
  reg                 io_B_Valid_1_delay_4_3;
  reg                 io_B_Valid_1_delay_5_2;
  reg                 io_B_Valid_1_delay_6_1;
  reg                 io_B_Valid_1_delay_7;
  reg                 io_A_Valid_7_delay_1_1;
  reg                 io_A_Valid_7_delay_2;
  reg                 io_B_Valid_2_delay_1_6;
  reg                 io_B_Valid_2_delay_2_5;
  reg                 io_B_Valid_2_delay_3_4;
  reg                 io_B_Valid_2_delay_4_3;
  reg                 io_B_Valid_2_delay_5_2;
  reg                 io_B_Valid_2_delay_6_1;
  reg                 io_B_Valid_2_delay_7;
  reg                 io_A_Valid_7_delay_1_2;
  reg                 io_A_Valid_7_delay_2_1;
  reg                 io_A_Valid_7_delay_3;
  reg                 io_B_Valid_3_delay_1_6;
  reg                 io_B_Valid_3_delay_2_5;
  reg                 io_B_Valid_3_delay_3_4;
  reg                 io_B_Valid_3_delay_4_3;
  reg                 io_B_Valid_3_delay_5_2;
  reg                 io_B_Valid_3_delay_6_1;
  reg                 io_B_Valid_3_delay_7;
  reg                 io_A_Valid_7_delay_1_3;
  reg                 io_A_Valid_7_delay_2_2;
  reg                 io_A_Valid_7_delay_3_1;
  reg                 io_A_Valid_7_delay_4;
  reg                 io_B_Valid_4_delay_1_6;
  reg                 io_B_Valid_4_delay_2_5;
  reg                 io_B_Valid_4_delay_3_4;
  reg                 io_B_Valid_4_delay_4_3;
  reg                 io_B_Valid_4_delay_5_2;
  reg                 io_B_Valid_4_delay_6_1;
  reg                 io_B_Valid_4_delay_7;
  reg                 io_A_Valid_7_delay_1_4;
  reg                 io_A_Valid_7_delay_2_3;
  reg                 io_A_Valid_7_delay_3_2;
  reg                 io_A_Valid_7_delay_4_1;
  reg                 io_A_Valid_7_delay_5;
  reg                 io_B_Valid_5_delay_1_6;
  reg                 io_B_Valid_5_delay_2_5;
  reg                 io_B_Valid_5_delay_3_4;
  reg                 io_B_Valid_5_delay_4_3;
  reg                 io_B_Valid_5_delay_5_2;
  reg                 io_B_Valid_5_delay_6_1;
  reg                 io_B_Valid_5_delay_7;
  reg                 io_A_Valid_7_delay_1_5;
  reg                 io_A_Valid_7_delay_2_4;
  reg                 io_A_Valid_7_delay_3_3;
  reg                 io_A_Valid_7_delay_4_2;
  reg                 io_A_Valid_7_delay_5_1;
  reg                 io_A_Valid_7_delay_6;
  reg                 io_B_Valid_6_delay_1_6;
  reg                 io_B_Valid_6_delay_2_5;
  reg                 io_B_Valid_6_delay_3_4;
  reg                 io_B_Valid_6_delay_4_3;
  reg                 io_B_Valid_6_delay_5_2;
  reg                 io_B_Valid_6_delay_6_1;
  reg                 io_B_Valid_6_delay_7;
  reg                 io_A_Valid_7_delay_1_6;
  reg                 io_A_Valid_7_delay_2_5;
  reg                 io_A_Valid_7_delay_3_4;
  reg                 io_A_Valid_7_delay_4_3;
  reg                 io_A_Valid_7_delay_5_2;
  reg                 io_A_Valid_7_delay_6_1;
  reg                 io_A_Valid_7_delay_7;
  reg                 io_B_Valid_7_delay_1_6;
  reg                 io_B_Valid_7_delay_2_5;
  reg                 io_B_Valid_7_delay_3_4;
  reg                 io_B_Valid_7_delay_4_3;
  reg                 io_B_Valid_7_delay_5_2;
  reg                 io_B_Valid_7_delay_6_1;
  reg                 io_B_Valid_7_delay_7;

  PE_448 pE_512 (
    .activate  (io_MatrixA_0[7:0]             ), //i
    .weight    (io_MatrixB_0[7:0]             ), //i
    .valid     (pE_512_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_512_acount[7:0]            ), //o
    .bcount    (pE_512_bcount[7:0]            ), //o
    .PE_OUT    (pE_512_PE_OUT[31:0]           ), //o
    .finish    (pE_512_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_513 (
    .activate  (pE_512_acount[7:0]            ), //i
    .weight    (io_MatrixB_1[7:0]             ), //i
    .valid     (pE_513_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_513_acount[7:0]            ), //o
    .bcount    (pE_513_bcount[7:0]            ), //o
    .PE_OUT    (pE_513_PE_OUT[31:0]           ), //o
    .finish    (pE_513_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_514 (
    .activate  (pE_513_acount[7:0]            ), //i
    .weight    (io_MatrixB_2[7:0]             ), //i
    .valid     (pE_514_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_514_acount[7:0]            ), //o
    .bcount    (pE_514_bcount[7:0]            ), //o
    .PE_OUT    (pE_514_PE_OUT[31:0]           ), //o
    .finish    (pE_514_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_515 (
    .activate  (pE_514_acount[7:0]            ), //i
    .weight    (io_MatrixB_3[7:0]             ), //i
    .valid     (pE_515_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_515_acount[7:0]            ), //o
    .bcount    (pE_515_bcount[7:0]            ), //o
    .PE_OUT    (pE_515_PE_OUT[31:0]           ), //o
    .finish    (pE_515_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_516 (
    .activate  (pE_515_acount[7:0]            ), //i
    .weight    (io_MatrixB_4[7:0]             ), //i
    .valid     (pE_516_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_516_acount[7:0]            ), //o
    .bcount    (pE_516_bcount[7:0]            ), //o
    .PE_OUT    (pE_516_PE_OUT[31:0]           ), //o
    .finish    (pE_516_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_517 (
    .activate  (pE_516_acount[7:0]            ), //i
    .weight    (io_MatrixB_5[7:0]             ), //i
    .valid     (pE_517_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_517_acount[7:0]            ), //o
    .bcount    (pE_517_bcount[7:0]            ), //o
    .PE_OUT    (pE_517_PE_OUT[31:0]           ), //o
    .finish    (pE_517_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_518 (
    .activate  (pE_517_acount[7:0]            ), //i
    .weight    (io_MatrixB_6[7:0]             ), //i
    .valid     (pE_518_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_518_acount[7:0]            ), //o
    .bcount    (pE_518_bcount[7:0]            ), //o
    .PE_OUT    (pE_518_PE_OUT[31:0]           ), //o
    .finish    (pE_518_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_519 (
    .activate  (pE_518_acount[7:0]            ), //i
    .weight    (io_MatrixB_7[7:0]             ), //i
    .valid     (pE_519_valid                  ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (pE_519_acount[7:0]            ), //o
    .bcount    (pE_519_bcount[7:0]            ), //o
    .PE_OUT    (pE_519_PE_OUT[31:0]           ), //o
    .finish    (pE_519_finish                 ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE_448 pE_520 (
    .activate  (pE_520_acount[7:0]              ), //i
    .weight    (pE_512_bcount[7:0]              ), //i
    .valid     (pE_520_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_520_acount[7:0]              ), //o
    .bcount    (pE_520_bcount[7:0]              ), //o
    .PE_OUT    (pE_520_PE_OUT[31:0]             ), //o
    .finish    (pE_520_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_521 (
    .activate  (pE_512_acount[7:0]              ), //i
    .weight    (pE_512_bcount[7:0]              ), //i
    .valid     (pE_521_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_521_acount[7:0]              ), //o
    .bcount    (pE_521_bcount[7:0]              ), //o
    .PE_OUT    (pE_521_PE_OUT[31:0]             ), //o
    .finish    (pE_521_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_522 (
    .activate  (pE_513_acount[7:0]              ), //i
    .weight    (pE_513_bcount[7:0]              ), //i
    .valid     (pE_522_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_522_acount[7:0]              ), //o
    .bcount    (pE_522_bcount[7:0]              ), //o
    .PE_OUT    (pE_522_PE_OUT[31:0]             ), //o
    .finish    (pE_522_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_523 (
    .activate  (pE_514_acount[7:0]              ), //i
    .weight    (pE_514_bcount[7:0]              ), //i
    .valid     (pE_523_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_523_acount[7:0]              ), //o
    .bcount    (pE_523_bcount[7:0]              ), //o
    .PE_OUT    (pE_523_PE_OUT[31:0]             ), //o
    .finish    (pE_523_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_524 (
    .activate  (pE_515_acount[7:0]              ), //i
    .weight    (pE_515_bcount[7:0]              ), //i
    .valid     (pE_524_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_524_acount[7:0]              ), //o
    .bcount    (pE_524_bcount[7:0]              ), //o
    .PE_OUT    (pE_524_PE_OUT[31:0]             ), //o
    .finish    (pE_524_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_525 (
    .activate  (pE_516_acount[7:0]              ), //i
    .weight    (pE_516_bcount[7:0]              ), //i
    .valid     (pE_525_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_525_acount[7:0]              ), //o
    .bcount    (pE_525_bcount[7:0]              ), //o
    .PE_OUT    (pE_525_PE_OUT[31:0]             ), //o
    .finish    (pE_525_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_526 (
    .activate  (pE_517_acount[7:0]              ), //i
    .weight    (pE_517_bcount[7:0]              ), //i
    .valid     (pE_526_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_526_acount[7:0]              ), //o
    .bcount    (pE_526_bcount[7:0]              ), //o
    .PE_OUT    (pE_526_PE_OUT[31:0]             ), //o
    .finish    (pE_526_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_527 (
    .activate  (pE_518_acount[7:0]              ), //i
    .weight    (pE_518_bcount[7:0]              ), //i
    .valid     (pE_527_valid                    ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (pE_527_acount[7:0]              ), //o
    .bcount    (pE_527_bcount[7:0]              ), //o
    .PE_OUT    (pE_527_PE_OUT[31:0]             ), //o
    .finish    (pE_527_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_528 (
    .activate  (pE_528_acount[7:0]              ), //i
    .weight    (pE_520_bcount[7:0]              ), //i
    .valid     (pE_528_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_528_acount[7:0]              ), //o
    .bcount    (pE_528_bcount[7:0]              ), //o
    .PE_OUT    (pE_528_PE_OUT[31:0]             ), //o
    .finish    (pE_528_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_529 (
    .activate  (pE_520_acount[7:0]              ), //i
    .weight    (pE_520_bcount[7:0]              ), //i
    .valid     (pE_529_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_529_acount[7:0]              ), //o
    .bcount    (pE_529_bcount[7:0]              ), //o
    .PE_OUT    (pE_529_PE_OUT[31:0]             ), //o
    .finish    (pE_529_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_530 (
    .activate  (pE_521_acount[7:0]              ), //i
    .weight    (pE_521_bcount[7:0]              ), //i
    .valid     (pE_530_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_530_acount[7:0]              ), //o
    .bcount    (pE_530_bcount[7:0]              ), //o
    .PE_OUT    (pE_530_PE_OUT[31:0]             ), //o
    .finish    (pE_530_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_531 (
    .activate  (pE_522_acount[7:0]              ), //i
    .weight    (pE_522_bcount[7:0]              ), //i
    .valid     (pE_531_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_531_acount[7:0]              ), //o
    .bcount    (pE_531_bcount[7:0]              ), //o
    .PE_OUT    (pE_531_PE_OUT[31:0]             ), //o
    .finish    (pE_531_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_532 (
    .activate  (pE_523_acount[7:0]              ), //i
    .weight    (pE_523_bcount[7:0]              ), //i
    .valid     (pE_532_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_532_acount[7:0]              ), //o
    .bcount    (pE_532_bcount[7:0]              ), //o
    .PE_OUT    (pE_532_PE_OUT[31:0]             ), //o
    .finish    (pE_532_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_533 (
    .activate  (pE_524_acount[7:0]              ), //i
    .weight    (pE_524_bcount[7:0]              ), //i
    .valid     (pE_533_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_533_acount[7:0]              ), //o
    .bcount    (pE_533_bcount[7:0]              ), //o
    .PE_OUT    (pE_533_PE_OUT[31:0]             ), //o
    .finish    (pE_533_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_534 (
    .activate  (pE_525_acount[7:0]              ), //i
    .weight    (pE_525_bcount[7:0]              ), //i
    .valid     (pE_534_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_534_acount[7:0]              ), //o
    .bcount    (pE_534_bcount[7:0]              ), //o
    .PE_OUT    (pE_534_PE_OUT[31:0]             ), //o
    .finish    (pE_534_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_535 (
    .activate  (pE_526_acount[7:0]              ), //i
    .weight    (pE_526_bcount[7:0]              ), //i
    .valid     (pE_535_valid                    ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (pE_535_acount[7:0]              ), //o
    .bcount    (pE_535_bcount[7:0]              ), //o
    .PE_OUT    (pE_535_PE_OUT[31:0]             ), //o
    .finish    (pE_535_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_536 (
    .activate  (pE_536_acount[7:0]              ), //i
    .weight    (pE_528_bcount[7:0]              ), //i
    .valid     (pE_536_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_536_acount[7:0]              ), //o
    .bcount    (pE_536_bcount[7:0]              ), //o
    .PE_OUT    (pE_536_PE_OUT[31:0]             ), //o
    .finish    (pE_536_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_537 (
    .activate  (pE_528_acount[7:0]              ), //i
    .weight    (pE_528_bcount[7:0]              ), //i
    .valid     (pE_537_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_537_acount[7:0]              ), //o
    .bcount    (pE_537_bcount[7:0]              ), //o
    .PE_OUT    (pE_537_PE_OUT[31:0]             ), //o
    .finish    (pE_537_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_538 (
    .activate  (pE_529_acount[7:0]              ), //i
    .weight    (pE_529_bcount[7:0]              ), //i
    .valid     (pE_538_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_538_acount[7:0]              ), //o
    .bcount    (pE_538_bcount[7:0]              ), //o
    .PE_OUT    (pE_538_PE_OUT[31:0]             ), //o
    .finish    (pE_538_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_539 (
    .activate  (pE_530_acount[7:0]              ), //i
    .weight    (pE_530_bcount[7:0]              ), //i
    .valid     (pE_539_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_539_acount[7:0]              ), //o
    .bcount    (pE_539_bcount[7:0]              ), //o
    .PE_OUT    (pE_539_PE_OUT[31:0]             ), //o
    .finish    (pE_539_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_540 (
    .activate  (pE_531_acount[7:0]              ), //i
    .weight    (pE_531_bcount[7:0]              ), //i
    .valid     (pE_540_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_540_acount[7:0]              ), //o
    .bcount    (pE_540_bcount[7:0]              ), //o
    .PE_OUT    (pE_540_PE_OUT[31:0]             ), //o
    .finish    (pE_540_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_541 (
    .activate  (pE_532_acount[7:0]              ), //i
    .weight    (pE_532_bcount[7:0]              ), //i
    .valid     (pE_541_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_541_acount[7:0]              ), //o
    .bcount    (pE_541_bcount[7:0]              ), //o
    .PE_OUT    (pE_541_PE_OUT[31:0]             ), //o
    .finish    (pE_541_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_542 (
    .activate  (pE_533_acount[7:0]              ), //i
    .weight    (pE_533_bcount[7:0]              ), //i
    .valid     (pE_542_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_542_acount[7:0]              ), //o
    .bcount    (pE_542_bcount[7:0]              ), //o
    .PE_OUT    (pE_542_PE_OUT[31:0]             ), //o
    .finish    (pE_542_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_543 (
    .activate  (pE_534_acount[7:0]              ), //i
    .weight    (pE_534_bcount[7:0]              ), //i
    .valid     (pE_543_valid                    ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (pE_543_acount[7:0]              ), //o
    .bcount    (pE_543_bcount[7:0]              ), //o
    .PE_OUT    (pE_543_PE_OUT[31:0]             ), //o
    .finish    (pE_543_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_544 (
    .activate  (pE_544_acount[7:0]              ), //i
    .weight    (pE_536_bcount[7:0]              ), //i
    .valid     (pE_544_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_544_acount[7:0]              ), //o
    .bcount    (pE_544_bcount[7:0]              ), //o
    .PE_OUT    (pE_544_PE_OUT[31:0]             ), //o
    .finish    (pE_544_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_545 (
    .activate  (pE_536_acount[7:0]              ), //i
    .weight    (pE_536_bcount[7:0]              ), //i
    .valid     (pE_545_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_545_acount[7:0]              ), //o
    .bcount    (pE_545_bcount[7:0]              ), //o
    .PE_OUT    (pE_545_PE_OUT[31:0]             ), //o
    .finish    (pE_545_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_546 (
    .activate  (pE_537_acount[7:0]              ), //i
    .weight    (pE_537_bcount[7:0]              ), //i
    .valid     (pE_546_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_546_acount[7:0]              ), //o
    .bcount    (pE_546_bcount[7:0]              ), //o
    .PE_OUT    (pE_546_PE_OUT[31:0]             ), //o
    .finish    (pE_546_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_547 (
    .activate  (pE_538_acount[7:0]              ), //i
    .weight    (pE_538_bcount[7:0]              ), //i
    .valid     (pE_547_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_547_acount[7:0]              ), //o
    .bcount    (pE_547_bcount[7:0]              ), //o
    .PE_OUT    (pE_547_PE_OUT[31:0]             ), //o
    .finish    (pE_547_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_548 (
    .activate  (pE_539_acount[7:0]              ), //i
    .weight    (pE_539_bcount[7:0]              ), //i
    .valid     (pE_548_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_548_acount[7:0]              ), //o
    .bcount    (pE_548_bcount[7:0]              ), //o
    .PE_OUT    (pE_548_PE_OUT[31:0]             ), //o
    .finish    (pE_548_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_549 (
    .activate  (pE_540_acount[7:0]              ), //i
    .weight    (pE_540_bcount[7:0]              ), //i
    .valid     (pE_549_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_549_acount[7:0]              ), //o
    .bcount    (pE_549_bcount[7:0]              ), //o
    .PE_OUT    (pE_549_PE_OUT[31:0]             ), //o
    .finish    (pE_549_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_550 (
    .activate  (pE_541_acount[7:0]              ), //i
    .weight    (pE_541_bcount[7:0]              ), //i
    .valid     (pE_550_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_550_acount[7:0]              ), //o
    .bcount    (pE_550_bcount[7:0]              ), //o
    .PE_OUT    (pE_550_PE_OUT[31:0]             ), //o
    .finish    (pE_550_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_551 (
    .activate  (pE_542_acount[7:0]              ), //i
    .weight    (pE_542_bcount[7:0]              ), //i
    .valid     (pE_551_valid                    ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (pE_551_acount[7:0]              ), //o
    .bcount    (pE_551_bcount[7:0]              ), //o
    .PE_OUT    (pE_551_PE_OUT[31:0]             ), //o
    .finish    (pE_551_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_552 (
    .activate  (pE_552_acount[7:0]              ), //i
    .weight    (pE_544_bcount[7:0]              ), //i
    .valid     (pE_552_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_552_acount[7:0]              ), //o
    .bcount    (pE_552_bcount[7:0]              ), //o
    .PE_OUT    (pE_552_PE_OUT[31:0]             ), //o
    .finish    (pE_552_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_553 (
    .activate  (pE_544_acount[7:0]              ), //i
    .weight    (pE_544_bcount[7:0]              ), //i
    .valid     (pE_553_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_553_acount[7:0]              ), //o
    .bcount    (pE_553_bcount[7:0]              ), //o
    .PE_OUT    (pE_553_PE_OUT[31:0]             ), //o
    .finish    (pE_553_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_554 (
    .activate  (pE_545_acount[7:0]              ), //i
    .weight    (pE_545_bcount[7:0]              ), //i
    .valid     (pE_554_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_554_acount[7:0]              ), //o
    .bcount    (pE_554_bcount[7:0]              ), //o
    .PE_OUT    (pE_554_PE_OUT[31:0]             ), //o
    .finish    (pE_554_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_555 (
    .activate  (pE_546_acount[7:0]              ), //i
    .weight    (pE_546_bcount[7:0]              ), //i
    .valid     (pE_555_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_555_acount[7:0]              ), //o
    .bcount    (pE_555_bcount[7:0]              ), //o
    .PE_OUT    (pE_555_PE_OUT[31:0]             ), //o
    .finish    (pE_555_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_556 (
    .activate  (pE_547_acount[7:0]              ), //i
    .weight    (pE_547_bcount[7:0]              ), //i
    .valid     (pE_556_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_556_acount[7:0]              ), //o
    .bcount    (pE_556_bcount[7:0]              ), //o
    .PE_OUT    (pE_556_PE_OUT[31:0]             ), //o
    .finish    (pE_556_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_557 (
    .activate  (pE_548_acount[7:0]              ), //i
    .weight    (pE_548_bcount[7:0]              ), //i
    .valid     (pE_557_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_557_acount[7:0]              ), //o
    .bcount    (pE_557_bcount[7:0]              ), //o
    .PE_OUT    (pE_557_PE_OUT[31:0]             ), //o
    .finish    (pE_557_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_558 (
    .activate  (pE_549_acount[7:0]              ), //i
    .weight    (pE_549_bcount[7:0]              ), //i
    .valid     (pE_558_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_558_acount[7:0]              ), //o
    .bcount    (pE_558_bcount[7:0]              ), //o
    .PE_OUT    (pE_558_PE_OUT[31:0]             ), //o
    .finish    (pE_558_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_559 (
    .activate  (pE_550_acount[7:0]              ), //i
    .weight    (pE_550_bcount[7:0]              ), //i
    .valid     (pE_559_valid                    ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (pE_559_acount[7:0]              ), //o
    .bcount    (pE_559_bcount[7:0]              ), //o
    .PE_OUT    (pE_559_PE_OUT[31:0]             ), //o
    .finish    (pE_559_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_560 (
    .activate  (pE_560_acount[7:0]              ), //i
    .weight    (pE_552_bcount[7:0]              ), //i
    .valid     (pE_560_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_560_acount[7:0]              ), //o
    .bcount    (pE_560_bcount[7:0]              ), //o
    .PE_OUT    (pE_560_PE_OUT[31:0]             ), //o
    .finish    (pE_560_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_561 (
    .activate  (pE_552_acount[7:0]              ), //i
    .weight    (pE_552_bcount[7:0]              ), //i
    .valid     (pE_561_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_561_acount[7:0]              ), //o
    .bcount    (pE_561_bcount[7:0]              ), //o
    .PE_OUT    (pE_561_PE_OUT[31:0]             ), //o
    .finish    (pE_561_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_562 (
    .activate  (pE_553_acount[7:0]              ), //i
    .weight    (pE_553_bcount[7:0]              ), //i
    .valid     (pE_562_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_562_acount[7:0]              ), //o
    .bcount    (pE_562_bcount[7:0]              ), //o
    .PE_OUT    (pE_562_PE_OUT[31:0]             ), //o
    .finish    (pE_562_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_563 (
    .activate  (pE_554_acount[7:0]              ), //i
    .weight    (pE_554_bcount[7:0]              ), //i
    .valid     (pE_563_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_563_acount[7:0]              ), //o
    .bcount    (pE_563_bcount[7:0]              ), //o
    .PE_OUT    (pE_563_PE_OUT[31:0]             ), //o
    .finish    (pE_563_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_564 (
    .activate  (pE_555_acount[7:0]              ), //i
    .weight    (pE_555_bcount[7:0]              ), //i
    .valid     (pE_564_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_564_acount[7:0]              ), //o
    .bcount    (pE_564_bcount[7:0]              ), //o
    .PE_OUT    (pE_564_PE_OUT[31:0]             ), //o
    .finish    (pE_564_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_565 (
    .activate  (pE_556_acount[7:0]              ), //i
    .weight    (pE_556_bcount[7:0]              ), //i
    .valid     (pE_565_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_565_acount[7:0]              ), //o
    .bcount    (pE_565_bcount[7:0]              ), //o
    .PE_OUT    (pE_565_PE_OUT[31:0]             ), //o
    .finish    (pE_565_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_566 (
    .activate  (pE_557_acount[7:0]              ), //i
    .weight    (pE_557_bcount[7:0]              ), //i
    .valid     (pE_566_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_566_acount[7:0]              ), //o
    .bcount    (pE_566_bcount[7:0]              ), //o
    .PE_OUT    (pE_566_PE_OUT[31:0]             ), //o
    .finish    (pE_566_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_567 (
    .activate  (pE_558_acount[7:0]              ), //i
    .weight    (pE_558_bcount[7:0]              ), //i
    .valid     (pE_567_valid                    ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (pE_567_acount[7:0]              ), //o
    .bcount    (pE_567_bcount[7:0]              ), //o
    .PE_OUT    (pE_567_PE_OUT[31:0]             ), //o
    .finish    (pE_567_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_568 (
    .activate  (pE_568_acount[7:0]              ), //i
    .weight    (pE_560_bcount[7:0]              ), //i
    .valid     (pE_568_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_568_acount[7:0]              ), //o
    .bcount    (pE_568_bcount[7:0]              ), //o
    .PE_OUT    (pE_568_PE_OUT[31:0]             ), //o
    .finish    (pE_568_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_569 (
    .activate  (pE_560_acount[7:0]              ), //i
    .weight    (pE_560_bcount[7:0]              ), //i
    .valid     (pE_569_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_569_acount[7:0]              ), //o
    .bcount    (pE_569_bcount[7:0]              ), //o
    .PE_OUT    (pE_569_PE_OUT[31:0]             ), //o
    .finish    (pE_569_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_570 (
    .activate  (pE_561_acount[7:0]              ), //i
    .weight    (pE_561_bcount[7:0]              ), //i
    .valid     (pE_570_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_570_acount[7:0]              ), //o
    .bcount    (pE_570_bcount[7:0]              ), //o
    .PE_OUT    (pE_570_PE_OUT[31:0]             ), //o
    .finish    (pE_570_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_571 (
    .activate  (pE_562_acount[7:0]              ), //i
    .weight    (pE_562_bcount[7:0]              ), //i
    .valid     (pE_571_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_571_acount[7:0]              ), //o
    .bcount    (pE_571_bcount[7:0]              ), //o
    .PE_OUT    (pE_571_PE_OUT[31:0]             ), //o
    .finish    (pE_571_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_572 (
    .activate  (pE_563_acount[7:0]              ), //i
    .weight    (pE_563_bcount[7:0]              ), //i
    .valid     (pE_572_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_572_acount[7:0]              ), //o
    .bcount    (pE_572_bcount[7:0]              ), //o
    .PE_OUT    (pE_572_PE_OUT[31:0]             ), //o
    .finish    (pE_572_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_573 (
    .activate  (pE_564_acount[7:0]              ), //i
    .weight    (pE_564_bcount[7:0]              ), //i
    .valid     (pE_573_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_573_acount[7:0]              ), //o
    .bcount    (pE_573_bcount[7:0]              ), //o
    .PE_OUT    (pE_573_PE_OUT[31:0]             ), //o
    .finish    (pE_573_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_574 (
    .activate  (pE_565_acount[7:0]              ), //i
    .weight    (pE_565_bcount[7:0]              ), //i
    .valid     (pE_574_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_574_acount[7:0]              ), //o
    .bcount    (pE_574_bcount[7:0]              ), //o
    .PE_OUT    (pE_574_PE_OUT[31:0]             ), //o
    .finish    (pE_574_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE_448 pE_575 (
    .activate  (pE_566_acount[7:0]              ), //i
    .weight    (pE_566_bcount[7:0]              ), //i
    .valid     (pE_575_valid                    ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (pE_575_acount[7:0]              ), //o
    .bcount    (pE_575_bcount[7:0]              ), //o
    .PE_OUT    (pE_575_PE_OUT[31:0]             ), //o
    .finish    (pE_575_finish                   ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  always @(*) begin
    MatrixC_0 = 32'h0;
    if(when_SA_3D_l80) begin
      MatrixC_0 = pE_512_PE_OUT;
    end
    if(when_SA_3D_l80_1) begin
      MatrixC_0 = pE_513_PE_OUT;
    end
    if(when_SA_3D_l80_2) begin
      MatrixC_0 = pE_514_PE_OUT;
    end
    if(when_SA_3D_l80_3) begin
      MatrixC_0 = pE_515_PE_OUT;
    end
    if(when_SA_3D_l80_4) begin
      MatrixC_0 = pE_516_PE_OUT;
    end
    if(when_SA_3D_l80_5) begin
      MatrixC_0 = pE_517_PE_OUT;
    end
    if(when_SA_3D_l80_6) begin
      MatrixC_0 = pE_518_PE_OUT;
    end
    if(when_SA_3D_l80_7) begin
      MatrixC_0 = pE_519_PE_OUT;
    end
  end

  always @(*) begin
    tmp[0] = pE_512_valid;
    tmp[0] = pE_513_valid;
    tmp[0] = pE_514_valid;
    tmp[0] = pE_515_valid;
    tmp[0] = pE_516_valid;
    tmp[0] = pE_517_valid;
    tmp[0] = pE_518_valid;
    tmp[0] = pE_519_valid;
    tmp[1] = pE_520_valid;
    tmp[1] = pE_521_valid;
    tmp[1] = pE_522_valid;
    tmp[1] = pE_523_valid;
    tmp[1] = pE_524_valid;
    tmp[1] = pE_525_valid;
    tmp[1] = pE_526_valid;
    tmp[1] = pE_527_valid;
    tmp[2] = pE_528_valid;
    tmp[2] = pE_529_valid;
    tmp[2] = pE_530_valid;
    tmp[2] = pE_531_valid;
    tmp[2] = pE_532_valid;
    tmp[2] = pE_533_valid;
    tmp[2] = pE_534_valid;
    tmp[2] = pE_535_valid;
    tmp[3] = pE_536_valid;
    tmp[3] = pE_537_valid;
    tmp[3] = pE_538_valid;
    tmp[3] = pE_539_valid;
    tmp[3] = pE_540_valid;
    tmp[3] = pE_541_valid;
    tmp[3] = pE_542_valid;
    tmp[3] = pE_543_valid;
    tmp[4] = pE_544_valid;
    tmp[4] = pE_545_valid;
    tmp[4] = pE_546_valid;
    tmp[4] = pE_547_valid;
    tmp[4] = pE_548_valid;
    tmp[4] = pE_549_valid;
    tmp[4] = pE_550_valid;
    tmp[4] = pE_551_valid;
    tmp[5] = pE_552_valid;
    tmp[5] = pE_553_valid;
    tmp[5] = pE_554_valid;
    tmp[5] = pE_555_valid;
    tmp[5] = pE_556_valid;
    tmp[5] = pE_557_valid;
    tmp[5] = pE_558_valid;
    tmp[5] = pE_559_valid;
    tmp[6] = pE_560_valid;
    tmp[6] = pE_561_valid;
    tmp[6] = pE_562_valid;
    tmp[6] = pE_563_valid;
    tmp[6] = pE_564_valid;
    tmp[6] = pE_565_valid;
    tmp[6] = pE_566_valid;
    tmp[6] = pE_567_valid;
    tmp[7] = pE_568_valid;
    tmp[7] = pE_569_valid;
    tmp[7] = pE_570_valid;
    tmp[7] = pE_571_valid;
    tmp[7] = pE_572_valid;
    tmp[7] = pE_573_valid;
    tmp[7] = pE_574_valid;
    tmp[7] = pE_575_valid;
  end

  assign when_SA_3D_l80 = tmp[0];
  assign when_SA_3D_l80_1 = tmp[1];
  assign when_SA_3D_l80_2 = tmp[2];
  assign when_SA_3D_l80_3 = tmp[3];
  assign when_SA_3D_l80_4 = tmp[4];
  assign when_SA_3D_l80_5 = tmp[5];
  assign when_SA_3D_l80_6 = tmp[6];
  assign when_SA_3D_l80_7 = tmp[7];
  assign C_Valid_0 = (|tmp);
  always @(*) begin
    MatrixC_1 = 32'h0;
    if(when_SA_3D_l80_8) begin
      MatrixC_1 = pE_520_PE_OUT;
    end
    if(when_SA_3D_l80_9) begin
      MatrixC_1 = pE_521_PE_OUT;
    end
    if(when_SA_3D_l80_10) begin
      MatrixC_1 = pE_522_PE_OUT;
    end
    if(when_SA_3D_l80_11) begin
      MatrixC_1 = pE_523_PE_OUT;
    end
    if(when_SA_3D_l80_12) begin
      MatrixC_1 = pE_524_PE_OUT;
    end
    if(when_SA_3D_l80_13) begin
      MatrixC_1 = pE_525_PE_OUT;
    end
    if(when_SA_3D_l80_14) begin
      MatrixC_1 = pE_526_PE_OUT;
    end
    if(when_SA_3D_l80_15) begin
      MatrixC_1 = pE_527_PE_OUT;
    end
  end

  assign when_SA_3D_l80_8 = tmp[0];
  assign when_SA_3D_l80_9 = tmp[1];
  assign when_SA_3D_l80_10 = tmp[2];
  assign when_SA_3D_l80_11 = tmp[3];
  assign when_SA_3D_l80_12 = tmp[4];
  assign when_SA_3D_l80_13 = tmp[5];
  assign when_SA_3D_l80_14 = tmp[6];
  assign when_SA_3D_l80_15 = tmp[7];
  assign C_Valid_1 = (|tmp);
  always @(*) begin
    MatrixC_2 = 32'h0;
    if(when_SA_3D_l80_16) begin
      MatrixC_2 = pE_528_PE_OUT;
    end
    if(when_SA_3D_l80_17) begin
      MatrixC_2 = pE_529_PE_OUT;
    end
    if(when_SA_3D_l80_18) begin
      MatrixC_2 = pE_530_PE_OUT;
    end
    if(when_SA_3D_l80_19) begin
      MatrixC_2 = pE_531_PE_OUT;
    end
    if(when_SA_3D_l80_20) begin
      MatrixC_2 = pE_532_PE_OUT;
    end
    if(when_SA_3D_l80_21) begin
      MatrixC_2 = pE_533_PE_OUT;
    end
    if(when_SA_3D_l80_22) begin
      MatrixC_2 = pE_534_PE_OUT;
    end
    if(when_SA_3D_l80_23) begin
      MatrixC_2 = pE_535_PE_OUT;
    end
  end

  assign when_SA_3D_l80_16 = tmp[0];
  assign when_SA_3D_l80_17 = tmp[1];
  assign when_SA_3D_l80_18 = tmp[2];
  assign when_SA_3D_l80_19 = tmp[3];
  assign when_SA_3D_l80_20 = tmp[4];
  assign when_SA_3D_l80_21 = tmp[5];
  assign when_SA_3D_l80_22 = tmp[6];
  assign when_SA_3D_l80_23 = tmp[7];
  assign C_Valid_2 = (|tmp);
  always @(*) begin
    MatrixC_3 = 32'h0;
    if(when_SA_3D_l80_24) begin
      MatrixC_3 = pE_536_PE_OUT;
    end
    if(when_SA_3D_l80_25) begin
      MatrixC_3 = pE_537_PE_OUT;
    end
    if(when_SA_3D_l80_26) begin
      MatrixC_3 = pE_538_PE_OUT;
    end
    if(when_SA_3D_l80_27) begin
      MatrixC_3 = pE_539_PE_OUT;
    end
    if(when_SA_3D_l80_28) begin
      MatrixC_3 = pE_540_PE_OUT;
    end
    if(when_SA_3D_l80_29) begin
      MatrixC_3 = pE_541_PE_OUT;
    end
    if(when_SA_3D_l80_30) begin
      MatrixC_3 = pE_542_PE_OUT;
    end
    if(when_SA_3D_l80_31) begin
      MatrixC_3 = pE_543_PE_OUT;
    end
  end

  assign when_SA_3D_l80_24 = tmp[0];
  assign when_SA_3D_l80_25 = tmp[1];
  assign when_SA_3D_l80_26 = tmp[2];
  assign when_SA_3D_l80_27 = tmp[3];
  assign when_SA_3D_l80_28 = tmp[4];
  assign when_SA_3D_l80_29 = tmp[5];
  assign when_SA_3D_l80_30 = tmp[6];
  assign when_SA_3D_l80_31 = tmp[7];
  assign C_Valid_3 = (|tmp);
  always @(*) begin
    MatrixC_4 = 32'h0;
    if(when_SA_3D_l80_32) begin
      MatrixC_4 = pE_544_PE_OUT;
    end
    if(when_SA_3D_l80_33) begin
      MatrixC_4 = pE_545_PE_OUT;
    end
    if(when_SA_3D_l80_34) begin
      MatrixC_4 = pE_546_PE_OUT;
    end
    if(when_SA_3D_l80_35) begin
      MatrixC_4 = pE_547_PE_OUT;
    end
    if(when_SA_3D_l80_36) begin
      MatrixC_4 = pE_548_PE_OUT;
    end
    if(when_SA_3D_l80_37) begin
      MatrixC_4 = pE_549_PE_OUT;
    end
    if(when_SA_3D_l80_38) begin
      MatrixC_4 = pE_550_PE_OUT;
    end
    if(when_SA_3D_l80_39) begin
      MatrixC_4 = pE_551_PE_OUT;
    end
  end

  assign when_SA_3D_l80_32 = tmp[0];
  assign when_SA_3D_l80_33 = tmp[1];
  assign when_SA_3D_l80_34 = tmp[2];
  assign when_SA_3D_l80_35 = tmp[3];
  assign when_SA_3D_l80_36 = tmp[4];
  assign when_SA_3D_l80_37 = tmp[5];
  assign when_SA_3D_l80_38 = tmp[6];
  assign when_SA_3D_l80_39 = tmp[7];
  assign C_Valid_4 = (|tmp);
  always @(*) begin
    MatrixC_5 = 32'h0;
    if(when_SA_3D_l80_40) begin
      MatrixC_5 = pE_552_PE_OUT;
    end
    if(when_SA_3D_l80_41) begin
      MatrixC_5 = pE_553_PE_OUT;
    end
    if(when_SA_3D_l80_42) begin
      MatrixC_5 = pE_554_PE_OUT;
    end
    if(when_SA_3D_l80_43) begin
      MatrixC_5 = pE_555_PE_OUT;
    end
    if(when_SA_3D_l80_44) begin
      MatrixC_5 = pE_556_PE_OUT;
    end
    if(when_SA_3D_l80_45) begin
      MatrixC_5 = pE_557_PE_OUT;
    end
    if(when_SA_3D_l80_46) begin
      MatrixC_5 = pE_558_PE_OUT;
    end
    if(when_SA_3D_l80_47) begin
      MatrixC_5 = pE_559_PE_OUT;
    end
  end

  assign when_SA_3D_l80_40 = tmp[0];
  assign when_SA_3D_l80_41 = tmp[1];
  assign when_SA_3D_l80_42 = tmp[2];
  assign when_SA_3D_l80_43 = tmp[3];
  assign when_SA_3D_l80_44 = tmp[4];
  assign when_SA_3D_l80_45 = tmp[5];
  assign when_SA_3D_l80_46 = tmp[6];
  assign when_SA_3D_l80_47 = tmp[7];
  assign C_Valid_5 = (|tmp);
  always @(*) begin
    MatrixC_6 = 32'h0;
    if(when_SA_3D_l80_48) begin
      MatrixC_6 = pE_560_PE_OUT;
    end
    if(when_SA_3D_l80_49) begin
      MatrixC_6 = pE_561_PE_OUT;
    end
    if(when_SA_3D_l80_50) begin
      MatrixC_6 = pE_562_PE_OUT;
    end
    if(when_SA_3D_l80_51) begin
      MatrixC_6 = pE_563_PE_OUT;
    end
    if(when_SA_3D_l80_52) begin
      MatrixC_6 = pE_564_PE_OUT;
    end
    if(when_SA_3D_l80_53) begin
      MatrixC_6 = pE_565_PE_OUT;
    end
    if(when_SA_3D_l80_54) begin
      MatrixC_6 = pE_566_PE_OUT;
    end
    if(when_SA_3D_l80_55) begin
      MatrixC_6 = pE_567_PE_OUT;
    end
  end

  assign when_SA_3D_l80_48 = tmp[0];
  assign when_SA_3D_l80_49 = tmp[1];
  assign when_SA_3D_l80_50 = tmp[2];
  assign when_SA_3D_l80_51 = tmp[3];
  assign when_SA_3D_l80_52 = tmp[4];
  assign when_SA_3D_l80_53 = tmp[5];
  assign when_SA_3D_l80_54 = tmp[6];
  assign when_SA_3D_l80_55 = tmp[7];
  assign C_Valid_6 = (|tmp);
  always @(*) begin
    MatrixC_7 = 32'h0;
    if(when_SA_3D_l80_56) begin
      MatrixC_7 = pE_568_PE_OUT;
    end
    if(when_SA_3D_l80_57) begin
      MatrixC_7 = pE_569_PE_OUT;
    end
    if(when_SA_3D_l80_58) begin
      MatrixC_7 = pE_570_PE_OUT;
    end
    if(when_SA_3D_l80_59) begin
      MatrixC_7 = pE_571_PE_OUT;
    end
    if(when_SA_3D_l80_60) begin
      MatrixC_7 = pE_572_PE_OUT;
    end
    if(when_SA_3D_l80_61) begin
      MatrixC_7 = pE_573_PE_OUT;
    end
    if(when_SA_3D_l80_62) begin
      MatrixC_7 = pE_574_PE_OUT;
    end
    if(when_SA_3D_l80_63) begin
      MatrixC_7 = pE_575_PE_OUT;
    end
  end

  assign when_SA_3D_l80_56 = tmp[0];
  assign when_SA_3D_l80_57 = tmp[1];
  assign when_SA_3D_l80_58 = tmp[2];
  assign when_SA_3D_l80_59 = tmp[3];
  assign when_SA_3D_l80_60 = tmp[4];
  assign when_SA_3D_l80_61 = tmp[5];
  assign when_SA_3D_l80_62 = tmp[6];
  assign when_SA_3D_l80_63 = tmp[7];
  assign C_Valid_7 = (|tmp);
  assign pE_512_valid = (io_A_Valid_0 && io_B_Valid_0);
  assign pE_513_valid = (io_A_Valid_0_delay_1 && io_B_Valid_1);
  assign pE_514_valid = (io_A_Valid_0_delay_2 && io_B_Valid_2);
  assign pE_515_valid = (io_A_Valid_0_delay_3 && io_B_Valid_3);
  assign pE_516_valid = (io_A_Valid_0_delay_4 && io_B_Valid_4);
  assign pE_517_valid = (io_A_Valid_0_delay_5 && io_B_Valid_5);
  assign pE_518_valid = (io_A_Valid_0_delay_6 && io_B_Valid_6);
  assign pE_519_valid = (io_A_Valid_0_delay_7 && io_B_Valid_7);
  assign pE_520_valid = (io_A_Valid_1 && io_B_Valid_0_delay_1);
  assign pE_521_valid = (io_A_Valid_1_delay_1 && io_B_Valid_1_delay_1);
  assign pE_522_valid = (io_A_Valid_1_delay_2 && io_B_Valid_2_delay_1);
  assign pE_523_valid = (io_A_Valid_1_delay_3 && io_B_Valid_3_delay_1);
  assign pE_524_valid = (io_A_Valid_1_delay_4 && io_B_Valid_4_delay_1);
  assign pE_525_valid = (io_A_Valid_1_delay_5 && io_B_Valid_5_delay_1);
  assign pE_526_valid = (io_A_Valid_1_delay_6 && io_B_Valid_6_delay_1);
  assign pE_527_valid = (io_A_Valid_1_delay_7 && io_B_Valid_7_delay_1);
  assign pE_528_valid = (io_A_Valid_2 && io_B_Valid_0_delay_2);
  assign pE_529_valid = (io_A_Valid_2_delay_1 && io_B_Valid_1_delay_2);
  assign pE_530_valid = (io_A_Valid_2_delay_2 && io_B_Valid_2_delay_2);
  assign pE_531_valid = (io_A_Valid_2_delay_3 && io_B_Valid_3_delay_2);
  assign pE_532_valid = (io_A_Valid_2_delay_4 && io_B_Valid_4_delay_2);
  assign pE_533_valid = (io_A_Valid_2_delay_5 && io_B_Valid_5_delay_2);
  assign pE_534_valid = (io_A_Valid_2_delay_6 && io_B_Valid_6_delay_2);
  assign pE_535_valid = (io_A_Valid_2_delay_7 && io_B_Valid_7_delay_2);
  assign pE_536_valid = (io_A_Valid_3 && io_B_Valid_0_delay_3);
  assign pE_537_valid = (io_A_Valid_3_delay_1 && io_B_Valid_1_delay_3);
  assign pE_538_valid = (io_A_Valid_3_delay_2 && io_B_Valid_2_delay_3);
  assign pE_539_valid = (io_A_Valid_3_delay_3 && io_B_Valid_3_delay_3);
  assign pE_540_valid = (io_A_Valid_3_delay_4 && io_B_Valid_4_delay_3);
  assign pE_541_valid = (io_A_Valid_3_delay_5 && io_B_Valid_5_delay_3);
  assign pE_542_valid = (io_A_Valid_3_delay_6 && io_B_Valid_6_delay_3);
  assign pE_543_valid = (io_A_Valid_3_delay_7 && io_B_Valid_7_delay_3);
  assign pE_544_valid = (io_A_Valid_4 && io_B_Valid_0_delay_4);
  assign pE_545_valid = (io_A_Valid_4_delay_1 && io_B_Valid_1_delay_4);
  assign pE_546_valid = (io_A_Valid_4_delay_2 && io_B_Valid_2_delay_4);
  assign pE_547_valid = (io_A_Valid_4_delay_3 && io_B_Valid_3_delay_4);
  assign pE_548_valid = (io_A_Valid_4_delay_4 && io_B_Valid_4_delay_4);
  assign pE_549_valid = (io_A_Valid_4_delay_5 && io_B_Valid_5_delay_4);
  assign pE_550_valid = (io_A_Valid_4_delay_6 && io_B_Valid_6_delay_4);
  assign pE_551_valid = (io_A_Valid_4_delay_7 && io_B_Valid_7_delay_4);
  assign pE_552_valid = (io_A_Valid_5 && io_B_Valid_0_delay_5);
  assign pE_553_valid = (io_A_Valid_5_delay_1 && io_B_Valid_1_delay_5);
  assign pE_554_valid = (io_A_Valid_5_delay_2 && io_B_Valid_2_delay_5);
  assign pE_555_valid = (io_A_Valid_5_delay_3 && io_B_Valid_3_delay_5);
  assign pE_556_valid = (io_A_Valid_5_delay_4 && io_B_Valid_4_delay_5);
  assign pE_557_valid = (io_A_Valid_5_delay_5 && io_B_Valid_5_delay_5);
  assign pE_558_valid = (io_A_Valid_5_delay_6 && io_B_Valid_6_delay_5);
  assign pE_559_valid = (io_A_Valid_5_delay_7 && io_B_Valid_7_delay_5);
  assign pE_560_valid = (io_A_Valid_6 && io_B_Valid_0_delay_6);
  assign pE_561_valid = (io_A_Valid_6_delay_1 && io_B_Valid_1_delay_6);
  assign pE_562_valid = (io_A_Valid_6_delay_2 && io_B_Valid_2_delay_6);
  assign pE_563_valid = (io_A_Valid_6_delay_3 && io_B_Valid_3_delay_6);
  assign pE_564_valid = (io_A_Valid_6_delay_4 && io_B_Valid_4_delay_6);
  assign pE_565_valid = (io_A_Valid_6_delay_5 && io_B_Valid_5_delay_6);
  assign pE_566_valid = (io_A_Valid_6_delay_6 && io_B_Valid_6_delay_6);
  assign pE_567_valid = (io_A_Valid_6_delay_7 && io_B_Valid_7_delay_6);
  assign pE_568_valid = (io_A_Valid_7 && io_B_Valid_0_delay_7);
  assign pE_569_valid = (io_A_Valid_7_delay_1 && io_B_Valid_1_delay_7);
  assign pE_570_valid = (io_A_Valid_7_delay_2 && io_B_Valid_2_delay_7);
  assign pE_571_valid = (io_A_Valid_7_delay_3 && io_B_Valid_3_delay_7);
  assign pE_572_valid = (io_A_Valid_7_delay_4 && io_B_Valid_4_delay_7);
  assign pE_573_valid = (io_A_Valid_7_delay_5 && io_B_Valid_5_delay_7);
  assign pE_574_valid = (io_A_Valid_7_delay_6 && io_B_Valid_6_delay_7);
  assign pE_575_valid = (io_A_Valid_7_delay_7 && io_B_Valid_7_delay_7);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      io_signCount_regNextWhen <= 16'h0;
      io_signCount_regNextWhen_1 <= 16'h0;
      io_signCount_regNextWhen_2 <= 16'h0;
      io_signCount_regNextWhen_3 <= 16'h0;
      io_signCount_regNextWhen_4 <= 16'h0;
      io_signCount_regNextWhen_5 <= 16'h0;
      io_signCount_regNextWhen_6 <= 16'h0;
      io_signCount_regNextWhen_7 <= 16'h0;
    end else begin
      if(start) begin
        io_signCount_regNextWhen <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_1 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_2 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_3 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_4 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_5 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_6 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_7 <= io_signCount;
      end
    end
  end

  always @(posedge clk) begin
    io_A_Valid_0_delay_1 <= io_A_Valid_0;
    io_A_Valid_0_delay_1_1 <= io_A_Valid_0;
    io_A_Valid_0_delay_2 <= io_A_Valid_0_delay_1_1;
    io_A_Valid_0_delay_1_2 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_1 <= io_A_Valid_0_delay_1_2;
    io_A_Valid_0_delay_3 <= io_A_Valid_0_delay_2_1;
    io_A_Valid_0_delay_1_3 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_2 <= io_A_Valid_0_delay_1_3;
    io_A_Valid_0_delay_3_1 <= io_A_Valid_0_delay_2_2;
    io_A_Valid_0_delay_4 <= io_A_Valid_0_delay_3_1;
    io_A_Valid_0_delay_1_4 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_3 <= io_A_Valid_0_delay_1_4;
    io_A_Valid_0_delay_3_2 <= io_A_Valid_0_delay_2_3;
    io_A_Valid_0_delay_4_1 <= io_A_Valid_0_delay_3_2;
    io_A_Valid_0_delay_5 <= io_A_Valid_0_delay_4_1;
    io_A_Valid_0_delay_1_5 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_4 <= io_A_Valid_0_delay_1_5;
    io_A_Valid_0_delay_3_3 <= io_A_Valid_0_delay_2_4;
    io_A_Valid_0_delay_4_2 <= io_A_Valid_0_delay_3_3;
    io_A_Valid_0_delay_5_1 <= io_A_Valid_0_delay_4_2;
    io_A_Valid_0_delay_6 <= io_A_Valid_0_delay_5_1;
    io_A_Valid_0_delay_1_6 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_5 <= io_A_Valid_0_delay_1_6;
    io_A_Valid_0_delay_3_4 <= io_A_Valid_0_delay_2_5;
    io_A_Valid_0_delay_4_3 <= io_A_Valid_0_delay_3_4;
    io_A_Valid_0_delay_5_2 <= io_A_Valid_0_delay_4_3;
    io_A_Valid_0_delay_6_1 <= io_A_Valid_0_delay_5_2;
    io_A_Valid_0_delay_7 <= io_A_Valid_0_delay_6_1;
    io_B_Valid_0_delay_1 <= io_B_Valid_0;
    io_A_Valid_1_delay_1 <= io_A_Valid_1;
    io_B_Valid_1_delay_1 <= io_B_Valid_1;
    io_A_Valid_1_delay_1_1 <= io_A_Valid_1;
    io_A_Valid_1_delay_2 <= io_A_Valid_1_delay_1_1;
    io_B_Valid_2_delay_1 <= io_B_Valid_2;
    io_A_Valid_1_delay_1_2 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_1 <= io_A_Valid_1_delay_1_2;
    io_A_Valid_1_delay_3 <= io_A_Valid_1_delay_2_1;
    io_B_Valid_3_delay_1 <= io_B_Valid_3;
    io_A_Valid_1_delay_1_3 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_2 <= io_A_Valid_1_delay_1_3;
    io_A_Valid_1_delay_3_1 <= io_A_Valid_1_delay_2_2;
    io_A_Valid_1_delay_4 <= io_A_Valid_1_delay_3_1;
    io_B_Valid_4_delay_1 <= io_B_Valid_4;
    io_A_Valid_1_delay_1_4 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_3 <= io_A_Valid_1_delay_1_4;
    io_A_Valid_1_delay_3_2 <= io_A_Valid_1_delay_2_3;
    io_A_Valid_1_delay_4_1 <= io_A_Valid_1_delay_3_2;
    io_A_Valid_1_delay_5 <= io_A_Valid_1_delay_4_1;
    io_B_Valid_5_delay_1 <= io_B_Valid_5;
    io_A_Valid_1_delay_1_5 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_4 <= io_A_Valid_1_delay_1_5;
    io_A_Valid_1_delay_3_3 <= io_A_Valid_1_delay_2_4;
    io_A_Valid_1_delay_4_2 <= io_A_Valid_1_delay_3_3;
    io_A_Valid_1_delay_5_1 <= io_A_Valid_1_delay_4_2;
    io_A_Valid_1_delay_6 <= io_A_Valid_1_delay_5_1;
    io_B_Valid_6_delay_1 <= io_B_Valid_6;
    io_A_Valid_1_delay_1_6 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_5 <= io_A_Valid_1_delay_1_6;
    io_A_Valid_1_delay_3_4 <= io_A_Valid_1_delay_2_5;
    io_A_Valid_1_delay_4_3 <= io_A_Valid_1_delay_3_4;
    io_A_Valid_1_delay_5_2 <= io_A_Valid_1_delay_4_3;
    io_A_Valid_1_delay_6_1 <= io_A_Valid_1_delay_5_2;
    io_A_Valid_1_delay_7 <= io_A_Valid_1_delay_6_1;
    io_B_Valid_7_delay_1 <= io_B_Valid_7;
    io_B_Valid_0_delay_1_1 <= io_B_Valid_0;
    io_B_Valid_0_delay_2 <= io_B_Valid_0_delay_1_1;
    io_A_Valid_2_delay_1 <= io_A_Valid_2;
    io_B_Valid_1_delay_1_1 <= io_B_Valid_1;
    io_B_Valid_1_delay_2 <= io_B_Valid_1_delay_1_1;
    io_A_Valid_2_delay_1_1 <= io_A_Valid_2;
    io_A_Valid_2_delay_2 <= io_A_Valid_2_delay_1_1;
    io_B_Valid_2_delay_1_1 <= io_B_Valid_2;
    io_B_Valid_2_delay_2 <= io_B_Valid_2_delay_1_1;
    io_A_Valid_2_delay_1_2 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_1 <= io_A_Valid_2_delay_1_2;
    io_A_Valid_2_delay_3 <= io_A_Valid_2_delay_2_1;
    io_B_Valid_3_delay_1_1 <= io_B_Valid_3;
    io_B_Valid_3_delay_2 <= io_B_Valid_3_delay_1_1;
    io_A_Valid_2_delay_1_3 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_2 <= io_A_Valid_2_delay_1_3;
    io_A_Valid_2_delay_3_1 <= io_A_Valid_2_delay_2_2;
    io_A_Valid_2_delay_4 <= io_A_Valid_2_delay_3_1;
    io_B_Valid_4_delay_1_1 <= io_B_Valid_4;
    io_B_Valid_4_delay_2 <= io_B_Valid_4_delay_1_1;
    io_A_Valid_2_delay_1_4 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_3 <= io_A_Valid_2_delay_1_4;
    io_A_Valid_2_delay_3_2 <= io_A_Valid_2_delay_2_3;
    io_A_Valid_2_delay_4_1 <= io_A_Valid_2_delay_3_2;
    io_A_Valid_2_delay_5 <= io_A_Valid_2_delay_4_1;
    io_B_Valid_5_delay_1_1 <= io_B_Valid_5;
    io_B_Valid_5_delay_2 <= io_B_Valid_5_delay_1_1;
    io_A_Valid_2_delay_1_5 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_4 <= io_A_Valid_2_delay_1_5;
    io_A_Valid_2_delay_3_3 <= io_A_Valid_2_delay_2_4;
    io_A_Valid_2_delay_4_2 <= io_A_Valid_2_delay_3_3;
    io_A_Valid_2_delay_5_1 <= io_A_Valid_2_delay_4_2;
    io_A_Valid_2_delay_6 <= io_A_Valid_2_delay_5_1;
    io_B_Valid_6_delay_1_1 <= io_B_Valid_6;
    io_B_Valid_6_delay_2 <= io_B_Valid_6_delay_1_1;
    io_A_Valid_2_delay_1_6 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_5 <= io_A_Valid_2_delay_1_6;
    io_A_Valid_2_delay_3_4 <= io_A_Valid_2_delay_2_5;
    io_A_Valid_2_delay_4_3 <= io_A_Valid_2_delay_3_4;
    io_A_Valid_2_delay_5_2 <= io_A_Valid_2_delay_4_3;
    io_A_Valid_2_delay_6_1 <= io_A_Valid_2_delay_5_2;
    io_A_Valid_2_delay_7 <= io_A_Valid_2_delay_6_1;
    io_B_Valid_7_delay_1_1 <= io_B_Valid_7;
    io_B_Valid_7_delay_2 <= io_B_Valid_7_delay_1_1;
    io_B_Valid_0_delay_1_2 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_1 <= io_B_Valid_0_delay_1_2;
    io_B_Valid_0_delay_3 <= io_B_Valid_0_delay_2_1;
    io_A_Valid_3_delay_1 <= io_A_Valid_3;
    io_B_Valid_1_delay_1_2 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_1 <= io_B_Valid_1_delay_1_2;
    io_B_Valid_1_delay_3 <= io_B_Valid_1_delay_2_1;
    io_A_Valid_3_delay_1_1 <= io_A_Valid_3;
    io_A_Valid_3_delay_2 <= io_A_Valid_3_delay_1_1;
    io_B_Valid_2_delay_1_2 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_1 <= io_B_Valid_2_delay_1_2;
    io_B_Valid_2_delay_3 <= io_B_Valid_2_delay_2_1;
    io_A_Valid_3_delay_1_2 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_1 <= io_A_Valid_3_delay_1_2;
    io_A_Valid_3_delay_3 <= io_A_Valid_3_delay_2_1;
    io_B_Valid_3_delay_1_2 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_1 <= io_B_Valid_3_delay_1_2;
    io_B_Valid_3_delay_3 <= io_B_Valid_3_delay_2_1;
    io_A_Valid_3_delay_1_3 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_2 <= io_A_Valid_3_delay_1_3;
    io_A_Valid_3_delay_3_1 <= io_A_Valid_3_delay_2_2;
    io_A_Valid_3_delay_4 <= io_A_Valid_3_delay_3_1;
    io_B_Valid_4_delay_1_2 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_1 <= io_B_Valid_4_delay_1_2;
    io_B_Valid_4_delay_3 <= io_B_Valid_4_delay_2_1;
    io_A_Valid_3_delay_1_4 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_3 <= io_A_Valid_3_delay_1_4;
    io_A_Valid_3_delay_3_2 <= io_A_Valid_3_delay_2_3;
    io_A_Valid_3_delay_4_1 <= io_A_Valid_3_delay_3_2;
    io_A_Valid_3_delay_5 <= io_A_Valid_3_delay_4_1;
    io_B_Valid_5_delay_1_2 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_1 <= io_B_Valid_5_delay_1_2;
    io_B_Valid_5_delay_3 <= io_B_Valid_5_delay_2_1;
    io_A_Valid_3_delay_1_5 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_4 <= io_A_Valid_3_delay_1_5;
    io_A_Valid_3_delay_3_3 <= io_A_Valid_3_delay_2_4;
    io_A_Valid_3_delay_4_2 <= io_A_Valid_3_delay_3_3;
    io_A_Valid_3_delay_5_1 <= io_A_Valid_3_delay_4_2;
    io_A_Valid_3_delay_6 <= io_A_Valid_3_delay_5_1;
    io_B_Valid_6_delay_1_2 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_1 <= io_B_Valid_6_delay_1_2;
    io_B_Valid_6_delay_3 <= io_B_Valid_6_delay_2_1;
    io_A_Valid_3_delay_1_6 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_5 <= io_A_Valid_3_delay_1_6;
    io_A_Valid_3_delay_3_4 <= io_A_Valid_3_delay_2_5;
    io_A_Valid_3_delay_4_3 <= io_A_Valid_3_delay_3_4;
    io_A_Valid_3_delay_5_2 <= io_A_Valid_3_delay_4_3;
    io_A_Valid_3_delay_6_1 <= io_A_Valid_3_delay_5_2;
    io_A_Valid_3_delay_7 <= io_A_Valid_3_delay_6_1;
    io_B_Valid_7_delay_1_2 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_1 <= io_B_Valid_7_delay_1_2;
    io_B_Valid_7_delay_3 <= io_B_Valid_7_delay_2_1;
    io_B_Valid_0_delay_1_3 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_2 <= io_B_Valid_0_delay_1_3;
    io_B_Valid_0_delay_3_1 <= io_B_Valid_0_delay_2_2;
    io_B_Valid_0_delay_4 <= io_B_Valid_0_delay_3_1;
    io_A_Valid_4_delay_1 <= io_A_Valid_4;
    io_B_Valid_1_delay_1_3 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_2 <= io_B_Valid_1_delay_1_3;
    io_B_Valid_1_delay_3_1 <= io_B_Valid_1_delay_2_2;
    io_B_Valid_1_delay_4 <= io_B_Valid_1_delay_3_1;
    io_A_Valid_4_delay_1_1 <= io_A_Valid_4;
    io_A_Valid_4_delay_2 <= io_A_Valid_4_delay_1_1;
    io_B_Valid_2_delay_1_3 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_2 <= io_B_Valid_2_delay_1_3;
    io_B_Valid_2_delay_3_1 <= io_B_Valid_2_delay_2_2;
    io_B_Valid_2_delay_4 <= io_B_Valid_2_delay_3_1;
    io_A_Valid_4_delay_1_2 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_1 <= io_A_Valid_4_delay_1_2;
    io_A_Valid_4_delay_3 <= io_A_Valid_4_delay_2_1;
    io_B_Valid_3_delay_1_3 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_2 <= io_B_Valid_3_delay_1_3;
    io_B_Valid_3_delay_3_1 <= io_B_Valid_3_delay_2_2;
    io_B_Valid_3_delay_4 <= io_B_Valid_3_delay_3_1;
    io_A_Valid_4_delay_1_3 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_2 <= io_A_Valid_4_delay_1_3;
    io_A_Valid_4_delay_3_1 <= io_A_Valid_4_delay_2_2;
    io_A_Valid_4_delay_4 <= io_A_Valid_4_delay_3_1;
    io_B_Valid_4_delay_1_3 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_2 <= io_B_Valid_4_delay_1_3;
    io_B_Valid_4_delay_3_1 <= io_B_Valid_4_delay_2_2;
    io_B_Valid_4_delay_4 <= io_B_Valid_4_delay_3_1;
    io_A_Valid_4_delay_1_4 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_3 <= io_A_Valid_4_delay_1_4;
    io_A_Valid_4_delay_3_2 <= io_A_Valid_4_delay_2_3;
    io_A_Valid_4_delay_4_1 <= io_A_Valid_4_delay_3_2;
    io_A_Valid_4_delay_5 <= io_A_Valid_4_delay_4_1;
    io_B_Valid_5_delay_1_3 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_2 <= io_B_Valid_5_delay_1_3;
    io_B_Valid_5_delay_3_1 <= io_B_Valid_5_delay_2_2;
    io_B_Valid_5_delay_4 <= io_B_Valid_5_delay_3_1;
    io_A_Valid_4_delay_1_5 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_4 <= io_A_Valid_4_delay_1_5;
    io_A_Valid_4_delay_3_3 <= io_A_Valid_4_delay_2_4;
    io_A_Valid_4_delay_4_2 <= io_A_Valid_4_delay_3_3;
    io_A_Valid_4_delay_5_1 <= io_A_Valid_4_delay_4_2;
    io_A_Valid_4_delay_6 <= io_A_Valid_4_delay_5_1;
    io_B_Valid_6_delay_1_3 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_2 <= io_B_Valid_6_delay_1_3;
    io_B_Valid_6_delay_3_1 <= io_B_Valid_6_delay_2_2;
    io_B_Valid_6_delay_4 <= io_B_Valid_6_delay_3_1;
    io_A_Valid_4_delay_1_6 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_5 <= io_A_Valid_4_delay_1_6;
    io_A_Valid_4_delay_3_4 <= io_A_Valid_4_delay_2_5;
    io_A_Valid_4_delay_4_3 <= io_A_Valid_4_delay_3_4;
    io_A_Valid_4_delay_5_2 <= io_A_Valid_4_delay_4_3;
    io_A_Valid_4_delay_6_1 <= io_A_Valid_4_delay_5_2;
    io_A_Valid_4_delay_7 <= io_A_Valid_4_delay_6_1;
    io_B_Valid_7_delay_1_3 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_2 <= io_B_Valid_7_delay_1_3;
    io_B_Valid_7_delay_3_1 <= io_B_Valid_7_delay_2_2;
    io_B_Valid_7_delay_4 <= io_B_Valid_7_delay_3_1;
    io_B_Valid_0_delay_1_4 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_3 <= io_B_Valid_0_delay_1_4;
    io_B_Valid_0_delay_3_2 <= io_B_Valid_0_delay_2_3;
    io_B_Valid_0_delay_4_1 <= io_B_Valid_0_delay_3_2;
    io_B_Valid_0_delay_5 <= io_B_Valid_0_delay_4_1;
    io_A_Valid_5_delay_1 <= io_A_Valid_5;
    io_B_Valid_1_delay_1_4 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_3 <= io_B_Valid_1_delay_1_4;
    io_B_Valid_1_delay_3_2 <= io_B_Valid_1_delay_2_3;
    io_B_Valid_1_delay_4_1 <= io_B_Valid_1_delay_3_2;
    io_B_Valid_1_delay_5 <= io_B_Valid_1_delay_4_1;
    io_A_Valid_5_delay_1_1 <= io_A_Valid_5;
    io_A_Valid_5_delay_2 <= io_A_Valid_5_delay_1_1;
    io_B_Valid_2_delay_1_4 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_3 <= io_B_Valid_2_delay_1_4;
    io_B_Valid_2_delay_3_2 <= io_B_Valid_2_delay_2_3;
    io_B_Valid_2_delay_4_1 <= io_B_Valid_2_delay_3_2;
    io_B_Valid_2_delay_5 <= io_B_Valid_2_delay_4_1;
    io_A_Valid_5_delay_1_2 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_1 <= io_A_Valid_5_delay_1_2;
    io_A_Valid_5_delay_3 <= io_A_Valid_5_delay_2_1;
    io_B_Valid_3_delay_1_4 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_3 <= io_B_Valid_3_delay_1_4;
    io_B_Valid_3_delay_3_2 <= io_B_Valid_3_delay_2_3;
    io_B_Valid_3_delay_4_1 <= io_B_Valid_3_delay_3_2;
    io_B_Valid_3_delay_5 <= io_B_Valid_3_delay_4_1;
    io_A_Valid_5_delay_1_3 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_2 <= io_A_Valid_5_delay_1_3;
    io_A_Valid_5_delay_3_1 <= io_A_Valid_5_delay_2_2;
    io_A_Valid_5_delay_4 <= io_A_Valid_5_delay_3_1;
    io_B_Valid_4_delay_1_4 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_3 <= io_B_Valid_4_delay_1_4;
    io_B_Valid_4_delay_3_2 <= io_B_Valid_4_delay_2_3;
    io_B_Valid_4_delay_4_1 <= io_B_Valid_4_delay_3_2;
    io_B_Valid_4_delay_5 <= io_B_Valid_4_delay_4_1;
    io_A_Valid_5_delay_1_4 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_3 <= io_A_Valid_5_delay_1_4;
    io_A_Valid_5_delay_3_2 <= io_A_Valid_5_delay_2_3;
    io_A_Valid_5_delay_4_1 <= io_A_Valid_5_delay_3_2;
    io_A_Valid_5_delay_5 <= io_A_Valid_5_delay_4_1;
    io_B_Valid_5_delay_1_4 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_3 <= io_B_Valid_5_delay_1_4;
    io_B_Valid_5_delay_3_2 <= io_B_Valid_5_delay_2_3;
    io_B_Valid_5_delay_4_1 <= io_B_Valid_5_delay_3_2;
    io_B_Valid_5_delay_5 <= io_B_Valid_5_delay_4_1;
    io_A_Valid_5_delay_1_5 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_4 <= io_A_Valid_5_delay_1_5;
    io_A_Valid_5_delay_3_3 <= io_A_Valid_5_delay_2_4;
    io_A_Valid_5_delay_4_2 <= io_A_Valid_5_delay_3_3;
    io_A_Valid_5_delay_5_1 <= io_A_Valid_5_delay_4_2;
    io_A_Valid_5_delay_6 <= io_A_Valid_5_delay_5_1;
    io_B_Valid_6_delay_1_4 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_3 <= io_B_Valid_6_delay_1_4;
    io_B_Valid_6_delay_3_2 <= io_B_Valid_6_delay_2_3;
    io_B_Valid_6_delay_4_1 <= io_B_Valid_6_delay_3_2;
    io_B_Valid_6_delay_5 <= io_B_Valid_6_delay_4_1;
    io_A_Valid_5_delay_1_6 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_5 <= io_A_Valid_5_delay_1_6;
    io_A_Valid_5_delay_3_4 <= io_A_Valid_5_delay_2_5;
    io_A_Valid_5_delay_4_3 <= io_A_Valid_5_delay_3_4;
    io_A_Valid_5_delay_5_2 <= io_A_Valid_5_delay_4_3;
    io_A_Valid_5_delay_6_1 <= io_A_Valid_5_delay_5_2;
    io_A_Valid_5_delay_7 <= io_A_Valid_5_delay_6_1;
    io_B_Valid_7_delay_1_4 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_3 <= io_B_Valid_7_delay_1_4;
    io_B_Valid_7_delay_3_2 <= io_B_Valid_7_delay_2_3;
    io_B_Valid_7_delay_4_1 <= io_B_Valid_7_delay_3_2;
    io_B_Valid_7_delay_5 <= io_B_Valid_7_delay_4_1;
    io_B_Valid_0_delay_1_5 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_4 <= io_B_Valid_0_delay_1_5;
    io_B_Valid_0_delay_3_3 <= io_B_Valid_0_delay_2_4;
    io_B_Valid_0_delay_4_2 <= io_B_Valid_0_delay_3_3;
    io_B_Valid_0_delay_5_1 <= io_B_Valid_0_delay_4_2;
    io_B_Valid_0_delay_6 <= io_B_Valid_0_delay_5_1;
    io_A_Valid_6_delay_1 <= io_A_Valid_6;
    io_B_Valid_1_delay_1_5 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_4 <= io_B_Valid_1_delay_1_5;
    io_B_Valid_1_delay_3_3 <= io_B_Valid_1_delay_2_4;
    io_B_Valid_1_delay_4_2 <= io_B_Valid_1_delay_3_3;
    io_B_Valid_1_delay_5_1 <= io_B_Valid_1_delay_4_2;
    io_B_Valid_1_delay_6 <= io_B_Valid_1_delay_5_1;
    io_A_Valid_6_delay_1_1 <= io_A_Valid_6;
    io_A_Valid_6_delay_2 <= io_A_Valid_6_delay_1_1;
    io_B_Valid_2_delay_1_5 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_4 <= io_B_Valid_2_delay_1_5;
    io_B_Valid_2_delay_3_3 <= io_B_Valid_2_delay_2_4;
    io_B_Valid_2_delay_4_2 <= io_B_Valid_2_delay_3_3;
    io_B_Valid_2_delay_5_1 <= io_B_Valid_2_delay_4_2;
    io_B_Valid_2_delay_6 <= io_B_Valid_2_delay_5_1;
    io_A_Valid_6_delay_1_2 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_1 <= io_A_Valid_6_delay_1_2;
    io_A_Valid_6_delay_3 <= io_A_Valid_6_delay_2_1;
    io_B_Valid_3_delay_1_5 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_4 <= io_B_Valid_3_delay_1_5;
    io_B_Valid_3_delay_3_3 <= io_B_Valid_3_delay_2_4;
    io_B_Valid_3_delay_4_2 <= io_B_Valid_3_delay_3_3;
    io_B_Valid_3_delay_5_1 <= io_B_Valid_3_delay_4_2;
    io_B_Valid_3_delay_6 <= io_B_Valid_3_delay_5_1;
    io_A_Valid_6_delay_1_3 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_2 <= io_A_Valid_6_delay_1_3;
    io_A_Valid_6_delay_3_1 <= io_A_Valid_6_delay_2_2;
    io_A_Valid_6_delay_4 <= io_A_Valid_6_delay_3_1;
    io_B_Valid_4_delay_1_5 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_4 <= io_B_Valid_4_delay_1_5;
    io_B_Valid_4_delay_3_3 <= io_B_Valid_4_delay_2_4;
    io_B_Valid_4_delay_4_2 <= io_B_Valid_4_delay_3_3;
    io_B_Valid_4_delay_5_1 <= io_B_Valid_4_delay_4_2;
    io_B_Valid_4_delay_6 <= io_B_Valid_4_delay_5_1;
    io_A_Valid_6_delay_1_4 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_3 <= io_A_Valid_6_delay_1_4;
    io_A_Valid_6_delay_3_2 <= io_A_Valid_6_delay_2_3;
    io_A_Valid_6_delay_4_1 <= io_A_Valid_6_delay_3_2;
    io_A_Valid_6_delay_5 <= io_A_Valid_6_delay_4_1;
    io_B_Valid_5_delay_1_5 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_4 <= io_B_Valid_5_delay_1_5;
    io_B_Valid_5_delay_3_3 <= io_B_Valid_5_delay_2_4;
    io_B_Valid_5_delay_4_2 <= io_B_Valid_5_delay_3_3;
    io_B_Valid_5_delay_5_1 <= io_B_Valid_5_delay_4_2;
    io_B_Valid_5_delay_6 <= io_B_Valid_5_delay_5_1;
    io_A_Valid_6_delay_1_5 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_4 <= io_A_Valid_6_delay_1_5;
    io_A_Valid_6_delay_3_3 <= io_A_Valid_6_delay_2_4;
    io_A_Valid_6_delay_4_2 <= io_A_Valid_6_delay_3_3;
    io_A_Valid_6_delay_5_1 <= io_A_Valid_6_delay_4_2;
    io_A_Valid_6_delay_6 <= io_A_Valid_6_delay_5_1;
    io_B_Valid_6_delay_1_5 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_4 <= io_B_Valid_6_delay_1_5;
    io_B_Valid_6_delay_3_3 <= io_B_Valid_6_delay_2_4;
    io_B_Valid_6_delay_4_2 <= io_B_Valid_6_delay_3_3;
    io_B_Valid_6_delay_5_1 <= io_B_Valid_6_delay_4_2;
    io_B_Valid_6_delay_6 <= io_B_Valid_6_delay_5_1;
    io_A_Valid_6_delay_1_6 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_5 <= io_A_Valid_6_delay_1_6;
    io_A_Valid_6_delay_3_4 <= io_A_Valid_6_delay_2_5;
    io_A_Valid_6_delay_4_3 <= io_A_Valid_6_delay_3_4;
    io_A_Valid_6_delay_5_2 <= io_A_Valid_6_delay_4_3;
    io_A_Valid_6_delay_6_1 <= io_A_Valid_6_delay_5_2;
    io_A_Valid_6_delay_7 <= io_A_Valid_6_delay_6_1;
    io_B_Valid_7_delay_1_5 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_4 <= io_B_Valid_7_delay_1_5;
    io_B_Valid_7_delay_3_3 <= io_B_Valid_7_delay_2_4;
    io_B_Valid_7_delay_4_2 <= io_B_Valid_7_delay_3_3;
    io_B_Valid_7_delay_5_1 <= io_B_Valid_7_delay_4_2;
    io_B_Valid_7_delay_6 <= io_B_Valid_7_delay_5_1;
    io_B_Valid_0_delay_1_6 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_5 <= io_B_Valid_0_delay_1_6;
    io_B_Valid_0_delay_3_4 <= io_B_Valid_0_delay_2_5;
    io_B_Valid_0_delay_4_3 <= io_B_Valid_0_delay_3_4;
    io_B_Valid_0_delay_5_2 <= io_B_Valid_0_delay_4_3;
    io_B_Valid_0_delay_6_1 <= io_B_Valid_0_delay_5_2;
    io_B_Valid_0_delay_7 <= io_B_Valid_0_delay_6_1;
    io_A_Valid_7_delay_1 <= io_A_Valid_7;
    io_B_Valid_1_delay_1_6 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_5 <= io_B_Valid_1_delay_1_6;
    io_B_Valid_1_delay_3_4 <= io_B_Valid_1_delay_2_5;
    io_B_Valid_1_delay_4_3 <= io_B_Valid_1_delay_3_4;
    io_B_Valid_1_delay_5_2 <= io_B_Valid_1_delay_4_3;
    io_B_Valid_1_delay_6_1 <= io_B_Valid_1_delay_5_2;
    io_B_Valid_1_delay_7 <= io_B_Valid_1_delay_6_1;
    io_A_Valid_7_delay_1_1 <= io_A_Valid_7;
    io_A_Valid_7_delay_2 <= io_A_Valid_7_delay_1_1;
    io_B_Valid_2_delay_1_6 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_5 <= io_B_Valid_2_delay_1_6;
    io_B_Valid_2_delay_3_4 <= io_B_Valid_2_delay_2_5;
    io_B_Valid_2_delay_4_3 <= io_B_Valid_2_delay_3_4;
    io_B_Valid_2_delay_5_2 <= io_B_Valid_2_delay_4_3;
    io_B_Valid_2_delay_6_1 <= io_B_Valid_2_delay_5_2;
    io_B_Valid_2_delay_7 <= io_B_Valid_2_delay_6_1;
    io_A_Valid_7_delay_1_2 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_1 <= io_A_Valid_7_delay_1_2;
    io_A_Valid_7_delay_3 <= io_A_Valid_7_delay_2_1;
    io_B_Valid_3_delay_1_6 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_5 <= io_B_Valid_3_delay_1_6;
    io_B_Valid_3_delay_3_4 <= io_B_Valid_3_delay_2_5;
    io_B_Valid_3_delay_4_3 <= io_B_Valid_3_delay_3_4;
    io_B_Valid_3_delay_5_2 <= io_B_Valid_3_delay_4_3;
    io_B_Valid_3_delay_6_1 <= io_B_Valid_3_delay_5_2;
    io_B_Valid_3_delay_7 <= io_B_Valid_3_delay_6_1;
    io_A_Valid_7_delay_1_3 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_2 <= io_A_Valid_7_delay_1_3;
    io_A_Valid_7_delay_3_1 <= io_A_Valid_7_delay_2_2;
    io_A_Valid_7_delay_4 <= io_A_Valid_7_delay_3_1;
    io_B_Valid_4_delay_1_6 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_5 <= io_B_Valid_4_delay_1_6;
    io_B_Valid_4_delay_3_4 <= io_B_Valid_4_delay_2_5;
    io_B_Valid_4_delay_4_3 <= io_B_Valid_4_delay_3_4;
    io_B_Valid_4_delay_5_2 <= io_B_Valid_4_delay_4_3;
    io_B_Valid_4_delay_6_1 <= io_B_Valid_4_delay_5_2;
    io_B_Valid_4_delay_7 <= io_B_Valid_4_delay_6_1;
    io_A_Valid_7_delay_1_4 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_3 <= io_A_Valid_7_delay_1_4;
    io_A_Valid_7_delay_3_2 <= io_A_Valid_7_delay_2_3;
    io_A_Valid_7_delay_4_1 <= io_A_Valid_7_delay_3_2;
    io_A_Valid_7_delay_5 <= io_A_Valid_7_delay_4_1;
    io_B_Valid_5_delay_1_6 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_5 <= io_B_Valid_5_delay_1_6;
    io_B_Valid_5_delay_3_4 <= io_B_Valid_5_delay_2_5;
    io_B_Valid_5_delay_4_3 <= io_B_Valid_5_delay_3_4;
    io_B_Valid_5_delay_5_2 <= io_B_Valid_5_delay_4_3;
    io_B_Valid_5_delay_6_1 <= io_B_Valid_5_delay_5_2;
    io_B_Valid_5_delay_7 <= io_B_Valid_5_delay_6_1;
    io_A_Valid_7_delay_1_5 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_4 <= io_A_Valid_7_delay_1_5;
    io_A_Valid_7_delay_3_3 <= io_A_Valid_7_delay_2_4;
    io_A_Valid_7_delay_4_2 <= io_A_Valid_7_delay_3_3;
    io_A_Valid_7_delay_5_1 <= io_A_Valid_7_delay_4_2;
    io_A_Valid_7_delay_6 <= io_A_Valid_7_delay_5_1;
    io_B_Valid_6_delay_1_6 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_5 <= io_B_Valid_6_delay_1_6;
    io_B_Valid_6_delay_3_4 <= io_B_Valid_6_delay_2_5;
    io_B_Valid_6_delay_4_3 <= io_B_Valid_6_delay_3_4;
    io_B_Valid_6_delay_5_2 <= io_B_Valid_6_delay_4_3;
    io_B_Valid_6_delay_6_1 <= io_B_Valid_6_delay_5_2;
    io_B_Valid_6_delay_7 <= io_B_Valid_6_delay_6_1;
    io_A_Valid_7_delay_1_6 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_5 <= io_A_Valid_7_delay_1_6;
    io_A_Valid_7_delay_3_4 <= io_A_Valid_7_delay_2_5;
    io_A_Valid_7_delay_4_3 <= io_A_Valid_7_delay_3_4;
    io_A_Valid_7_delay_5_2 <= io_A_Valid_7_delay_4_3;
    io_A_Valid_7_delay_6_1 <= io_A_Valid_7_delay_5_2;
    io_A_Valid_7_delay_7 <= io_A_Valid_7_delay_6_1;
    io_B_Valid_7_delay_1_6 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_5 <= io_B_Valid_7_delay_1_6;
    io_B_Valid_7_delay_3_4 <= io_B_Valid_7_delay_2_5;
    io_B_Valid_7_delay_4_3 <= io_B_Valid_7_delay_3_4;
    io_B_Valid_7_delay_5_2 <= io_B_Valid_7_delay_4_3;
    io_B_Valid_7_delay_6_1 <= io_B_Valid_7_delay_5_2;
    io_B_Valid_7_delay_7 <= io_B_Valid_7_delay_6_1;
  end


endmodule

//PE_63 replaced by PE_448

//PE_62 replaced by PE_448

//PE_61 replaced by PE_448

//PE_60 replaced by PE_448

//PE_59 replaced by PE_448

//PE_58 replaced by PE_448

//PE_57 replaced by PE_448

//PE_56 replaced by PE_448

//PE_55 replaced by PE_448

//PE_54 replaced by PE_448

//PE_53 replaced by PE_448

//PE_52 replaced by PE_448

//PE_51 replaced by PE_448

//PE_50 replaced by PE_448

//PE_49 replaced by PE_448

//PE_48 replaced by PE_448

//PE_47 replaced by PE_448

//PE_46 replaced by PE_448

//PE_45 replaced by PE_448

//PE_44 replaced by PE_448

//PE_43 replaced by PE_448

//PE_42 replaced by PE_448

//PE_41 replaced by PE_448

//PE_40 replaced by PE_448

//PE_39 replaced by PE_448

//PE_38 replaced by PE_448

//PE_37 replaced by PE_448

//PE_36 replaced by PE_448

//PE_35 replaced by PE_448

//PE_34 replaced by PE_448

//PE_33 replaced by PE_448

//PE_32 replaced by PE_448

//PE_31 replaced by PE_448

//PE_30 replaced by PE_448

//PE_29 replaced by PE_448

//PE_28 replaced by PE_448

//PE_27 replaced by PE_448

//PE_26 replaced by PE_448

//PE_25 replaced by PE_448

//PE_24 replaced by PE_448

//PE_23 replaced by PE_448

//PE_22 replaced by PE_448

//PE_21 replaced by PE_448

//PE_20 replaced by PE_448

//PE_19 replaced by PE_448

//PE_18 replaced by PE_448

//PE_17 replaced by PE_448

//PE_16 replaced by PE_448

//PE_15 replaced by PE_448

//PE_14 replaced by PE_448

//PE_13 replaced by PE_448

//PE_12 replaced by PE_448

//PE_11 replaced by PE_448

//PE_10 replaced by PE_448

//PE_9 replaced by PE_448

//PE_8 replaced by PE_448

//PE_7 replaced by PE_448

//PE_6 replaced by PE_448

//PE_5 replaced by PE_448

//PE_4 replaced by PE_448

//PE_3 replaced by PE_448

//PE_2 replaced by PE_448

//PE_1 replaced by PE_448

//PE replaced by PE_448

//PE_127 replaced by PE_448

//PE_126 replaced by PE_448

//PE_125 replaced by PE_448

//PE_124 replaced by PE_448

//PE_123 replaced by PE_448

//PE_122 replaced by PE_448

//PE_121 replaced by PE_448

//PE_120 replaced by PE_448

//PE_119 replaced by PE_448

//PE_118 replaced by PE_448

//PE_117 replaced by PE_448

//PE_116 replaced by PE_448

//PE_115 replaced by PE_448

//PE_114 replaced by PE_448

//PE_113 replaced by PE_448

//PE_112 replaced by PE_448

//PE_111 replaced by PE_448

//PE_110 replaced by PE_448

//PE_109 replaced by PE_448

//PE_108 replaced by PE_448

//PE_107 replaced by PE_448

//PE_106 replaced by PE_448

//PE_105 replaced by PE_448

//PE_104 replaced by PE_448

//PE_103 replaced by PE_448

//PE_102 replaced by PE_448

//PE_101 replaced by PE_448

//PE_100 replaced by PE_448

//PE_99 replaced by PE_448

//PE_98 replaced by PE_448

//PE_97 replaced by PE_448

//PE_96 replaced by PE_448

//PE_95 replaced by PE_448

//PE_94 replaced by PE_448

//PE_93 replaced by PE_448

//PE_92 replaced by PE_448

//PE_91 replaced by PE_448

//PE_90 replaced by PE_448

//PE_89 replaced by PE_448

//PE_88 replaced by PE_448

//PE_87 replaced by PE_448

//PE_86 replaced by PE_448

//PE_85 replaced by PE_448

//PE_84 replaced by PE_448

//PE_83 replaced by PE_448

//PE_82 replaced by PE_448

//PE_81 replaced by PE_448

//PE_80 replaced by PE_448

//PE_79 replaced by PE_448

//PE_78 replaced by PE_448

//PE_77 replaced by PE_448

//PE_76 replaced by PE_448

//PE_75 replaced by PE_448

//PE_74 replaced by PE_448

//PE_73 replaced by PE_448

//PE_72 replaced by PE_448

//PE_71 replaced by PE_448

//PE_70 replaced by PE_448

//PE_69 replaced by PE_448

//PE_68 replaced by PE_448

//PE_67 replaced by PE_448

//PE_66 replaced by PE_448

//PE_65 replaced by PE_448

//PE_64 replaced by PE_448

//PE_191 replaced by PE_448

//PE_190 replaced by PE_448

//PE_189 replaced by PE_448

//PE_188 replaced by PE_448

//PE_187 replaced by PE_448

//PE_186 replaced by PE_448

//PE_185 replaced by PE_448

//PE_184 replaced by PE_448

//PE_183 replaced by PE_448

//PE_182 replaced by PE_448

//PE_181 replaced by PE_448

//PE_180 replaced by PE_448

//PE_179 replaced by PE_448

//PE_178 replaced by PE_448

//PE_177 replaced by PE_448

//PE_176 replaced by PE_448

//PE_175 replaced by PE_448

//PE_174 replaced by PE_448

//PE_173 replaced by PE_448

//PE_172 replaced by PE_448

//PE_171 replaced by PE_448

//PE_170 replaced by PE_448

//PE_169 replaced by PE_448

//PE_168 replaced by PE_448

//PE_167 replaced by PE_448

//PE_166 replaced by PE_448

//PE_165 replaced by PE_448

//PE_164 replaced by PE_448

//PE_163 replaced by PE_448

//PE_162 replaced by PE_448

//PE_161 replaced by PE_448

//PE_160 replaced by PE_448

//PE_159 replaced by PE_448

//PE_158 replaced by PE_448

//PE_157 replaced by PE_448

//PE_156 replaced by PE_448

//PE_155 replaced by PE_448

//PE_154 replaced by PE_448

//PE_153 replaced by PE_448

//PE_152 replaced by PE_448

//PE_151 replaced by PE_448

//PE_150 replaced by PE_448

//PE_149 replaced by PE_448

//PE_148 replaced by PE_448

//PE_147 replaced by PE_448

//PE_146 replaced by PE_448

//PE_145 replaced by PE_448

//PE_144 replaced by PE_448

//PE_143 replaced by PE_448

//PE_142 replaced by PE_448

//PE_141 replaced by PE_448

//PE_140 replaced by PE_448

//PE_139 replaced by PE_448

//PE_138 replaced by PE_448

//PE_137 replaced by PE_448

//PE_136 replaced by PE_448

//PE_135 replaced by PE_448

//PE_134 replaced by PE_448

//PE_133 replaced by PE_448

//PE_132 replaced by PE_448

//PE_131 replaced by PE_448

//PE_130 replaced by PE_448

//PE_129 replaced by PE_448

//PE_128 replaced by PE_448

//PE_255 replaced by PE_448

//PE_254 replaced by PE_448

//PE_253 replaced by PE_448

//PE_252 replaced by PE_448

//PE_251 replaced by PE_448

//PE_250 replaced by PE_448

//PE_249 replaced by PE_448

//PE_248 replaced by PE_448

//PE_247 replaced by PE_448

//PE_246 replaced by PE_448

//PE_245 replaced by PE_448

//PE_244 replaced by PE_448

//PE_243 replaced by PE_448

//PE_242 replaced by PE_448

//PE_241 replaced by PE_448

//PE_240 replaced by PE_448

//PE_239 replaced by PE_448

//PE_238 replaced by PE_448

//PE_237 replaced by PE_448

//PE_236 replaced by PE_448

//PE_235 replaced by PE_448

//PE_234 replaced by PE_448

//PE_233 replaced by PE_448

//PE_232 replaced by PE_448

//PE_231 replaced by PE_448

//PE_230 replaced by PE_448

//PE_229 replaced by PE_448

//PE_228 replaced by PE_448

//PE_227 replaced by PE_448

//PE_226 replaced by PE_448

//PE_225 replaced by PE_448

//PE_224 replaced by PE_448

//PE_223 replaced by PE_448

//PE_222 replaced by PE_448

//PE_221 replaced by PE_448

//PE_220 replaced by PE_448

//PE_219 replaced by PE_448

//PE_218 replaced by PE_448

//PE_217 replaced by PE_448

//PE_216 replaced by PE_448

//PE_215 replaced by PE_448

//PE_214 replaced by PE_448

//PE_213 replaced by PE_448

//PE_212 replaced by PE_448

//PE_211 replaced by PE_448

//PE_210 replaced by PE_448

//PE_209 replaced by PE_448

//PE_208 replaced by PE_448

//PE_207 replaced by PE_448

//PE_206 replaced by PE_448

//PE_205 replaced by PE_448

//PE_204 replaced by PE_448

//PE_203 replaced by PE_448

//PE_202 replaced by PE_448

//PE_201 replaced by PE_448

//PE_200 replaced by PE_448

//PE_199 replaced by PE_448

//PE_198 replaced by PE_448

//PE_197 replaced by PE_448

//PE_196 replaced by PE_448

//PE_195 replaced by PE_448

//PE_194 replaced by PE_448

//PE_193 replaced by PE_448

//PE_192 replaced by PE_448

//PE_319 replaced by PE_448

//PE_318 replaced by PE_448

//PE_317 replaced by PE_448

//PE_316 replaced by PE_448

//PE_315 replaced by PE_448

//PE_314 replaced by PE_448

//PE_313 replaced by PE_448

//PE_312 replaced by PE_448

//PE_311 replaced by PE_448

//PE_310 replaced by PE_448

//PE_309 replaced by PE_448

//PE_308 replaced by PE_448

//PE_307 replaced by PE_448

//PE_306 replaced by PE_448

//PE_305 replaced by PE_448

//PE_304 replaced by PE_448

//PE_303 replaced by PE_448

//PE_302 replaced by PE_448

//PE_301 replaced by PE_448

//PE_300 replaced by PE_448

//PE_299 replaced by PE_448

//PE_298 replaced by PE_448

//PE_297 replaced by PE_448

//PE_296 replaced by PE_448

//PE_295 replaced by PE_448

//PE_294 replaced by PE_448

//PE_293 replaced by PE_448

//PE_292 replaced by PE_448

//PE_291 replaced by PE_448

//PE_290 replaced by PE_448

//PE_289 replaced by PE_448

//PE_288 replaced by PE_448

//PE_287 replaced by PE_448

//PE_286 replaced by PE_448

//PE_285 replaced by PE_448

//PE_284 replaced by PE_448

//PE_283 replaced by PE_448

//PE_282 replaced by PE_448

//PE_281 replaced by PE_448

//PE_280 replaced by PE_448

//PE_279 replaced by PE_448

//PE_278 replaced by PE_448

//PE_277 replaced by PE_448

//PE_276 replaced by PE_448

//PE_275 replaced by PE_448

//PE_274 replaced by PE_448

//PE_273 replaced by PE_448

//PE_272 replaced by PE_448

//PE_271 replaced by PE_448

//PE_270 replaced by PE_448

//PE_269 replaced by PE_448

//PE_268 replaced by PE_448

//PE_267 replaced by PE_448

//PE_266 replaced by PE_448

//PE_265 replaced by PE_448

//PE_264 replaced by PE_448

//PE_263 replaced by PE_448

//PE_262 replaced by PE_448

//PE_261 replaced by PE_448

//PE_260 replaced by PE_448

//PE_259 replaced by PE_448

//PE_258 replaced by PE_448

//PE_257 replaced by PE_448

//PE_256 replaced by PE_448

//PE_383 replaced by PE_448

//PE_382 replaced by PE_448

//PE_381 replaced by PE_448

//PE_380 replaced by PE_448

//PE_379 replaced by PE_448

//PE_378 replaced by PE_448

//PE_377 replaced by PE_448

//PE_376 replaced by PE_448

//PE_375 replaced by PE_448

//PE_374 replaced by PE_448

//PE_373 replaced by PE_448

//PE_372 replaced by PE_448

//PE_371 replaced by PE_448

//PE_370 replaced by PE_448

//PE_369 replaced by PE_448

//PE_368 replaced by PE_448

//PE_367 replaced by PE_448

//PE_366 replaced by PE_448

//PE_365 replaced by PE_448

//PE_364 replaced by PE_448

//PE_363 replaced by PE_448

//PE_362 replaced by PE_448

//PE_361 replaced by PE_448

//PE_360 replaced by PE_448

//PE_359 replaced by PE_448

//PE_358 replaced by PE_448

//PE_357 replaced by PE_448

//PE_356 replaced by PE_448

//PE_355 replaced by PE_448

//PE_354 replaced by PE_448

//PE_353 replaced by PE_448

//PE_352 replaced by PE_448

//PE_351 replaced by PE_448

//PE_350 replaced by PE_448

//PE_349 replaced by PE_448

//PE_348 replaced by PE_448

//PE_347 replaced by PE_448

//PE_346 replaced by PE_448

//PE_345 replaced by PE_448

//PE_344 replaced by PE_448

//PE_343 replaced by PE_448

//PE_342 replaced by PE_448

//PE_341 replaced by PE_448

//PE_340 replaced by PE_448

//PE_339 replaced by PE_448

//PE_338 replaced by PE_448

//PE_337 replaced by PE_448

//PE_336 replaced by PE_448

//PE_335 replaced by PE_448

//PE_334 replaced by PE_448

//PE_333 replaced by PE_448

//PE_332 replaced by PE_448

//PE_331 replaced by PE_448

//PE_330 replaced by PE_448

//PE_329 replaced by PE_448

//PE_328 replaced by PE_448

//PE_327 replaced by PE_448

//PE_326 replaced by PE_448

//PE_325 replaced by PE_448

//PE_324 replaced by PE_448

//PE_323 replaced by PE_448

//PE_322 replaced by PE_448

//PE_321 replaced by PE_448

//PE_320 replaced by PE_448

//PE_447 replaced by PE_448

//PE_446 replaced by PE_448

//PE_445 replaced by PE_448

//PE_444 replaced by PE_448

//PE_443 replaced by PE_448

//PE_442 replaced by PE_448

//PE_441 replaced by PE_448

//PE_440 replaced by PE_448

//PE_439 replaced by PE_448

//PE_438 replaced by PE_448

//PE_437 replaced by PE_448

//PE_436 replaced by PE_448

//PE_435 replaced by PE_448

//PE_434 replaced by PE_448

//PE_433 replaced by PE_448

//PE_432 replaced by PE_448

//PE_431 replaced by PE_448

//PE_430 replaced by PE_448

//PE_429 replaced by PE_448

//PE_428 replaced by PE_448

//PE_427 replaced by PE_448

//PE_426 replaced by PE_448

//PE_425 replaced by PE_448

//PE_424 replaced by PE_448

//PE_423 replaced by PE_448

//PE_422 replaced by PE_448

//PE_421 replaced by PE_448

//PE_420 replaced by PE_448

//PE_419 replaced by PE_448

//PE_418 replaced by PE_448

//PE_417 replaced by PE_448

//PE_416 replaced by PE_448

//PE_415 replaced by PE_448

//PE_414 replaced by PE_448

//PE_413 replaced by PE_448

//PE_412 replaced by PE_448

//PE_411 replaced by PE_448

//PE_410 replaced by PE_448

//PE_409 replaced by PE_448

//PE_408 replaced by PE_448

//PE_407 replaced by PE_448

//PE_406 replaced by PE_448

//PE_405 replaced by PE_448

//PE_404 replaced by PE_448

//PE_403 replaced by PE_448

//PE_402 replaced by PE_448

//PE_401 replaced by PE_448

//PE_400 replaced by PE_448

//PE_399 replaced by PE_448

//PE_398 replaced by PE_448

//PE_397 replaced by PE_448

//PE_396 replaced by PE_448

//PE_395 replaced by PE_448

//PE_394 replaced by PE_448

//PE_393 replaced by PE_448

//PE_392 replaced by PE_448

//PE_391 replaced by PE_448

//PE_390 replaced by PE_448

//PE_389 replaced by PE_448

//PE_388 replaced by PE_448

//PE_387 replaced by PE_448

//PE_386 replaced by PE_448

//PE_385 replaced by PE_448

//PE_384 replaced by PE_448

//PE_511 replaced by PE_448

//PE_510 replaced by PE_448

//PE_509 replaced by PE_448

//PE_508 replaced by PE_448

//PE_507 replaced by PE_448

//PE_506 replaced by PE_448

//PE_505 replaced by PE_448

//PE_504 replaced by PE_448

//PE_503 replaced by PE_448

//PE_502 replaced by PE_448

//PE_501 replaced by PE_448

//PE_500 replaced by PE_448

//PE_499 replaced by PE_448

//PE_498 replaced by PE_448

//PE_497 replaced by PE_448

//PE_496 replaced by PE_448

//PE_495 replaced by PE_448

//PE_494 replaced by PE_448

//PE_493 replaced by PE_448

//PE_492 replaced by PE_448

//PE_491 replaced by PE_448

//PE_490 replaced by PE_448

//PE_489 replaced by PE_448

//PE_488 replaced by PE_448

//PE_487 replaced by PE_448

//PE_486 replaced by PE_448

//PE_485 replaced by PE_448

//PE_484 replaced by PE_448

//PE_483 replaced by PE_448

//PE_482 replaced by PE_448

//PE_481 replaced by PE_448

//PE_480 replaced by PE_448

//PE_479 replaced by PE_448

//PE_478 replaced by PE_448

//PE_477 replaced by PE_448

//PE_476 replaced by PE_448

//PE_475 replaced by PE_448

//PE_474 replaced by PE_448

//PE_473 replaced by PE_448

//PE_472 replaced by PE_448

//PE_471 replaced by PE_448

//PE_470 replaced by PE_448

//PE_469 replaced by PE_448

//PE_468 replaced by PE_448

//PE_467 replaced by PE_448

//PE_466 replaced by PE_448

//PE_465 replaced by PE_448

//PE_464 replaced by PE_448

//PE_463 replaced by PE_448

//PE_462 replaced by PE_448

//PE_461 replaced by PE_448

//PE_460 replaced by PE_448

//PE_459 replaced by PE_448

//PE_458 replaced by PE_448

//PE_457 replaced by PE_448

//PE_456 replaced by PE_448

//PE_455 replaced by PE_448

//PE_454 replaced by PE_448

//PE_453 replaced by PE_448

//PE_452 replaced by PE_448

//PE_451 replaced by PE_448

//PE_450 replaced by PE_448

//PE_449 replaced by PE_448

module PE_448 (
  input      [7:0]    activate,
  input      [7:0]    weight,
  input               valid,
  input      [15:0]   signCount,
  output     [7:0]    acount,
  output     [7:0]    bcount,
  output reg [31:0]   PE_OUT,
  output              finish,
  input               clk,
  input               reset
);

  wire       [15:0]   dsp_P;
  wire       [31:0]   _zz_reg1;
  wire       [31:0]   _zz_reg1_1;
  wire       [31:0]   _zz_reg1_2;
  reg        [31:0]   reg1;
  reg                 valid_regNext;
  reg                 valid_regNext_regNext;
  reg        [15:0]   finishCnt_count;
  wire                finishCnt_valid;
  reg                 valid_regNext_1;
  reg        [7:0]    activate_regNext;
  reg        [7:0]    weight_regNext;

  assign _zz_reg1 = {{16{dsp_P[15]}}, dsp_P};
  assign _zz_reg1_1 = 32'h0;
  assign _zz_reg1_2 = {{16{dsp_P[15]}}, dsp_P};
  dsp_marco dsp (
    .CLK (clk          ), //i
    .A   (activate[7:0]), //i
    .B   (weight[7:0]  ), //i
    .P   (dsp_P[15:0]  )  //o
  );
  assign finishCnt_valid = ((finishCnt_count == signCount) && valid_regNext_regNext);
  assign finish = finishCnt_valid;
  always @(*) begin
    PE_OUT = 32'h0;
    if(finishCnt_valid) begin
      PE_OUT = reg1;
    end
  end

  assign acount = activate_regNext;
  assign bcount = weight_regNext;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      reg1 <= 32'h0;
      finishCnt_count <= 16'h0;
    end else begin
      if(valid_regNext_regNext) begin
        if(finishCnt_valid) begin
          finishCnt_count <= 16'h0;
        end else begin
          finishCnt_count <= (finishCnt_count + 16'h0001);
        end
      end
      if(finishCnt_valid) begin
        reg1 <= (valid ? _zz_reg1 : _zz_reg1_1);
      end else begin
        if(valid_regNext_1) begin
          reg1 <= ($signed(_zz_reg1_2) + $signed(reg1));
        end
      end
    end
  end

  always @(posedge clk) begin
    valid_regNext <= valid;
    valid_regNext_regNext <= valid_regNext;
    valid_regNext_1 <= valid;
    activate_regNext <= activate;
    weight_regNext <= weight;
  end


endmodule
