// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : Weight_Cache
// Git hash  : 3ff479e98fb57df10a7ff9265112a692f55de7c4

`timescale 1ns/1ps

module Weight_Cache (
  input               start,
  input               sData_valid,
  output              sData_ready,
  input      [63:0]   sData_payload,
  input      [15:0]   Matrix_Row,
  input      [15:0]   Matrix_Col,
  output     [7:0]    mData_0,
  output     [7:0]    mData_1,
  output     [7:0]    mData_2,
  output     [7:0]    mData_3,
  output     [7:0]    mData_4,
  output     [7:0]    mData_5,
  output     [7:0]    mData_6,
  output     [7:0]    mData_7,
  output     [7:0]    mData_8,
  output     [7:0]    mData_9,
  output     [7:0]    mData_10,
  output     [7:0]    mData_11,
  output     [7:0]    mData_12,
  output     [7:0]    mData_13,
  output     [7:0]    mData_14,
  output     [7:0]    mData_15,
  output     [7:0]    mData_16,
  output     [7:0]    mData_17,
  output     [7:0]    mData_18,
  output     [7:0]    mData_19,
  output     [7:0]    mData_20,
  output     [7:0]    mData_21,
  output     [7:0]    mData_22,
  output     [7:0]    mData_23,
  output     [7:0]    mData_24,
  output     [7:0]    mData_25,
  output     [7:0]    mData_26,
  output     [7:0]    mData_27,
  output     [7:0]    mData_28,
  output     [7:0]    mData_29,
  output     [7:0]    mData_30,
  output     [7:0]    mData_31,
  output     [7:0]    mData_32,
  output     [7:0]    mData_33,
  output     [7:0]    mData_34,
  output     [7:0]    mData_35,
  output     [7:0]    mData_36,
  output     [7:0]    mData_37,
  output     [7:0]    mData_38,
  output     [7:0]    mData_39,
  output     [7:0]    mData_40,
  output     [7:0]    mData_41,
  output     [7:0]    mData_42,
  output     [7:0]    mData_43,
  output     [7:0]    mData_44,
  output     [7:0]    mData_45,
  output     [7:0]    mData_46,
  output     [7:0]    mData_47,
  output     [7:0]    mData_48,
  output     [7:0]    mData_49,
  output     [7:0]    mData_50,
  output     [7:0]    mData_51,
  output     [7:0]    mData_52,
  output     [7:0]    mData_53,
  output     [7:0]    mData_54,
  output     [7:0]    mData_55,
  output     [7:0]    mData_56,
  output     [7:0]    mData_57,
  output     [7:0]    mData_58,
  output     [7:0]    mData_59,
  output     [7:0]    mData_60,
  output     [7:0]    mData_61,
  output     [7:0]    mData_62,
  output     [7:0]    mData_63,
  output     [7:0]    mData_64,
  output     [7:0]    mData_65,
  output     [7:0]    mData_66,
  output     [7:0]    mData_67,
  output     [7:0]    mData_68,
  output     [7:0]    mData_69,
  output     [7:0]    mData_70,
  output     [7:0]    mData_71,
  output     [7:0]    mData_72,
  output     [7:0]    mData_73,
  output     [7:0]    mData_74,
  output     [7:0]    mData_75,
  output     [7:0]    mData_76,
  output     [7:0]    mData_77,
  output     [7:0]    mData_78,
  output     [7:0]    mData_79,
  output     [7:0]    mData_80,
  output     [7:0]    mData_81,
  output     [7:0]    mData_82,
  output     [7:0]    mData_83,
  output     [7:0]    mData_84,
  output     [7:0]    mData_85,
  output     [7:0]    mData_86,
  output     [7:0]    mData_87,
  output     [7:0]    mData_88,
  output     [7:0]    mData_89,
  output     [7:0]    mData_90,
  output     [7:0]    mData_91,
  output     [7:0]    mData_92,
  output     [7:0]    mData_93,
  output     [7:0]    mData_94,
  output     [7:0]    mData_95,
  output     [7:0]    mData_96,
  output     [7:0]    mData_97,
  output     [7:0]    mData_98,
  output     [7:0]    mData_99,
  output     [7:0]    mData_100,
  output     [7:0]    mData_101,
  output     [7:0]    mData_102,
  output     [7:0]    mData_103,
  output     [7:0]    mData_104,
  output     [7:0]    mData_105,
  output     [7:0]    mData_106,
  output     [7:0]    mData_107,
  output     [7:0]    mData_108,
  output     [7:0]    mData_109,
  output     [7:0]    mData_110,
  output     [7:0]    mData_111,
  output     [7:0]    mData_112,
  output     [7:0]    mData_113,
  output     [7:0]    mData_114,
  output     [7:0]    mData_115,
  output     [7:0]    mData_116,
  output     [7:0]    mData_117,
  output     [7:0]    mData_118,
  output     [7:0]    mData_119,
  output     [7:0]    mData_120,
  output     [7:0]    mData_121,
  output     [7:0]    mData_122,
  output     [7:0]    mData_123,
  output     [7:0]    mData_124,
  output     [7:0]    mData_125,
  output     [7:0]    mData_126,
  output     [7:0]    mData_127,
  output     [7:0]    mData_128,
  output     [7:0]    mData_129,
  output     [7:0]    mData_130,
  output     [7:0]    mData_131,
  output     [7:0]    mData_132,
  output     [7:0]    mData_133,
  output     [7:0]    mData_134,
  output     [7:0]    mData_135,
  output     [7:0]    mData_136,
  output     [7:0]    mData_137,
  output     [7:0]    mData_138,
  output     [7:0]    mData_139,
  output     [7:0]    mData_140,
  output     [7:0]    mData_141,
  output     [7:0]    mData_142,
  output     [7:0]    mData_143,
  output     [7:0]    mData_144,
  output     [7:0]    mData_145,
  output     [7:0]    mData_146,
  output     [7:0]    mData_147,
  output     [7:0]    mData_148,
  output     [7:0]    mData_149,
  output     [7:0]    mData_150,
  output     [7:0]    mData_151,
  output     [7:0]    mData_152,
  output     [7:0]    mData_153,
  output     [7:0]    mData_154,
  output     [7:0]    mData_155,
  output     [7:0]    mData_156,
  output     [7:0]    mData_157,
  output     [7:0]    mData_158,
  output     [7:0]    mData_159,
  output     [7:0]    mData_160,
  output     [7:0]    mData_161,
  output     [7:0]    mData_162,
  output     [7:0]    mData_163,
  output     [7:0]    mData_164,
  output     [7:0]    mData_165,
  output     [7:0]    mData_166,
  output     [7:0]    mData_167,
  output     [7:0]    mData_168,
  output     [7:0]    mData_169,
  output     [7:0]    mData_170,
  output     [7:0]    mData_171,
  output     [7:0]    mData_172,
  output     [7:0]    mData_173,
  output     [7:0]    mData_174,
  output     [7:0]    mData_175,
  output     [7:0]    mData_176,
  output     [7:0]    mData_177,
  output     [7:0]    mData_178,
  output     [7:0]    mData_179,
  output     [7:0]    mData_180,
  output     [7:0]    mData_181,
  output     [7:0]    mData_182,
  output     [7:0]    mData_183,
  output     [7:0]    mData_184,
  output     [7:0]    mData_185,
  output     [7:0]    mData_186,
  output     [7:0]    mData_187,
  output     [7:0]    mData_188,
  output     [7:0]    mData_189,
  output     [7:0]    mData_190,
  output     [7:0]    mData_191,
  output     [7:0]    mData_192,
  output     [7:0]    mData_193,
  output     [7:0]    mData_194,
  output     [7:0]    mData_195,
  output     [7:0]    mData_196,
  output     [7:0]    mData_197,
  output     [7:0]    mData_198,
  output     [7:0]    mData_199,
  output     [7:0]    mData_200,
  output     [7:0]    mData_201,
  output     [7:0]    mData_202,
  output     [7:0]    mData_203,
  output     [7:0]    mData_204,
  output     [7:0]    mData_205,
  output     [7:0]    mData_206,
  output     [7:0]    mData_207,
  output     [7:0]    mData_208,
  output     [7:0]    mData_209,
  output     [7:0]    mData_210,
  output     [7:0]    mData_211,
  output     [7:0]    mData_212,
  output     [7:0]    mData_213,
  output     [7:0]    mData_214,
  output     [7:0]    mData_215,
  output     [7:0]    mData_216,
  output     [7:0]    mData_217,
  output     [7:0]    mData_218,
  output     [7:0]    mData_219,
  output     [7:0]    mData_220,
  output     [7:0]    mData_221,
  output     [7:0]    mData_222,
  output     [7:0]    mData_223,
  output     [7:0]    mData_224,
  output     [7:0]    mData_225,
  output     [7:0]    mData_226,
  output     [7:0]    mData_227,
  output     [7:0]    mData_228,
  output     [7:0]    mData_229,
  output     [7:0]    mData_230,
  output     [7:0]    mData_231,
  output     [7:0]    mData_232,
  output     [7:0]    mData_233,
  output     [7:0]    mData_234,
  output     [7:0]    mData_235,
  output     [7:0]    mData_236,
  output     [7:0]    mData_237,
  output     [7:0]    mData_238,
  output     [7:0]    mData_239,
  output     [7:0]    mData_240,
  output     [7:0]    mData_241,
  output     [7:0]    mData_242,
  output     [7:0]    mData_243,
  output     [7:0]    mData_244,
  output     [7:0]    mData_245,
  output     [7:0]    mData_246,
  output     [7:0]    mData_247,
  output     [7:0]    mData_248,
  output     [7:0]    mData_249,
  output     [7:0]    mData_250,
  output     [7:0]    mData_251,
  output     [7:0]    mData_252,
  output     [7:0]    mData_253,
  output     [7:0]    mData_254,
  output     [7:0]    mData_255,
  output     [7:0]    mData_256,
  output     [7:0]    mData_257,
  output     [7:0]    mData_258,
  output     [7:0]    mData_259,
  output     [7:0]    mData_260,
  output     [7:0]    mData_261,
  output     [7:0]    mData_262,
  output     [7:0]    mData_263,
  output     [7:0]    mData_264,
  output     [7:0]    mData_265,
  output     [7:0]    mData_266,
  output     [7:0]    mData_267,
  output     [7:0]    mData_268,
  output     [7:0]    mData_269,
  output     [7:0]    mData_270,
  output     [7:0]    mData_271,
  output     [7:0]    mData_272,
  output     [7:0]    mData_273,
  output     [7:0]    mData_274,
  output     [7:0]    mData_275,
  output     [7:0]    mData_276,
  output     [7:0]    mData_277,
  output     [7:0]    mData_278,
  output     [7:0]    mData_279,
  output     [7:0]    mData_280,
  output     [7:0]    mData_281,
  output     [7:0]    mData_282,
  output     [7:0]    mData_283,
  output     [7:0]    mData_284,
  output     [7:0]    mData_285,
  output     [7:0]    mData_286,
  output     [7:0]    mData_287,
  output     [7:0]    mData_288,
  output     [7:0]    mData_289,
  output     [7:0]    mData_290,
  output     [7:0]    mData_291,
  output     [7:0]    mData_292,
  output     [7:0]    mData_293,
  output     [7:0]    mData_294,
  output     [7:0]    mData_295,
  output     [7:0]    mData_296,
  output     [7:0]    mData_297,
  output     [7:0]    mData_298,
  output     [7:0]    mData_299,
  output     [7:0]    mData_300,
  output     [7:0]    mData_301,
  output     [7:0]    mData_302,
  output     [7:0]    mData_303,
  output     [7:0]    mData_304,
  output     [7:0]    mData_305,
  output     [7:0]    mData_306,
  output     [7:0]    mData_307,
  output     [7:0]    mData_308,
  output     [7:0]    mData_309,
  output     [7:0]    mData_310,
  output     [7:0]    mData_311,
  output     [7:0]    mData_312,
  output     [7:0]    mData_313,
  output     [7:0]    mData_314,
  output     [7:0]    mData_315,
  output     [7:0]    mData_316,
  output     [7:0]    mData_317,
  output     [7:0]    mData_318,
  output     [7:0]    mData_319,
  output     [7:0]    mData_320,
  output     [7:0]    mData_321,
  output     [7:0]    mData_322,
  output     [7:0]    mData_323,
  output     [7:0]    mData_324,
  output     [7:0]    mData_325,
  output     [7:0]    mData_326,
  output     [7:0]    mData_327,
  output     [7:0]    mData_328,
  output     [7:0]    mData_329,
  output     [7:0]    mData_330,
  output     [7:0]    mData_331,
  output     [7:0]    mData_332,
  output     [7:0]    mData_333,
  output     [7:0]    mData_334,
  output     [7:0]    mData_335,
  output     [7:0]    mData_336,
  output     [7:0]    mData_337,
  output     [7:0]    mData_338,
  output     [7:0]    mData_339,
  output     [7:0]    mData_340,
  output     [7:0]    mData_341,
  output     [7:0]    mData_342,
  output     [7:0]    mData_343,
  output     [7:0]    mData_344,
  output     [7:0]    mData_345,
  output     [7:0]    mData_346,
  output     [7:0]    mData_347,
  output     [7:0]    mData_348,
  output     [7:0]    mData_349,
  output     [7:0]    mData_350,
  output     [7:0]    mData_351,
  output     [7:0]    mData_352,
  output     [7:0]    mData_353,
  output     [7:0]    mData_354,
  output     [7:0]    mData_355,
  output     [7:0]    mData_356,
  output     [7:0]    mData_357,
  output     [7:0]    mData_358,
  output     [7:0]    mData_359,
  output     [7:0]    mData_360,
  output     [7:0]    mData_361,
  output     [7:0]    mData_362,
  output     [7:0]    mData_363,
  output     [7:0]    mData_364,
  output     [7:0]    mData_365,
  output     [7:0]    mData_366,
  output     [7:0]    mData_367,
  output     [7:0]    mData_368,
  output     [7:0]    mData_369,
  output     [7:0]    mData_370,
  output     [7:0]    mData_371,
  output     [7:0]    mData_372,
  output     [7:0]    mData_373,
  output     [7:0]    mData_374,
  output     [7:0]    mData_375,
  output     [7:0]    mData_376,
  output     [7:0]    mData_377,
  output     [7:0]    mData_378,
  output     [7:0]    mData_379,
  output     [7:0]    mData_380,
  output     [7:0]    mData_381,
  output     [7:0]    mData_382,
  output     [7:0]    mData_383,
  output     [7:0]    mData_384,
  output     [7:0]    mData_385,
  output     [7:0]    mData_386,
  output     [7:0]    mData_387,
  output     [7:0]    mData_388,
  output     [7:0]    mData_389,
  output     [7:0]    mData_390,
  output     [7:0]    mData_391,
  output     [7:0]    mData_392,
  output     [7:0]    mData_393,
  output     [7:0]    mData_394,
  output     [7:0]    mData_395,
  output     [7:0]    mData_396,
  output     [7:0]    mData_397,
  output     [7:0]    mData_398,
  output     [7:0]    mData_399,
  output     [7:0]    mData_400,
  output     [7:0]    mData_401,
  output     [7:0]    mData_402,
  output     [7:0]    mData_403,
  output     [7:0]    mData_404,
  output     [7:0]    mData_405,
  output     [7:0]    mData_406,
  output     [7:0]    mData_407,
  output     [7:0]    mData_408,
  output     [7:0]    mData_409,
  output     [7:0]    mData_410,
  output     [7:0]    mData_411,
  output     [7:0]    mData_412,
  output     [7:0]    mData_413,
  output     [7:0]    mData_414,
  output     [7:0]    mData_415,
  output     [7:0]    mData_416,
  output     [7:0]    mData_417,
  output     [7:0]    mData_418,
  output     [7:0]    mData_419,
  output     [7:0]    mData_420,
  output     [7:0]    mData_421,
  output     [7:0]    mData_422,
  output     [7:0]    mData_423,
  output     [7:0]    mData_424,
  output     [7:0]    mData_425,
  output     [7:0]    mData_426,
  output     [7:0]    mData_427,
  output     [7:0]    mData_428,
  output     [7:0]    mData_429,
  output     [7:0]    mData_430,
  output     [7:0]    mData_431,
  output     [7:0]    mData_432,
  output     [7:0]    mData_433,
  output     [7:0]    mData_434,
  output     [7:0]    mData_435,
  output     [7:0]    mData_436,
  output     [7:0]    mData_437,
  output     [7:0]    mData_438,
  output     [7:0]    mData_439,
  output     [7:0]    mData_440,
  output     [7:0]    mData_441,
  output     [7:0]    mData_442,
  output     [7:0]    mData_443,
  output     [7:0]    mData_444,
  output     [7:0]    mData_445,
  output     [7:0]    mData_446,
  output     [7:0]    mData_447,
  output     [7:0]    mData_448,
  output     [7:0]    mData_449,
  output     [7:0]    mData_450,
  output     [7:0]    mData_451,
  output     [7:0]    mData_452,
  output     [7:0]    mData_453,
  output     [7:0]    mData_454,
  output     [7:0]    mData_455,
  output     [7:0]    mData_456,
  output     [7:0]    mData_457,
  output     [7:0]    mData_458,
  output     [7:0]    mData_459,
  output     [7:0]    mData_460,
  output     [7:0]    mData_461,
  output     [7:0]    mData_462,
  output     [7:0]    mData_463,
  output     [7:0]    mData_464,
  output     [7:0]    mData_465,
  output     [7:0]    mData_466,
  output     [7:0]    mData_467,
  output     [7:0]    mData_468,
  output     [7:0]    mData_469,
  output     [7:0]    mData_470,
  output     [7:0]    mData_471,
  output     [7:0]    mData_472,
  output     [7:0]    mData_473,
  output     [7:0]    mData_474,
  output     [7:0]    mData_475,
  output     [7:0]    mData_476,
  output     [7:0]    mData_477,
  output     [7:0]    mData_478,
  output     [7:0]    mData_479,
  output     [7:0]    mData_480,
  output     [7:0]    mData_481,
  output     [7:0]    mData_482,
  output     [7:0]    mData_483,
  output     [7:0]    mData_484,
  output     [7:0]    mData_485,
  output     [7:0]    mData_486,
  output     [7:0]    mData_487,
  output     [7:0]    mData_488,
  output     [7:0]    mData_489,
  output     [7:0]    mData_490,
  output     [7:0]    mData_491,
  output     [7:0]    mData_492,
  output     [7:0]    mData_493,
  output     [7:0]    mData_494,
  output     [7:0]    mData_495,
  output     [7:0]    mData_496,
  output     [7:0]    mData_497,
  output     [7:0]    mData_498,
  output     [7:0]    mData_499,
  output     [7:0]    mData_500,
  output     [7:0]    mData_501,
  output     [7:0]    mData_502,
  output     [7:0]    mData_503,
  output     [7:0]    mData_504,
  output     [7:0]    mData_505,
  output     [7:0]    mData_506,
  output     [7:0]    mData_507,
  output     [7:0]    mData_508,
  output     [7:0]    mData_509,
  output     [7:0]    mData_510,
  output     [7:0]    mData_511,
  input               Raddr_Valid,
  output              Weight_Cached,
  input               LayerEnd,
  output     [7:0]    MatrixCol_Switch,
  input               clk,
  input               reset
);
  localparam WEIGHT_CACHE_STATUS_IDLE = 4'd1;
  localparam WEIGHT_CACHE_STATUS_INIT = 4'd2;
  localparam WEIGHT_CACHE_STATUS_CACHE_WEIGHT = 4'd4;
  localparam WEIGHT_CACHE_STATUS_SA_COMPUTE = 4'd8;

  wire       [10:0]   xil_SimpleDualBram_addra;
  wire                xil_SimpleDualBram_ena;
  wire       [13:0]   xil_SimpleDualBram_addrb;
  wire       [10:0]   xil_SimpleDualBram_1_addra;
  wire                xil_SimpleDualBram_1_ena;
  wire       [13:0]   xil_SimpleDualBram_1_addrb;
  wire       [10:0]   xil_SimpleDualBram_2_addra;
  wire                xil_SimpleDualBram_2_ena;
  wire       [13:0]   xil_SimpleDualBram_2_addrb;
  wire       [10:0]   xil_SimpleDualBram_3_addra;
  wire                xil_SimpleDualBram_3_ena;
  wire       [13:0]   xil_SimpleDualBram_3_addrb;
  wire       [10:0]   xil_SimpleDualBram_4_addra;
  wire                xil_SimpleDualBram_4_ena;
  wire       [13:0]   xil_SimpleDualBram_4_addrb;
  wire       [10:0]   xil_SimpleDualBram_5_addra;
  wire                xil_SimpleDualBram_5_ena;
  wire       [13:0]   xil_SimpleDualBram_5_addrb;
  wire       [10:0]   xil_SimpleDualBram_6_addra;
  wire                xil_SimpleDualBram_6_ena;
  wire       [13:0]   xil_SimpleDualBram_6_addrb;
  wire       [10:0]   xil_SimpleDualBram_7_addra;
  wire                xil_SimpleDualBram_7_ena;
  wire       [13:0]   xil_SimpleDualBram_7_addrb;
  wire       [10:0]   xil_SimpleDualBram_8_addra;
  wire                xil_SimpleDualBram_8_ena;
  wire       [13:0]   xil_SimpleDualBram_8_addrb;
  wire       [10:0]   xil_SimpleDualBram_9_addra;
  wire                xil_SimpleDualBram_9_ena;
  wire       [13:0]   xil_SimpleDualBram_9_addrb;
  wire       [10:0]   xil_SimpleDualBram_10_addra;
  wire                xil_SimpleDualBram_10_ena;
  wire       [13:0]   xil_SimpleDualBram_10_addrb;
  wire       [10:0]   xil_SimpleDualBram_11_addra;
  wire                xil_SimpleDualBram_11_ena;
  wire       [13:0]   xil_SimpleDualBram_11_addrb;
  wire       [10:0]   xil_SimpleDualBram_12_addra;
  wire                xil_SimpleDualBram_12_ena;
  wire       [13:0]   xil_SimpleDualBram_12_addrb;
  wire       [10:0]   xil_SimpleDualBram_13_addra;
  wire                xil_SimpleDualBram_13_ena;
  wire       [13:0]   xil_SimpleDualBram_13_addrb;
  wire       [10:0]   xil_SimpleDualBram_14_addra;
  wire                xil_SimpleDualBram_14_ena;
  wire       [13:0]   xil_SimpleDualBram_14_addrb;
  wire       [10:0]   xil_SimpleDualBram_15_addra;
  wire                xil_SimpleDualBram_15_ena;
  wire       [13:0]   xil_SimpleDualBram_15_addrb;
  wire       [10:0]   xil_SimpleDualBram_16_addra;
  wire                xil_SimpleDualBram_16_ena;
  wire       [13:0]   xil_SimpleDualBram_16_addrb;
  wire       [10:0]   xil_SimpleDualBram_17_addra;
  wire                xil_SimpleDualBram_17_ena;
  wire       [13:0]   xil_SimpleDualBram_17_addrb;
  wire       [10:0]   xil_SimpleDualBram_18_addra;
  wire                xil_SimpleDualBram_18_ena;
  wire       [13:0]   xil_SimpleDualBram_18_addrb;
  wire       [10:0]   xil_SimpleDualBram_19_addra;
  wire                xil_SimpleDualBram_19_ena;
  wire       [13:0]   xil_SimpleDualBram_19_addrb;
  wire       [10:0]   xil_SimpleDualBram_20_addra;
  wire                xil_SimpleDualBram_20_ena;
  wire       [13:0]   xil_SimpleDualBram_20_addrb;
  wire       [10:0]   xil_SimpleDualBram_21_addra;
  wire                xil_SimpleDualBram_21_ena;
  wire       [13:0]   xil_SimpleDualBram_21_addrb;
  wire       [10:0]   xil_SimpleDualBram_22_addra;
  wire                xil_SimpleDualBram_22_ena;
  wire       [13:0]   xil_SimpleDualBram_22_addrb;
  wire       [10:0]   xil_SimpleDualBram_23_addra;
  wire                xil_SimpleDualBram_23_ena;
  wire       [13:0]   xil_SimpleDualBram_23_addrb;
  wire       [10:0]   xil_SimpleDualBram_24_addra;
  wire                xil_SimpleDualBram_24_ena;
  wire       [13:0]   xil_SimpleDualBram_24_addrb;
  wire       [10:0]   xil_SimpleDualBram_25_addra;
  wire                xil_SimpleDualBram_25_ena;
  wire       [13:0]   xil_SimpleDualBram_25_addrb;
  wire       [10:0]   xil_SimpleDualBram_26_addra;
  wire                xil_SimpleDualBram_26_ena;
  wire       [13:0]   xil_SimpleDualBram_26_addrb;
  wire       [10:0]   xil_SimpleDualBram_27_addra;
  wire                xil_SimpleDualBram_27_ena;
  wire       [13:0]   xil_SimpleDualBram_27_addrb;
  wire       [10:0]   xil_SimpleDualBram_28_addra;
  wire                xil_SimpleDualBram_28_ena;
  wire       [13:0]   xil_SimpleDualBram_28_addrb;
  wire       [10:0]   xil_SimpleDualBram_29_addra;
  wire                xil_SimpleDualBram_29_ena;
  wire       [13:0]   xil_SimpleDualBram_29_addrb;
  wire       [10:0]   xil_SimpleDualBram_30_addra;
  wire                xil_SimpleDualBram_30_ena;
  wire       [13:0]   xil_SimpleDualBram_30_addrb;
  wire       [10:0]   xil_SimpleDualBram_31_addra;
  wire                xil_SimpleDualBram_31_ena;
  wire       [13:0]   xil_SimpleDualBram_31_addrb;
  wire       [10:0]   xil_SimpleDualBram_32_addra;
  wire                xil_SimpleDualBram_32_ena;
  wire       [13:0]   xil_SimpleDualBram_32_addrb;
  wire       [10:0]   xil_SimpleDualBram_33_addra;
  wire                xil_SimpleDualBram_33_ena;
  wire       [13:0]   xil_SimpleDualBram_33_addrb;
  wire       [10:0]   xil_SimpleDualBram_34_addra;
  wire                xil_SimpleDualBram_34_ena;
  wire       [13:0]   xil_SimpleDualBram_34_addrb;
  wire       [10:0]   xil_SimpleDualBram_35_addra;
  wire                xil_SimpleDualBram_35_ena;
  wire       [13:0]   xil_SimpleDualBram_35_addrb;
  wire       [10:0]   xil_SimpleDualBram_36_addra;
  wire                xil_SimpleDualBram_36_ena;
  wire       [13:0]   xil_SimpleDualBram_36_addrb;
  wire       [10:0]   xil_SimpleDualBram_37_addra;
  wire                xil_SimpleDualBram_37_ena;
  wire       [13:0]   xil_SimpleDualBram_37_addrb;
  wire       [10:0]   xil_SimpleDualBram_38_addra;
  wire                xil_SimpleDualBram_38_ena;
  wire       [13:0]   xil_SimpleDualBram_38_addrb;
  wire       [10:0]   xil_SimpleDualBram_39_addra;
  wire                xil_SimpleDualBram_39_ena;
  wire       [13:0]   xil_SimpleDualBram_39_addrb;
  wire       [10:0]   xil_SimpleDualBram_40_addra;
  wire                xil_SimpleDualBram_40_ena;
  wire       [13:0]   xil_SimpleDualBram_40_addrb;
  wire       [10:0]   xil_SimpleDualBram_41_addra;
  wire                xil_SimpleDualBram_41_ena;
  wire       [13:0]   xil_SimpleDualBram_41_addrb;
  wire       [10:0]   xil_SimpleDualBram_42_addra;
  wire                xil_SimpleDualBram_42_ena;
  wire       [13:0]   xil_SimpleDualBram_42_addrb;
  wire       [10:0]   xil_SimpleDualBram_43_addra;
  wire                xil_SimpleDualBram_43_ena;
  wire       [13:0]   xil_SimpleDualBram_43_addrb;
  wire       [10:0]   xil_SimpleDualBram_44_addra;
  wire                xil_SimpleDualBram_44_ena;
  wire       [13:0]   xil_SimpleDualBram_44_addrb;
  wire       [10:0]   xil_SimpleDualBram_45_addra;
  wire                xil_SimpleDualBram_45_ena;
  wire       [13:0]   xil_SimpleDualBram_45_addrb;
  wire       [10:0]   xil_SimpleDualBram_46_addra;
  wire                xil_SimpleDualBram_46_ena;
  wire       [13:0]   xil_SimpleDualBram_46_addrb;
  wire       [10:0]   xil_SimpleDualBram_47_addra;
  wire                xil_SimpleDualBram_47_ena;
  wire       [13:0]   xil_SimpleDualBram_47_addrb;
  wire       [10:0]   xil_SimpleDualBram_48_addra;
  wire                xil_SimpleDualBram_48_ena;
  wire       [13:0]   xil_SimpleDualBram_48_addrb;
  wire       [10:0]   xil_SimpleDualBram_49_addra;
  wire                xil_SimpleDualBram_49_ena;
  wire       [13:0]   xil_SimpleDualBram_49_addrb;
  wire       [10:0]   xil_SimpleDualBram_50_addra;
  wire                xil_SimpleDualBram_50_ena;
  wire       [13:0]   xil_SimpleDualBram_50_addrb;
  wire       [10:0]   xil_SimpleDualBram_51_addra;
  wire                xil_SimpleDualBram_51_ena;
  wire       [13:0]   xil_SimpleDualBram_51_addrb;
  wire       [10:0]   xil_SimpleDualBram_52_addra;
  wire                xil_SimpleDualBram_52_ena;
  wire       [13:0]   xil_SimpleDualBram_52_addrb;
  wire       [10:0]   xil_SimpleDualBram_53_addra;
  wire                xil_SimpleDualBram_53_ena;
  wire       [13:0]   xil_SimpleDualBram_53_addrb;
  wire       [10:0]   xil_SimpleDualBram_54_addra;
  wire                xil_SimpleDualBram_54_ena;
  wire       [13:0]   xil_SimpleDualBram_54_addrb;
  wire       [10:0]   xil_SimpleDualBram_55_addra;
  wire                xil_SimpleDualBram_55_ena;
  wire       [13:0]   xil_SimpleDualBram_55_addrb;
  wire       [10:0]   xil_SimpleDualBram_56_addra;
  wire                xil_SimpleDualBram_56_ena;
  wire       [13:0]   xil_SimpleDualBram_56_addrb;
  wire       [10:0]   xil_SimpleDualBram_57_addra;
  wire                xil_SimpleDualBram_57_ena;
  wire       [13:0]   xil_SimpleDualBram_57_addrb;
  wire       [10:0]   xil_SimpleDualBram_58_addra;
  wire                xil_SimpleDualBram_58_ena;
  wire       [13:0]   xil_SimpleDualBram_58_addrb;
  wire       [10:0]   xil_SimpleDualBram_59_addra;
  wire                xil_SimpleDualBram_59_ena;
  wire       [13:0]   xil_SimpleDualBram_59_addrb;
  wire       [10:0]   xil_SimpleDualBram_60_addra;
  wire                xil_SimpleDualBram_60_ena;
  wire       [13:0]   xil_SimpleDualBram_60_addrb;
  wire       [10:0]   xil_SimpleDualBram_61_addra;
  wire                xil_SimpleDualBram_61_ena;
  wire       [13:0]   xil_SimpleDualBram_61_addrb;
  wire       [10:0]   xil_SimpleDualBram_62_addra;
  wire                xil_SimpleDualBram_62_ena;
  wire       [13:0]   xil_SimpleDualBram_62_addrb;
  wire       [10:0]   xil_SimpleDualBram_63_addra;
  wire                xil_SimpleDualBram_63_ena;
  wire       [13:0]   xil_SimpleDualBram_63_addrb;
  wire       [10:0]   xil_SimpleDualBram_64_addra;
  wire                xil_SimpleDualBram_64_ena;
  wire       [13:0]   xil_SimpleDualBram_64_addrb;
  wire       [10:0]   xil_SimpleDualBram_65_addra;
  wire                xil_SimpleDualBram_65_ena;
  wire       [13:0]   xil_SimpleDualBram_65_addrb;
  wire       [10:0]   xil_SimpleDualBram_66_addra;
  wire                xil_SimpleDualBram_66_ena;
  wire       [13:0]   xil_SimpleDualBram_66_addrb;
  wire       [10:0]   xil_SimpleDualBram_67_addra;
  wire                xil_SimpleDualBram_67_ena;
  wire       [13:0]   xil_SimpleDualBram_67_addrb;
  wire       [10:0]   xil_SimpleDualBram_68_addra;
  wire                xil_SimpleDualBram_68_ena;
  wire       [13:0]   xil_SimpleDualBram_68_addrb;
  wire       [10:0]   xil_SimpleDualBram_69_addra;
  wire                xil_SimpleDualBram_69_ena;
  wire       [13:0]   xil_SimpleDualBram_69_addrb;
  wire       [10:0]   xil_SimpleDualBram_70_addra;
  wire                xil_SimpleDualBram_70_ena;
  wire       [13:0]   xil_SimpleDualBram_70_addrb;
  wire       [10:0]   xil_SimpleDualBram_71_addra;
  wire                xil_SimpleDualBram_71_ena;
  wire       [13:0]   xil_SimpleDualBram_71_addrb;
  wire       [10:0]   xil_SimpleDualBram_72_addra;
  wire                xil_SimpleDualBram_72_ena;
  wire       [13:0]   xil_SimpleDualBram_72_addrb;
  wire       [10:0]   xil_SimpleDualBram_73_addra;
  wire                xil_SimpleDualBram_73_ena;
  wire       [13:0]   xil_SimpleDualBram_73_addrb;
  wire       [10:0]   xil_SimpleDualBram_74_addra;
  wire                xil_SimpleDualBram_74_ena;
  wire       [13:0]   xil_SimpleDualBram_74_addrb;
  wire       [10:0]   xil_SimpleDualBram_75_addra;
  wire                xil_SimpleDualBram_75_ena;
  wire       [13:0]   xil_SimpleDualBram_75_addrb;
  wire       [10:0]   xil_SimpleDualBram_76_addra;
  wire                xil_SimpleDualBram_76_ena;
  wire       [13:0]   xil_SimpleDualBram_76_addrb;
  wire       [10:0]   xil_SimpleDualBram_77_addra;
  wire                xil_SimpleDualBram_77_ena;
  wire       [13:0]   xil_SimpleDualBram_77_addrb;
  wire       [10:0]   xil_SimpleDualBram_78_addra;
  wire                xil_SimpleDualBram_78_ena;
  wire       [13:0]   xil_SimpleDualBram_78_addrb;
  wire       [10:0]   xil_SimpleDualBram_79_addra;
  wire                xil_SimpleDualBram_79_ena;
  wire       [13:0]   xil_SimpleDualBram_79_addrb;
  wire       [10:0]   xil_SimpleDualBram_80_addra;
  wire                xil_SimpleDualBram_80_ena;
  wire       [13:0]   xil_SimpleDualBram_80_addrb;
  wire       [10:0]   xil_SimpleDualBram_81_addra;
  wire                xil_SimpleDualBram_81_ena;
  wire       [13:0]   xil_SimpleDualBram_81_addrb;
  wire       [10:0]   xil_SimpleDualBram_82_addra;
  wire                xil_SimpleDualBram_82_ena;
  wire       [13:0]   xil_SimpleDualBram_82_addrb;
  wire       [10:0]   xil_SimpleDualBram_83_addra;
  wire                xil_SimpleDualBram_83_ena;
  wire       [13:0]   xil_SimpleDualBram_83_addrb;
  wire       [10:0]   xil_SimpleDualBram_84_addra;
  wire                xil_SimpleDualBram_84_ena;
  wire       [13:0]   xil_SimpleDualBram_84_addrb;
  wire       [10:0]   xil_SimpleDualBram_85_addra;
  wire                xil_SimpleDualBram_85_ena;
  wire       [13:0]   xil_SimpleDualBram_85_addrb;
  wire       [10:0]   xil_SimpleDualBram_86_addra;
  wire                xil_SimpleDualBram_86_ena;
  wire       [13:0]   xil_SimpleDualBram_86_addrb;
  wire       [10:0]   xil_SimpleDualBram_87_addra;
  wire                xil_SimpleDualBram_87_ena;
  wire       [13:0]   xil_SimpleDualBram_87_addrb;
  wire       [10:0]   xil_SimpleDualBram_88_addra;
  wire                xil_SimpleDualBram_88_ena;
  wire       [13:0]   xil_SimpleDualBram_88_addrb;
  wire       [10:0]   xil_SimpleDualBram_89_addra;
  wire                xil_SimpleDualBram_89_ena;
  wire       [13:0]   xil_SimpleDualBram_89_addrb;
  wire       [10:0]   xil_SimpleDualBram_90_addra;
  wire                xil_SimpleDualBram_90_ena;
  wire       [13:0]   xil_SimpleDualBram_90_addrb;
  wire       [10:0]   xil_SimpleDualBram_91_addra;
  wire                xil_SimpleDualBram_91_ena;
  wire       [13:0]   xil_SimpleDualBram_91_addrb;
  wire       [10:0]   xil_SimpleDualBram_92_addra;
  wire                xil_SimpleDualBram_92_ena;
  wire       [13:0]   xil_SimpleDualBram_92_addrb;
  wire       [10:0]   xil_SimpleDualBram_93_addra;
  wire                xil_SimpleDualBram_93_ena;
  wire       [13:0]   xil_SimpleDualBram_93_addrb;
  wire       [10:0]   xil_SimpleDualBram_94_addra;
  wire                xil_SimpleDualBram_94_ena;
  wire       [13:0]   xil_SimpleDualBram_94_addrb;
  wire       [10:0]   xil_SimpleDualBram_95_addra;
  wire                xil_SimpleDualBram_95_ena;
  wire       [13:0]   xil_SimpleDualBram_95_addrb;
  wire       [10:0]   xil_SimpleDualBram_96_addra;
  wire                xil_SimpleDualBram_96_ena;
  wire       [13:0]   xil_SimpleDualBram_96_addrb;
  wire       [10:0]   xil_SimpleDualBram_97_addra;
  wire                xil_SimpleDualBram_97_ena;
  wire       [13:0]   xil_SimpleDualBram_97_addrb;
  wire       [10:0]   xil_SimpleDualBram_98_addra;
  wire                xil_SimpleDualBram_98_ena;
  wire       [13:0]   xil_SimpleDualBram_98_addrb;
  wire       [10:0]   xil_SimpleDualBram_99_addra;
  wire                xil_SimpleDualBram_99_ena;
  wire       [13:0]   xil_SimpleDualBram_99_addrb;
  wire       [10:0]   xil_SimpleDualBram_100_addra;
  wire                xil_SimpleDualBram_100_ena;
  wire       [13:0]   xil_SimpleDualBram_100_addrb;
  wire       [10:0]   xil_SimpleDualBram_101_addra;
  wire                xil_SimpleDualBram_101_ena;
  wire       [13:0]   xil_SimpleDualBram_101_addrb;
  wire       [10:0]   xil_SimpleDualBram_102_addra;
  wire                xil_SimpleDualBram_102_ena;
  wire       [13:0]   xil_SimpleDualBram_102_addrb;
  wire       [10:0]   xil_SimpleDualBram_103_addra;
  wire                xil_SimpleDualBram_103_ena;
  wire       [13:0]   xil_SimpleDualBram_103_addrb;
  wire       [10:0]   xil_SimpleDualBram_104_addra;
  wire                xil_SimpleDualBram_104_ena;
  wire       [13:0]   xil_SimpleDualBram_104_addrb;
  wire       [10:0]   xil_SimpleDualBram_105_addra;
  wire                xil_SimpleDualBram_105_ena;
  wire       [13:0]   xil_SimpleDualBram_105_addrb;
  wire       [10:0]   xil_SimpleDualBram_106_addra;
  wire                xil_SimpleDualBram_106_ena;
  wire       [13:0]   xil_SimpleDualBram_106_addrb;
  wire       [10:0]   xil_SimpleDualBram_107_addra;
  wire                xil_SimpleDualBram_107_ena;
  wire       [13:0]   xil_SimpleDualBram_107_addrb;
  wire       [10:0]   xil_SimpleDualBram_108_addra;
  wire                xil_SimpleDualBram_108_ena;
  wire       [13:0]   xil_SimpleDualBram_108_addrb;
  wire       [10:0]   xil_SimpleDualBram_109_addra;
  wire                xil_SimpleDualBram_109_ena;
  wire       [13:0]   xil_SimpleDualBram_109_addrb;
  wire       [10:0]   xil_SimpleDualBram_110_addra;
  wire                xil_SimpleDualBram_110_ena;
  wire       [13:0]   xil_SimpleDualBram_110_addrb;
  wire       [10:0]   xil_SimpleDualBram_111_addra;
  wire                xil_SimpleDualBram_111_ena;
  wire       [13:0]   xil_SimpleDualBram_111_addrb;
  wire       [10:0]   xil_SimpleDualBram_112_addra;
  wire                xil_SimpleDualBram_112_ena;
  wire       [13:0]   xil_SimpleDualBram_112_addrb;
  wire       [10:0]   xil_SimpleDualBram_113_addra;
  wire                xil_SimpleDualBram_113_ena;
  wire       [13:0]   xil_SimpleDualBram_113_addrb;
  wire       [10:0]   xil_SimpleDualBram_114_addra;
  wire                xil_SimpleDualBram_114_ena;
  wire       [13:0]   xil_SimpleDualBram_114_addrb;
  wire       [10:0]   xil_SimpleDualBram_115_addra;
  wire                xil_SimpleDualBram_115_ena;
  wire       [13:0]   xil_SimpleDualBram_115_addrb;
  wire       [10:0]   xil_SimpleDualBram_116_addra;
  wire                xil_SimpleDualBram_116_ena;
  wire       [13:0]   xil_SimpleDualBram_116_addrb;
  wire       [10:0]   xil_SimpleDualBram_117_addra;
  wire                xil_SimpleDualBram_117_ena;
  wire       [13:0]   xil_SimpleDualBram_117_addrb;
  wire       [10:0]   xil_SimpleDualBram_118_addra;
  wire                xil_SimpleDualBram_118_ena;
  wire       [13:0]   xil_SimpleDualBram_118_addrb;
  wire       [10:0]   xil_SimpleDualBram_119_addra;
  wire                xil_SimpleDualBram_119_ena;
  wire       [13:0]   xil_SimpleDualBram_119_addrb;
  wire       [10:0]   xil_SimpleDualBram_120_addra;
  wire                xil_SimpleDualBram_120_ena;
  wire       [13:0]   xil_SimpleDualBram_120_addrb;
  wire       [10:0]   xil_SimpleDualBram_121_addra;
  wire                xil_SimpleDualBram_121_ena;
  wire       [13:0]   xil_SimpleDualBram_121_addrb;
  wire       [10:0]   xil_SimpleDualBram_122_addra;
  wire                xil_SimpleDualBram_122_ena;
  wire       [13:0]   xil_SimpleDualBram_122_addrb;
  wire       [10:0]   xil_SimpleDualBram_123_addra;
  wire                xil_SimpleDualBram_123_ena;
  wire       [13:0]   xil_SimpleDualBram_123_addrb;
  wire       [10:0]   xil_SimpleDualBram_124_addra;
  wire                xil_SimpleDualBram_124_ena;
  wire       [13:0]   xil_SimpleDualBram_124_addrb;
  wire       [10:0]   xil_SimpleDualBram_125_addra;
  wire                xil_SimpleDualBram_125_ena;
  wire       [13:0]   xil_SimpleDualBram_125_addrb;
  wire       [10:0]   xil_SimpleDualBram_126_addra;
  wire                xil_SimpleDualBram_126_ena;
  wire       [13:0]   xil_SimpleDualBram_126_addrb;
  wire       [10:0]   xil_SimpleDualBram_127_addra;
  wire                xil_SimpleDualBram_127_ena;
  wire       [13:0]   xil_SimpleDualBram_127_addrb;
  wire       [10:0]   xil_SimpleDualBram_128_addra;
  wire                xil_SimpleDualBram_128_ena;
  wire       [13:0]   xil_SimpleDualBram_128_addrb;
  wire       [10:0]   xil_SimpleDualBram_129_addra;
  wire                xil_SimpleDualBram_129_ena;
  wire       [13:0]   xil_SimpleDualBram_129_addrb;
  wire       [10:0]   xil_SimpleDualBram_130_addra;
  wire                xil_SimpleDualBram_130_ena;
  wire       [13:0]   xil_SimpleDualBram_130_addrb;
  wire       [10:0]   xil_SimpleDualBram_131_addra;
  wire                xil_SimpleDualBram_131_ena;
  wire       [13:0]   xil_SimpleDualBram_131_addrb;
  wire       [10:0]   xil_SimpleDualBram_132_addra;
  wire                xil_SimpleDualBram_132_ena;
  wire       [13:0]   xil_SimpleDualBram_132_addrb;
  wire       [10:0]   xil_SimpleDualBram_133_addra;
  wire                xil_SimpleDualBram_133_ena;
  wire       [13:0]   xil_SimpleDualBram_133_addrb;
  wire       [10:0]   xil_SimpleDualBram_134_addra;
  wire                xil_SimpleDualBram_134_ena;
  wire       [13:0]   xil_SimpleDualBram_134_addrb;
  wire       [10:0]   xil_SimpleDualBram_135_addra;
  wire                xil_SimpleDualBram_135_ena;
  wire       [13:0]   xil_SimpleDualBram_135_addrb;
  wire       [10:0]   xil_SimpleDualBram_136_addra;
  wire                xil_SimpleDualBram_136_ena;
  wire       [13:0]   xil_SimpleDualBram_136_addrb;
  wire       [10:0]   xil_SimpleDualBram_137_addra;
  wire                xil_SimpleDualBram_137_ena;
  wire       [13:0]   xil_SimpleDualBram_137_addrb;
  wire       [10:0]   xil_SimpleDualBram_138_addra;
  wire                xil_SimpleDualBram_138_ena;
  wire       [13:0]   xil_SimpleDualBram_138_addrb;
  wire       [10:0]   xil_SimpleDualBram_139_addra;
  wire                xil_SimpleDualBram_139_ena;
  wire       [13:0]   xil_SimpleDualBram_139_addrb;
  wire       [10:0]   xil_SimpleDualBram_140_addra;
  wire                xil_SimpleDualBram_140_ena;
  wire       [13:0]   xil_SimpleDualBram_140_addrb;
  wire       [10:0]   xil_SimpleDualBram_141_addra;
  wire                xil_SimpleDualBram_141_ena;
  wire       [13:0]   xil_SimpleDualBram_141_addrb;
  wire       [10:0]   xil_SimpleDualBram_142_addra;
  wire                xil_SimpleDualBram_142_ena;
  wire       [13:0]   xil_SimpleDualBram_142_addrb;
  wire       [10:0]   xil_SimpleDualBram_143_addra;
  wire                xil_SimpleDualBram_143_ena;
  wire       [13:0]   xil_SimpleDualBram_143_addrb;
  wire       [10:0]   xil_SimpleDualBram_144_addra;
  wire                xil_SimpleDualBram_144_ena;
  wire       [13:0]   xil_SimpleDualBram_144_addrb;
  wire       [10:0]   xil_SimpleDualBram_145_addra;
  wire                xil_SimpleDualBram_145_ena;
  wire       [13:0]   xil_SimpleDualBram_145_addrb;
  wire       [10:0]   xil_SimpleDualBram_146_addra;
  wire                xil_SimpleDualBram_146_ena;
  wire       [13:0]   xil_SimpleDualBram_146_addrb;
  wire       [10:0]   xil_SimpleDualBram_147_addra;
  wire                xil_SimpleDualBram_147_ena;
  wire       [13:0]   xil_SimpleDualBram_147_addrb;
  wire       [10:0]   xil_SimpleDualBram_148_addra;
  wire                xil_SimpleDualBram_148_ena;
  wire       [13:0]   xil_SimpleDualBram_148_addrb;
  wire       [10:0]   xil_SimpleDualBram_149_addra;
  wire                xil_SimpleDualBram_149_ena;
  wire       [13:0]   xil_SimpleDualBram_149_addrb;
  wire       [10:0]   xil_SimpleDualBram_150_addra;
  wire                xil_SimpleDualBram_150_ena;
  wire       [13:0]   xil_SimpleDualBram_150_addrb;
  wire       [10:0]   xil_SimpleDualBram_151_addra;
  wire                xil_SimpleDualBram_151_ena;
  wire       [13:0]   xil_SimpleDualBram_151_addrb;
  wire       [10:0]   xil_SimpleDualBram_152_addra;
  wire                xil_SimpleDualBram_152_ena;
  wire       [13:0]   xil_SimpleDualBram_152_addrb;
  wire       [10:0]   xil_SimpleDualBram_153_addra;
  wire                xil_SimpleDualBram_153_ena;
  wire       [13:0]   xil_SimpleDualBram_153_addrb;
  wire       [10:0]   xil_SimpleDualBram_154_addra;
  wire                xil_SimpleDualBram_154_ena;
  wire       [13:0]   xil_SimpleDualBram_154_addrb;
  wire       [10:0]   xil_SimpleDualBram_155_addra;
  wire                xil_SimpleDualBram_155_ena;
  wire       [13:0]   xil_SimpleDualBram_155_addrb;
  wire       [10:0]   xil_SimpleDualBram_156_addra;
  wire                xil_SimpleDualBram_156_ena;
  wire       [13:0]   xil_SimpleDualBram_156_addrb;
  wire       [10:0]   xil_SimpleDualBram_157_addra;
  wire                xil_SimpleDualBram_157_ena;
  wire       [13:0]   xil_SimpleDualBram_157_addrb;
  wire       [10:0]   xil_SimpleDualBram_158_addra;
  wire                xil_SimpleDualBram_158_ena;
  wire       [13:0]   xil_SimpleDualBram_158_addrb;
  wire       [10:0]   xil_SimpleDualBram_159_addra;
  wire                xil_SimpleDualBram_159_ena;
  wire       [13:0]   xil_SimpleDualBram_159_addrb;
  wire       [10:0]   xil_SimpleDualBram_160_addra;
  wire                xil_SimpleDualBram_160_ena;
  wire       [13:0]   xil_SimpleDualBram_160_addrb;
  wire       [10:0]   xil_SimpleDualBram_161_addra;
  wire                xil_SimpleDualBram_161_ena;
  wire       [13:0]   xil_SimpleDualBram_161_addrb;
  wire       [10:0]   xil_SimpleDualBram_162_addra;
  wire                xil_SimpleDualBram_162_ena;
  wire       [13:0]   xil_SimpleDualBram_162_addrb;
  wire       [10:0]   xil_SimpleDualBram_163_addra;
  wire                xil_SimpleDualBram_163_ena;
  wire       [13:0]   xil_SimpleDualBram_163_addrb;
  wire       [10:0]   xil_SimpleDualBram_164_addra;
  wire                xil_SimpleDualBram_164_ena;
  wire       [13:0]   xil_SimpleDualBram_164_addrb;
  wire       [10:0]   xil_SimpleDualBram_165_addra;
  wire                xil_SimpleDualBram_165_ena;
  wire       [13:0]   xil_SimpleDualBram_165_addrb;
  wire       [10:0]   xil_SimpleDualBram_166_addra;
  wire                xil_SimpleDualBram_166_ena;
  wire       [13:0]   xil_SimpleDualBram_166_addrb;
  wire       [10:0]   xil_SimpleDualBram_167_addra;
  wire                xil_SimpleDualBram_167_ena;
  wire       [13:0]   xil_SimpleDualBram_167_addrb;
  wire       [10:0]   xil_SimpleDualBram_168_addra;
  wire                xil_SimpleDualBram_168_ena;
  wire       [13:0]   xil_SimpleDualBram_168_addrb;
  wire       [10:0]   xil_SimpleDualBram_169_addra;
  wire                xil_SimpleDualBram_169_ena;
  wire       [13:0]   xil_SimpleDualBram_169_addrb;
  wire       [10:0]   xil_SimpleDualBram_170_addra;
  wire                xil_SimpleDualBram_170_ena;
  wire       [13:0]   xil_SimpleDualBram_170_addrb;
  wire       [10:0]   xil_SimpleDualBram_171_addra;
  wire                xil_SimpleDualBram_171_ena;
  wire       [13:0]   xil_SimpleDualBram_171_addrb;
  wire       [10:0]   xil_SimpleDualBram_172_addra;
  wire                xil_SimpleDualBram_172_ena;
  wire       [13:0]   xil_SimpleDualBram_172_addrb;
  wire       [10:0]   xil_SimpleDualBram_173_addra;
  wire                xil_SimpleDualBram_173_ena;
  wire       [13:0]   xil_SimpleDualBram_173_addrb;
  wire       [10:0]   xil_SimpleDualBram_174_addra;
  wire                xil_SimpleDualBram_174_ena;
  wire       [13:0]   xil_SimpleDualBram_174_addrb;
  wire       [10:0]   xil_SimpleDualBram_175_addra;
  wire                xil_SimpleDualBram_175_ena;
  wire       [13:0]   xil_SimpleDualBram_175_addrb;
  wire       [10:0]   xil_SimpleDualBram_176_addra;
  wire                xil_SimpleDualBram_176_ena;
  wire       [13:0]   xil_SimpleDualBram_176_addrb;
  wire       [10:0]   xil_SimpleDualBram_177_addra;
  wire                xil_SimpleDualBram_177_ena;
  wire       [13:0]   xil_SimpleDualBram_177_addrb;
  wire       [10:0]   xil_SimpleDualBram_178_addra;
  wire                xil_SimpleDualBram_178_ena;
  wire       [13:0]   xil_SimpleDualBram_178_addrb;
  wire       [10:0]   xil_SimpleDualBram_179_addra;
  wire                xil_SimpleDualBram_179_ena;
  wire       [13:0]   xil_SimpleDualBram_179_addrb;
  wire       [10:0]   xil_SimpleDualBram_180_addra;
  wire                xil_SimpleDualBram_180_ena;
  wire       [13:0]   xil_SimpleDualBram_180_addrb;
  wire       [10:0]   xil_SimpleDualBram_181_addra;
  wire                xil_SimpleDualBram_181_ena;
  wire       [13:0]   xil_SimpleDualBram_181_addrb;
  wire       [10:0]   xil_SimpleDualBram_182_addra;
  wire                xil_SimpleDualBram_182_ena;
  wire       [13:0]   xil_SimpleDualBram_182_addrb;
  wire       [10:0]   xil_SimpleDualBram_183_addra;
  wire                xil_SimpleDualBram_183_ena;
  wire       [13:0]   xil_SimpleDualBram_183_addrb;
  wire       [10:0]   xil_SimpleDualBram_184_addra;
  wire                xil_SimpleDualBram_184_ena;
  wire       [13:0]   xil_SimpleDualBram_184_addrb;
  wire       [10:0]   xil_SimpleDualBram_185_addra;
  wire                xil_SimpleDualBram_185_ena;
  wire       [13:0]   xil_SimpleDualBram_185_addrb;
  wire       [10:0]   xil_SimpleDualBram_186_addra;
  wire                xil_SimpleDualBram_186_ena;
  wire       [13:0]   xil_SimpleDualBram_186_addrb;
  wire       [10:0]   xil_SimpleDualBram_187_addra;
  wire                xil_SimpleDualBram_187_ena;
  wire       [13:0]   xil_SimpleDualBram_187_addrb;
  wire       [10:0]   xil_SimpleDualBram_188_addra;
  wire                xil_SimpleDualBram_188_ena;
  wire       [13:0]   xil_SimpleDualBram_188_addrb;
  wire       [10:0]   xil_SimpleDualBram_189_addra;
  wire                xil_SimpleDualBram_189_ena;
  wire       [13:0]   xil_SimpleDualBram_189_addrb;
  wire       [10:0]   xil_SimpleDualBram_190_addra;
  wire                xil_SimpleDualBram_190_ena;
  wire       [13:0]   xil_SimpleDualBram_190_addrb;
  wire       [10:0]   xil_SimpleDualBram_191_addra;
  wire                xil_SimpleDualBram_191_ena;
  wire       [13:0]   xil_SimpleDualBram_191_addrb;
  wire       [10:0]   xil_SimpleDualBram_192_addra;
  wire                xil_SimpleDualBram_192_ena;
  wire       [13:0]   xil_SimpleDualBram_192_addrb;
  wire       [10:0]   xil_SimpleDualBram_193_addra;
  wire                xil_SimpleDualBram_193_ena;
  wire       [13:0]   xil_SimpleDualBram_193_addrb;
  wire       [10:0]   xil_SimpleDualBram_194_addra;
  wire                xil_SimpleDualBram_194_ena;
  wire       [13:0]   xil_SimpleDualBram_194_addrb;
  wire       [10:0]   xil_SimpleDualBram_195_addra;
  wire                xil_SimpleDualBram_195_ena;
  wire       [13:0]   xil_SimpleDualBram_195_addrb;
  wire       [10:0]   xil_SimpleDualBram_196_addra;
  wire                xil_SimpleDualBram_196_ena;
  wire       [13:0]   xil_SimpleDualBram_196_addrb;
  wire       [10:0]   xil_SimpleDualBram_197_addra;
  wire                xil_SimpleDualBram_197_ena;
  wire       [13:0]   xil_SimpleDualBram_197_addrb;
  wire       [10:0]   xil_SimpleDualBram_198_addra;
  wire                xil_SimpleDualBram_198_ena;
  wire       [13:0]   xil_SimpleDualBram_198_addrb;
  wire       [10:0]   xil_SimpleDualBram_199_addra;
  wire                xil_SimpleDualBram_199_ena;
  wire       [13:0]   xil_SimpleDualBram_199_addrb;
  wire       [10:0]   xil_SimpleDualBram_200_addra;
  wire                xil_SimpleDualBram_200_ena;
  wire       [13:0]   xil_SimpleDualBram_200_addrb;
  wire       [10:0]   xil_SimpleDualBram_201_addra;
  wire                xil_SimpleDualBram_201_ena;
  wire       [13:0]   xil_SimpleDualBram_201_addrb;
  wire       [10:0]   xil_SimpleDualBram_202_addra;
  wire                xil_SimpleDualBram_202_ena;
  wire       [13:0]   xil_SimpleDualBram_202_addrb;
  wire       [10:0]   xil_SimpleDualBram_203_addra;
  wire                xil_SimpleDualBram_203_ena;
  wire       [13:0]   xil_SimpleDualBram_203_addrb;
  wire       [10:0]   xil_SimpleDualBram_204_addra;
  wire                xil_SimpleDualBram_204_ena;
  wire       [13:0]   xil_SimpleDualBram_204_addrb;
  wire       [10:0]   xil_SimpleDualBram_205_addra;
  wire                xil_SimpleDualBram_205_ena;
  wire       [13:0]   xil_SimpleDualBram_205_addrb;
  wire       [10:0]   xil_SimpleDualBram_206_addra;
  wire                xil_SimpleDualBram_206_ena;
  wire       [13:0]   xil_SimpleDualBram_206_addrb;
  wire       [10:0]   xil_SimpleDualBram_207_addra;
  wire                xil_SimpleDualBram_207_ena;
  wire       [13:0]   xil_SimpleDualBram_207_addrb;
  wire       [10:0]   xil_SimpleDualBram_208_addra;
  wire                xil_SimpleDualBram_208_ena;
  wire       [13:0]   xil_SimpleDualBram_208_addrb;
  wire       [10:0]   xil_SimpleDualBram_209_addra;
  wire                xil_SimpleDualBram_209_ena;
  wire       [13:0]   xil_SimpleDualBram_209_addrb;
  wire       [10:0]   xil_SimpleDualBram_210_addra;
  wire                xil_SimpleDualBram_210_ena;
  wire       [13:0]   xil_SimpleDualBram_210_addrb;
  wire       [10:0]   xil_SimpleDualBram_211_addra;
  wire                xil_SimpleDualBram_211_ena;
  wire       [13:0]   xil_SimpleDualBram_211_addrb;
  wire       [10:0]   xil_SimpleDualBram_212_addra;
  wire                xil_SimpleDualBram_212_ena;
  wire       [13:0]   xil_SimpleDualBram_212_addrb;
  wire       [10:0]   xil_SimpleDualBram_213_addra;
  wire                xil_SimpleDualBram_213_ena;
  wire       [13:0]   xil_SimpleDualBram_213_addrb;
  wire       [10:0]   xil_SimpleDualBram_214_addra;
  wire                xil_SimpleDualBram_214_ena;
  wire       [13:0]   xil_SimpleDualBram_214_addrb;
  wire       [10:0]   xil_SimpleDualBram_215_addra;
  wire                xil_SimpleDualBram_215_ena;
  wire       [13:0]   xil_SimpleDualBram_215_addrb;
  wire       [10:0]   xil_SimpleDualBram_216_addra;
  wire                xil_SimpleDualBram_216_ena;
  wire       [13:0]   xil_SimpleDualBram_216_addrb;
  wire       [10:0]   xil_SimpleDualBram_217_addra;
  wire                xil_SimpleDualBram_217_ena;
  wire       [13:0]   xil_SimpleDualBram_217_addrb;
  wire       [10:0]   xil_SimpleDualBram_218_addra;
  wire                xil_SimpleDualBram_218_ena;
  wire       [13:0]   xil_SimpleDualBram_218_addrb;
  wire       [10:0]   xil_SimpleDualBram_219_addra;
  wire                xil_SimpleDualBram_219_ena;
  wire       [13:0]   xil_SimpleDualBram_219_addrb;
  wire       [10:0]   xil_SimpleDualBram_220_addra;
  wire                xil_SimpleDualBram_220_ena;
  wire       [13:0]   xil_SimpleDualBram_220_addrb;
  wire       [10:0]   xil_SimpleDualBram_221_addra;
  wire                xil_SimpleDualBram_221_ena;
  wire       [13:0]   xil_SimpleDualBram_221_addrb;
  wire       [10:0]   xil_SimpleDualBram_222_addra;
  wire                xil_SimpleDualBram_222_ena;
  wire       [13:0]   xil_SimpleDualBram_222_addrb;
  wire       [10:0]   xil_SimpleDualBram_223_addra;
  wire                xil_SimpleDualBram_223_ena;
  wire       [13:0]   xil_SimpleDualBram_223_addrb;
  wire       [10:0]   xil_SimpleDualBram_224_addra;
  wire                xil_SimpleDualBram_224_ena;
  wire       [13:0]   xil_SimpleDualBram_224_addrb;
  wire       [10:0]   xil_SimpleDualBram_225_addra;
  wire                xil_SimpleDualBram_225_ena;
  wire       [13:0]   xil_SimpleDualBram_225_addrb;
  wire       [10:0]   xil_SimpleDualBram_226_addra;
  wire                xil_SimpleDualBram_226_ena;
  wire       [13:0]   xil_SimpleDualBram_226_addrb;
  wire       [10:0]   xil_SimpleDualBram_227_addra;
  wire                xil_SimpleDualBram_227_ena;
  wire       [13:0]   xil_SimpleDualBram_227_addrb;
  wire       [10:0]   xil_SimpleDualBram_228_addra;
  wire                xil_SimpleDualBram_228_ena;
  wire       [13:0]   xil_SimpleDualBram_228_addrb;
  wire       [10:0]   xil_SimpleDualBram_229_addra;
  wire                xil_SimpleDualBram_229_ena;
  wire       [13:0]   xil_SimpleDualBram_229_addrb;
  wire       [10:0]   xil_SimpleDualBram_230_addra;
  wire                xil_SimpleDualBram_230_ena;
  wire       [13:0]   xil_SimpleDualBram_230_addrb;
  wire       [10:0]   xil_SimpleDualBram_231_addra;
  wire                xil_SimpleDualBram_231_ena;
  wire       [13:0]   xil_SimpleDualBram_231_addrb;
  wire       [10:0]   xil_SimpleDualBram_232_addra;
  wire                xil_SimpleDualBram_232_ena;
  wire       [13:0]   xil_SimpleDualBram_232_addrb;
  wire       [10:0]   xil_SimpleDualBram_233_addra;
  wire                xil_SimpleDualBram_233_ena;
  wire       [13:0]   xil_SimpleDualBram_233_addrb;
  wire       [10:0]   xil_SimpleDualBram_234_addra;
  wire                xil_SimpleDualBram_234_ena;
  wire       [13:0]   xil_SimpleDualBram_234_addrb;
  wire       [10:0]   xil_SimpleDualBram_235_addra;
  wire                xil_SimpleDualBram_235_ena;
  wire       [13:0]   xil_SimpleDualBram_235_addrb;
  wire       [10:0]   xil_SimpleDualBram_236_addra;
  wire                xil_SimpleDualBram_236_ena;
  wire       [13:0]   xil_SimpleDualBram_236_addrb;
  wire       [10:0]   xil_SimpleDualBram_237_addra;
  wire                xil_SimpleDualBram_237_ena;
  wire       [13:0]   xil_SimpleDualBram_237_addrb;
  wire       [10:0]   xil_SimpleDualBram_238_addra;
  wire                xil_SimpleDualBram_238_ena;
  wire       [13:0]   xil_SimpleDualBram_238_addrb;
  wire       [10:0]   xil_SimpleDualBram_239_addra;
  wire                xil_SimpleDualBram_239_ena;
  wire       [13:0]   xil_SimpleDualBram_239_addrb;
  wire       [10:0]   xil_SimpleDualBram_240_addra;
  wire                xil_SimpleDualBram_240_ena;
  wire       [13:0]   xil_SimpleDualBram_240_addrb;
  wire       [10:0]   xil_SimpleDualBram_241_addra;
  wire                xil_SimpleDualBram_241_ena;
  wire       [13:0]   xil_SimpleDualBram_241_addrb;
  wire       [10:0]   xil_SimpleDualBram_242_addra;
  wire                xil_SimpleDualBram_242_ena;
  wire       [13:0]   xil_SimpleDualBram_242_addrb;
  wire       [10:0]   xil_SimpleDualBram_243_addra;
  wire                xil_SimpleDualBram_243_ena;
  wire       [13:0]   xil_SimpleDualBram_243_addrb;
  wire       [10:0]   xil_SimpleDualBram_244_addra;
  wire                xil_SimpleDualBram_244_ena;
  wire       [13:0]   xil_SimpleDualBram_244_addrb;
  wire       [10:0]   xil_SimpleDualBram_245_addra;
  wire                xil_SimpleDualBram_245_ena;
  wire       [13:0]   xil_SimpleDualBram_245_addrb;
  wire       [10:0]   xil_SimpleDualBram_246_addra;
  wire                xil_SimpleDualBram_246_ena;
  wire       [13:0]   xil_SimpleDualBram_246_addrb;
  wire       [10:0]   xil_SimpleDualBram_247_addra;
  wire                xil_SimpleDualBram_247_ena;
  wire       [13:0]   xil_SimpleDualBram_247_addrb;
  wire       [10:0]   xil_SimpleDualBram_248_addra;
  wire                xil_SimpleDualBram_248_ena;
  wire       [13:0]   xil_SimpleDualBram_248_addrb;
  wire       [10:0]   xil_SimpleDualBram_249_addra;
  wire                xil_SimpleDualBram_249_ena;
  wire       [13:0]   xil_SimpleDualBram_249_addrb;
  wire       [10:0]   xil_SimpleDualBram_250_addra;
  wire                xil_SimpleDualBram_250_ena;
  wire       [13:0]   xil_SimpleDualBram_250_addrb;
  wire       [10:0]   xil_SimpleDualBram_251_addra;
  wire                xil_SimpleDualBram_251_ena;
  wire       [13:0]   xil_SimpleDualBram_251_addrb;
  wire       [10:0]   xil_SimpleDualBram_252_addra;
  wire                xil_SimpleDualBram_252_ena;
  wire       [13:0]   xil_SimpleDualBram_252_addrb;
  wire       [10:0]   xil_SimpleDualBram_253_addra;
  wire                xil_SimpleDualBram_253_ena;
  wire       [13:0]   xil_SimpleDualBram_253_addrb;
  wire       [10:0]   xil_SimpleDualBram_254_addra;
  wire                xil_SimpleDualBram_254_ena;
  wire       [13:0]   xil_SimpleDualBram_254_addrb;
  wire       [10:0]   xil_SimpleDualBram_255_addra;
  wire                xil_SimpleDualBram_255_ena;
  wire       [13:0]   xil_SimpleDualBram_255_addrb;
  wire       [10:0]   xil_SimpleDualBram_256_addra;
  wire                xil_SimpleDualBram_256_ena;
  wire       [13:0]   xil_SimpleDualBram_256_addrb;
  wire       [10:0]   xil_SimpleDualBram_257_addra;
  wire                xil_SimpleDualBram_257_ena;
  wire       [13:0]   xil_SimpleDualBram_257_addrb;
  wire       [10:0]   xil_SimpleDualBram_258_addra;
  wire                xil_SimpleDualBram_258_ena;
  wire       [13:0]   xil_SimpleDualBram_258_addrb;
  wire       [10:0]   xil_SimpleDualBram_259_addra;
  wire                xil_SimpleDualBram_259_ena;
  wire       [13:0]   xil_SimpleDualBram_259_addrb;
  wire       [10:0]   xil_SimpleDualBram_260_addra;
  wire                xil_SimpleDualBram_260_ena;
  wire       [13:0]   xil_SimpleDualBram_260_addrb;
  wire       [10:0]   xil_SimpleDualBram_261_addra;
  wire                xil_SimpleDualBram_261_ena;
  wire       [13:0]   xil_SimpleDualBram_261_addrb;
  wire       [10:0]   xil_SimpleDualBram_262_addra;
  wire                xil_SimpleDualBram_262_ena;
  wire       [13:0]   xil_SimpleDualBram_262_addrb;
  wire       [10:0]   xil_SimpleDualBram_263_addra;
  wire                xil_SimpleDualBram_263_ena;
  wire       [13:0]   xil_SimpleDualBram_263_addrb;
  wire       [10:0]   xil_SimpleDualBram_264_addra;
  wire                xil_SimpleDualBram_264_ena;
  wire       [13:0]   xil_SimpleDualBram_264_addrb;
  wire       [10:0]   xil_SimpleDualBram_265_addra;
  wire                xil_SimpleDualBram_265_ena;
  wire       [13:0]   xil_SimpleDualBram_265_addrb;
  wire       [10:0]   xil_SimpleDualBram_266_addra;
  wire                xil_SimpleDualBram_266_ena;
  wire       [13:0]   xil_SimpleDualBram_266_addrb;
  wire       [10:0]   xil_SimpleDualBram_267_addra;
  wire                xil_SimpleDualBram_267_ena;
  wire       [13:0]   xil_SimpleDualBram_267_addrb;
  wire       [10:0]   xil_SimpleDualBram_268_addra;
  wire                xil_SimpleDualBram_268_ena;
  wire       [13:0]   xil_SimpleDualBram_268_addrb;
  wire       [10:0]   xil_SimpleDualBram_269_addra;
  wire                xil_SimpleDualBram_269_ena;
  wire       [13:0]   xil_SimpleDualBram_269_addrb;
  wire       [10:0]   xil_SimpleDualBram_270_addra;
  wire                xil_SimpleDualBram_270_ena;
  wire       [13:0]   xil_SimpleDualBram_270_addrb;
  wire       [10:0]   xil_SimpleDualBram_271_addra;
  wire                xil_SimpleDualBram_271_ena;
  wire       [13:0]   xil_SimpleDualBram_271_addrb;
  wire       [10:0]   xil_SimpleDualBram_272_addra;
  wire                xil_SimpleDualBram_272_ena;
  wire       [13:0]   xil_SimpleDualBram_272_addrb;
  wire       [10:0]   xil_SimpleDualBram_273_addra;
  wire                xil_SimpleDualBram_273_ena;
  wire       [13:0]   xil_SimpleDualBram_273_addrb;
  wire       [10:0]   xil_SimpleDualBram_274_addra;
  wire                xil_SimpleDualBram_274_ena;
  wire       [13:0]   xil_SimpleDualBram_274_addrb;
  wire       [10:0]   xil_SimpleDualBram_275_addra;
  wire                xil_SimpleDualBram_275_ena;
  wire       [13:0]   xil_SimpleDualBram_275_addrb;
  wire       [10:0]   xil_SimpleDualBram_276_addra;
  wire                xil_SimpleDualBram_276_ena;
  wire       [13:0]   xil_SimpleDualBram_276_addrb;
  wire       [10:0]   xil_SimpleDualBram_277_addra;
  wire                xil_SimpleDualBram_277_ena;
  wire       [13:0]   xil_SimpleDualBram_277_addrb;
  wire       [10:0]   xil_SimpleDualBram_278_addra;
  wire                xil_SimpleDualBram_278_ena;
  wire       [13:0]   xil_SimpleDualBram_278_addrb;
  wire       [10:0]   xil_SimpleDualBram_279_addra;
  wire                xil_SimpleDualBram_279_ena;
  wire       [13:0]   xil_SimpleDualBram_279_addrb;
  wire       [10:0]   xil_SimpleDualBram_280_addra;
  wire                xil_SimpleDualBram_280_ena;
  wire       [13:0]   xil_SimpleDualBram_280_addrb;
  wire       [10:0]   xil_SimpleDualBram_281_addra;
  wire                xil_SimpleDualBram_281_ena;
  wire       [13:0]   xil_SimpleDualBram_281_addrb;
  wire       [10:0]   xil_SimpleDualBram_282_addra;
  wire                xil_SimpleDualBram_282_ena;
  wire       [13:0]   xil_SimpleDualBram_282_addrb;
  wire       [10:0]   xil_SimpleDualBram_283_addra;
  wire                xil_SimpleDualBram_283_ena;
  wire       [13:0]   xil_SimpleDualBram_283_addrb;
  wire       [10:0]   xil_SimpleDualBram_284_addra;
  wire                xil_SimpleDualBram_284_ena;
  wire       [13:0]   xil_SimpleDualBram_284_addrb;
  wire       [10:0]   xil_SimpleDualBram_285_addra;
  wire                xil_SimpleDualBram_285_ena;
  wire       [13:0]   xil_SimpleDualBram_285_addrb;
  wire       [10:0]   xil_SimpleDualBram_286_addra;
  wire                xil_SimpleDualBram_286_ena;
  wire       [13:0]   xil_SimpleDualBram_286_addrb;
  wire       [10:0]   xil_SimpleDualBram_287_addra;
  wire                xil_SimpleDualBram_287_ena;
  wire       [13:0]   xil_SimpleDualBram_287_addrb;
  wire       [10:0]   xil_SimpleDualBram_288_addra;
  wire                xil_SimpleDualBram_288_ena;
  wire       [13:0]   xil_SimpleDualBram_288_addrb;
  wire       [10:0]   xil_SimpleDualBram_289_addra;
  wire                xil_SimpleDualBram_289_ena;
  wire       [13:0]   xil_SimpleDualBram_289_addrb;
  wire       [10:0]   xil_SimpleDualBram_290_addra;
  wire                xil_SimpleDualBram_290_ena;
  wire       [13:0]   xil_SimpleDualBram_290_addrb;
  wire       [10:0]   xil_SimpleDualBram_291_addra;
  wire                xil_SimpleDualBram_291_ena;
  wire       [13:0]   xil_SimpleDualBram_291_addrb;
  wire       [10:0]   xil_SimpleDualBram_292_addra;
  wire                xil_SimpleDualBram_292_ena;
  wire       [13:0]   xil_SimpleDualBram_292_addrb;
  wire       [10:0]   xil_SimpleDualBram_293_addra;
  wire                xil_SimpleDualBram_293_ena;
  wire       [13:0]   xil_SimpleDualBram_293_addrb;
  wire       [10:0]   xil_SimpleDualBram_294_addra;
  wire                xil_SimpleDualBram_294_ena;
  wire       [13:0]   xil_SimpleDualBram_294_addrb;
  wire       [10:0]   xil_SimpleDualBram_295_addra;
  wire                xil_SimpleDualBram_295_ena;
  wire       [13:0]   xil_SimpleDualBram_295_addrb;
  wire       [10:0]   xil_SimpleDualBram_296_addra;
  wire                xil_SimpleDualBram_296_ena;
  wire       [13:0]   xil_SimpleDualBram_296_addrb;
  wire       [10:0]   xil_SimpleDualBram_297_addra;
  wire                xil_SimpleDualBram_297_ena;
  wire       [13:0]   xil_SimpleDualBram_297_addrb;
  wire       [10:0]   xil_SimpleDualBram_298_addra;
  wire                xil_SimpleDualBram_298_ena;
  wire       [13:0]   xil_SimpleDualBram_298_addrb;
  wire       [10:0]   xil_SimpleDualBram_299_addra;
  wire                xil_SimpleDualBram_299_ena;
  wire       [13:0]   xil_SimpleDualBram_299_addrb;
  wire       [10:0]   xil_SimpleDualBram_300_addra;
  wire                xil_SimpleDualBram_300_ena;
  wire       [13:0]   xil_SimpleDualBram_300_addrb;
  wire       [10:0]   xil_SimpleDualBram_301_addra;
  wire                xil_SimpleDualBram_301_ena;
  wire       [13:0]   xil_SimpleDualBram_301_addrb;
  wire       [10:0]   xil_SimpleDualBram_302_addra;
  wire                xil_SimpleDualBram_302_ena;
  wire       [13:0]   xil_SimpleDualBram_302_addrb;
  wire       [10:0]   xil_SimpleDualBram_303_addra;
  wire                xil_SimpleDualBram_303_ena;
  wire       [13:0]   xil_SimpleDualBram_303_addrb;
  wire       [10:0]   xil_SimpleDualBram_304_addra;
  wire                xil_SimpleDualBram_304_ena;
  wire       [13:0]   xil_SimpleDualBram_304_addrb;
  wire       [10:0]   xil_SimpleDualBram_305_addra;
  wire                xil_SimpleDualBram_305_ena;
  wire       [13:0]   xil_SimpleDualBram_305_addrb;
  wire       [10:0]   xil_SimpleDualBram_306_addra;
  wire                xil_SimpleDualBram_306_ena;
  wire       [13:0]   xil_SimpleDualBram_306_addrb;
  wire       [10:0]   xil_SimpleDualBram_307_addra;
  wire                xil_SimpleDualBram_307_ena;
  wire       [13:0]   xil_SimpleDualBram_307_addrb;
  wire       [10:0]   xil_SimpleDualBram_308_addra;
  wire                xil_SimpleDualBram_308_ena;
  wire       [13:0]   xil_SimpleDualBram_308_addrb;
  wire       [10:0]   xil_SimpleDualBram_309_addra;
  wire                xil_SimpleDualBram_309_ena;
  wire       [13:0]   xil_SimpleDualBram_309_addrb;
  wire       [10:0]   xil_SimpleDualBram_310_addra;
  wire                xil_SimpleDualBram_310_ena;
  wire       [13:0]   xil_SimpleDualBram_310_addrb;
  wire       [10:0]   xil_SimpleDualBram_311_addra;
  wire                xil_SimpleDualBram_311_ena;
  wire       [13:0]   xil_SimpleDualBram_311_addrb;
  wire       [10:0]   xil_SimpleDualBram_312_addra;
  wire                xil_SimpleDualBram_312_ena;
  wire       [13:0]   xil_SimpleDualBram_312_addrb;
  wire       [10:0]   xil_SimpleDualBram_313_addra;
  wire                xil_SimpleDualBram_313_ena;
  wire       [13:0]   xil_SimpleDualBram_313_addrb;
  wire       [10:0]   xil_SimpleDualBram_314_addra;
  wire                xil_SimpleDualBram_314_ena;
  wire       [13:0]   xil_SimpleDualBram_314_addrb;
  wire       [10:0]   xil_SimpleDualBram_315_addra;
  wire                xil_SimpleDualBram_315_ena;
  wire       [13:0]   xil_SimpleDualBram_315_addrb;
  wire       [10:0]   xil_SimpleDualBram_316_addra;
  wire                xil_SimpleDualBram_316_ena;
  wire       [13:0]   xil_SimpleDualBram_316_addrb;
  wire       [10:0]   xil_SimpleDualBram_317_addra;
  wire                xil_SimpleDualBram_317_ena;
  wire       [13:0]   xil_SimpleDualBram_317_addrb;
  wire       [10:0]   xil_SimpleDualBram_318_addra;
  wire                xil_SimpleDualBram_318_ena;
  wire       [13:0]   xil_SimpleDualBram_318_addrb;
  wire       [10:0]   xil_SimpleDualBram_319_addra;
  wire                xil_SimpleDualBram_319_ena;
  wire       [13:0]   xil_SimpleDualBram_319_addrb;
  wire       [10:0]   xil_SimpleDualBram_320_addra;
  wire                xil_SimpleDualBram_320_ena;
  wire       [13:0]   xil_SimpleDualBram_320_addrb;
  wire       [10:0]   xil_SimpleDualBram_321_addra;
  wire                xil_SimpleDualBram_321_ena;
  wire       [13:0]   xil_SimpleDualBram_321_addrb;
  wire       [10:0]   xil_SimpleDualBram_322_addra;
  wire                xil_SimpleDualBram_322_ena;
  wire       [13:0]   xil_SimpleDualBram_322_addrb;
  wire       [10:0]   xil_SimpleDualBram_323_addra;
  wire                xil_SimpleDualBram_323_ena;
  wire       [13:0]   xil_SimpleDualBram_323_addrb;
  wire       [10:0]   xil_SimpleDualBram_324_addra;
  wire                xil_SimpleDualBram_324_ena;
  wire       [13:0]   xil_SimpleDualBram_324_addrb;
  wire       [10:0]   xil_SimpleDualBram_325_addra;
  wire                xil_SimpleDualBram_325_ena;
  wire       [13:0]   xil_SimpleDualBram_325_addrb;
  wire       [10:0]   xil_SimpleDualBram_326_addra;
  wire                xil_SimpleDualBram_326_ena;
  wire       [13:0]   xil_SimpleDualBram_326_addrb;
  wire       [10:0]   xil_SimpleDualBram_327_addra;
  wire                xil_SimpleDualBram_327_ena;
  wire       [13:0]   xil_SimpleDualBram_327_addrb;
  wire       [10:0]   xil_SimpleDualBram_328_addra;
  wire                xil_SimpleDualBram_328_ena;
  wire       [13:0]   xil_SimpleDualBram_328_addrb;
  wire       [10:0]   xil_SimpleDualBram_329_addra;
  wire                xil_SimpleDualBram_329_ena;
  wire       [13:0]   xil_SimpleDualBram_329_addrb;
  wire       [10:0]   xil_SimpleDualBram_330_addra;
  wire                xil_SimpleDualBram_330_ena;
  wire       [13:0]   xil_SimpleDualBram_330_addrb;
  wire       [10:0]   xil_SimpleDualBram_331_addra;
  wire                xil_SimpleDualBram_331_ena;
  wire       [13:0]   xil_SimpleDualBram_331_addrb;
  wire       [10:0]   xil_SimpleDualBram_332_addra;
  wire                xil_SimpleDualBram_332_ena;
  wire       [13:0]   xil_SimpleDualBram_332_addrb;
  wire       [10:0]   xil_SimpleDualBram_333_addra;
  wire                xil_SimpleDualBram_333_ena;
  wire       [13:0]   xil_SimpleDualBram_333_addrb;
  wire       [10:0]   xil_SimpleDualBram_334_addra;
  wire                xil_SimpleDualBram_334_ena;
  wire       [13:0]   xil_SimpleDualBram_334_addrb;
  wire       [10:0]   xil_SimpleDualBram_335_addra;
  wire                xil_SimpleDualBram_335_ena;
  wire       [13:0]   xil_SimpleDualBram_335_addrb;
  wire       [10:0]   xil_SimpleDualBram_336_addra;
  wire                xil_SimpleDualBram_336_ena;
  wire       [13:0]   xil_SimpleDualBram_336_addrb;
  wire       [10:0]   xil_SimpleDualBram_337_addra;
  wire                xil_SimpleDualBram_337_ena;
  wire       [13:0]   xil_SimpleDualBram_337_addrb;
  wire       [10:0]   xil_SimpleDualBram_338_addra;
  wire                xil_SimpleDualBram_338_ena;
  wire       [13:0]   xil_SimpleDualBram_338_addrb;
  wire       [10:0]   xil_SimpleDualBram_339_addra;
  wire                xil_SimpleDualBram_339_ena;
  wire       [13:0]   xil_SimpleDualBram_339_addrb;
  wire       [10:0]   xil_SimpleDualBram_340_addra;
  wire                xil_SimpleDualBram_340_ena;
  wire       [13:0]   xil_SimpleDualBram_340_addrb;
  wire       [10:0]   xil_SimpleDualBram_341_addra;
  wire                xil_SimpleDualBram_341_ena;
  wire       [13:0]   xil_SimpleDualBram_341_addrb;
  wire       [10:0]   xil_SimpleDualBram_342_addra;
  wire                xil_SimpleDualBram_342_ena;
  wire       [13:0]   xil_SimpleDualBram_342_addrb;
  wire       [10:0]   xil_SimpleDualBram_343_addra;
  wire                xil_SimpleDualBram_343_ena;
  wire       [13:0]   xil_SimpleDualBram_343_addrb;
  wire       [10:0]   xil_SimpleDualBram_344_addra;
  wire                xil_SimpleDualBram_344_ena;
  wire       [13:0]   xil_SimpleDualBram_344_addrb;
  wire       [10:0]   xil_SimpleDualBram_345_addra;
  wire                xil_SimpleDualBram_345_ena;
  wire       [13:0]   xil_SimpleDualBram_345_addrb;
  wire       [10:0]   xil_SimpleDualBram_346_addra;
  wire                xil_SimpleDualBram_346_ena;
  wire       [13:0]   xil_SimpleDualBram_346_addrb;
  wire       [10:0]   xil_SimpleDualBram_347_addra;
  wire                xil_SimpleDualBram_347_ena;
  wire       [13:0]   xil_SimpleDualBram_347_addrb;
  wire       [10:0]   xil_SimpleDualBram_348_addra;
  wire                xil_SimpleDualBram_348_ena;
  wire       [13:0]   xil_SimpleDualBram_348_addrb;
  wire       [10:0]   xil_SimpleDualBram_349_addra;
  wire                xil_SimpleDualBram_349_ena;
  wire       [13:0]   xil_SimpleDualBram_349_addrb;
  wire       [10:0]   xil_SimpleDualBram_350_addra;
  wire                xil_SimpleDualBram_350_ena;
  wire       [13:0]   xil_SimpleDualBram_350_addrb;
  wire       [10:0]   xil_SimpleDualBram_351_addra;
  wire                xil_SimpleDualBram_351_ena;
  wire       [13:0]   xil_SimpleDualBram_351_addrb;
  wire       [10:0]   xil_SimpleDualBram_352_addra;
  wire                xil_SimpleDualBram_352_ena;
  wire       [13:0]   xil_SimpleDualBram_352_addrb;
  wire       [10:0]   xil_SimpleDualBram_353_addra;
  wire                xil_SimpleDualBram_353_ena;
  wire       [13:0]   xil_SimpleDualBram_353_addrb;
  wire       [10:0]   xil_SimpleDualBram_354_addra;
  wire                xil_SimpleDualBram_354_ena;
  wire       [13:0]   xil_SimpleDualBram_354_addrb;
  wire       [10:0]   xil_SimpleDualBram_355_addra;
  wire                xil_SimpleDualBram_355_ena;
  wire       [13:0]   xil_SimpleDualBram_355_addrb;
  wire       [10:0]   xil_SimpleDualBram_356_addra;
  wire                xil_SimpleDualBram_356_ena;
  wire       [13:0]   xil_SimpleDualBram_356_addrb;
  wire       [10:0]   xil_SimpleDualBram_357_addra;
  wire                xil_SimpleDualBram_357_ena;
  wire       [13:0]   xil_SimpleDualBram_357_addrb;
  wire       [10:0]   xil_SimpleDualBram_358_addra;
  wire                xil_SimpleDualBram_358_ena;
  wire       [13:0]   xil_SimpleDualBram_358_addrb;
  wire       [10:0]   xil_SimpleDualBram_359_addra;
  wire                xil_SimpleDualBram_359_ena;
  wire       [13:0]   xil_SimpleDualBram_359_addrb;
  wire       [10:0]   xil_SimpleDualBram_360_addra;
  wire                xil_SimpleDualBram_360_ena;
  wire       [13:0]   xil_SimpleDualBram_360_addrb;
  wire       [10:0]   xil_SimpleDualBram_361_addra;
  wire                xil_SimpleDualBram_361_ena;
  wire       [13:0]   xil_SimpleDualBram_361_addrb;
  wire       [10:0]   xil_SimpleDualBram_362_addra;
  wire                xil_SimpleDualBram_362_ena;
  wire       [13:0]   xil_SimpleDualBram_362_addrb;
  wire       [10:0]   xil_SimpleDualBram_363_addra;
  wire                xil_SimpleDualBram_363_ena;
  wire       [13:0]   xil_SimpleDualBram_363_addrb;
  wire       [10:0]   xil_SimpleDualBram_364_addra;
  wire                xil_SimpleDualBram_364_ena;
  wire       [13:0]   xil_SimpleDualBram_364_addrb;
  wire       [10:0]   xil_SimpleDualBram_365_addra;
  wire                xil_SimpleDualBram_365_ena;
  wire       [13:0]   xil_SimpleDualBram_365_addrb;
  wire       [10:0]   xil_SimpleDualBram_366_addra;
  wire                xil_SimpleDualBram_366_ena;
  wire       [13:0]   xil_SimpleDualBram_366_addrb;
  wire       [10:0]   xil_SimpleDualBram_367_addra;
  wire                xil_SimpleDualBram_367_ena;
  wire       [13:0]   xil_SimpleDualBram_367_addrb;
  wire       [10:0]   xil_SimpleDualBram_368_addra;
  wire                xil_SimpleDualBram_368_ena;
  wire       [13:0]   xil_SimpleDualBram_368_addrb;
  wire       [10:0]   xil_SimpleDualBram_369_addra;
  wire                xil_SimpleDualBram_369_ena;
  wire       [13:0]   xil_SimpleDualBram_369_addrb;
  wire       [10:0]   xil_SimpleDualBram_370_addra;
  wire                xil_SimpleDualBram_370_ena;
  wire       [13:0]   xil_SimpleDualBram_370_addrb;
  wire       [10:0]   xil_SimpleDualBram_371_addra;
  wire                xil_SimpleDualBram_371_ena;
  wire       [13:0]   xil_SimpleDualBram_371_addrb;
  wire       [10:0]   xil_SimpleDualBram_372_addra;
  wire                xil_SimpleDualBram_372_ena;
  wire       [13:0]   xil_SimpleDualBram_372_addrb;
  wire       [10:0]   xil_SimpleDualBram_373_addra;
  wire                xil_SimpleDualBram_373_ena;
  wire       [13:0]   xil_SimpleDualBram_373_addrb;
  wire       [10:0]   xil_SimpleDualBram_374_addra;
  wire                xil_SimpleDualBram_374_ena;
  wire       [13:0]   xil_SimpleDualBram_374_addrb;
  wire       [10:0]   xil_SimpleDualBram_375_addra;
  wire                xil_SimpleDualBram_375_ena;
  wire       [13:0]   xil_SimpleDualBram_375_addrb;
  wire       [10:0]   xil_SimpleDualBram_376_addra;
  wire                xil_SimpleDualBram_376_ena;
  wire       [13:0]   xil_SimpleDualBram_376_addrb;
  wire       [10:0]   xil_SimpleDualBram_377_addra;
  wire                xil_SimpleDualBram_377_ena;
  wire       [13:0]   xil_SimpleDualBram_377_addrb;
  wire       [10:0]   xil_SimpleDualBram_378_addra;
  wire                xil_SimpleDualBram_378_ena;
  wire       [13:0]   xil_SimpleDualBram_378_addrb;
  wire       [10:0]   xil_SimpleDualBram_379_addra;
  wire                xil_SimpleDualBram_379_ena;
  wire       [13:0]   xil_SimpleDualBram_379_addrb;
  wire       [10:0]   xil_SimpleDualBram_380_addra;
  wire                xil_SimpleDualBram_380_ena;
  wire       [13:0]   xil_SimpleDualBram_380_addrb;
  wire       [10:0]   xil_SimpleDualBram_381_addra;
  wire                xil_SimpleDualBram_381_ena;
  wire       [13:0]   xil_SimpleDualBram_381_addrb;
  wire       [10:0]   xil_SimpleDualBram_382_addra;
  wire                xil_SimpleDualBram_382_ena;
  wire       [13:0]   xil_SimpleDualBram_382_addrb;
  wire       [10:0]   xil_SimpleDualBram_383_addra;
  wire                xil_SimpleDualBram_383_ena;
  wire       [13:0]   xil_SimpleDualBram_383_addrb;
  wire       [10:0]   xil_SimpleDualBram_384_addra;
  wire                xil_SimpleDualBram_384_ena;
  wire       [13:0]   xil_SimpleDualBram_384_addrb;
  wire       [10:0]   xil_SimpleDualBram_385_addra;
  wire                xil_SimpleDualBram_385_ena;
  wire       [13:0]   xil_SimpleDualBram_385_addrb;
  wire       [10:0]   xil_SimpleDualBram_386_addra;
  wire                xil_SimpleDualBram_386_ena;
  wire       [13:0]   xil_SimpleDualBram_386_addrb;
  wire       [10:0]   xil_SimpleDualBram_387_addra;
  wire                xil_SimpleDualBram_387_ena;
  wire       [13:0]   xil_SimpleDualBram_387_addrb;
  wire       [10:0]   xil_SimpleDualBram_388_addra;
  wire                xil_SimpleDualBram_388_ena;
  wire       [13:0]   xil_SimpleDualBram_388_addrb;
  wire       [10:0]   xil_SimpleDualBram_389_addra;
  wire                xil_SimpleDualBram_389_ena;
  wire       [13:0]   xil_SimpleDualBram_389_addrb;
  wire       [10:0]   xil_SimpleDualBram_390_addra;
  wire                xil_SimpleDualBram_390_ena;
  wire       [13:0]   xil_SimpleDualBram_390_addrb;
  wire       [10:0]   xil_SimpleDualBram_391_addra;
  wire                xil_SimpleDualBram_391_ena;
  wire       [13:0]   xil_SimpleDualBram_391_addrb;
  wire       [10:0]   xil_SimpleDualBram_392_addra;
  wire                xil_SimpleDualBram_392_ena;
  wire       [13:0]   xil_SimpleDualBram_392_addrb;
  wire       [10:0]   xil_SimpleDualBram_393_addra;
  wire                xil_SimpleDualBram_393_ena;
  wire       [13:0]   xil_SimpleDualBram_393_addrb;
  wire       [10:0]   xil_SimpleDualBram_394_addra;
  wire                xil_SimpleDualBram_394_ena;
  wire       [13:0]   xil_SimpleDualBram_394_addrb;
  wire       [10:0]   xil_SimpleDualBram_395_addra;
  wire                xil_SimpleDualBram_395_ena;
  wire       [13:0]   xil_SimpleDualBram_395_addrb;
  wire       [10:0]   xil_SimpleDualBram_396_addra;
  wire                xil_SimpleDualBram_396_ena;
  wire       [13:0]   xil_SimpleDualBram_396_addrb;
  wire       [10:0]   xil_SimpleDualBram_397_addra;
  wire                xil_SimpleDualBram_397_ena;
  wire       [13:0]   xil_SimpleDualBram_397_addrb;
  wire       [10:0]   xil_SimpleDualBram_398_addra;
  wire                xil_SimpleDualBram_398_ena;
  wire       [13:0]   xil_SimpleDualBram_398_addrb;
  wire       [10:0]   xil_SimpleDualBram_399_addra;
  wire                xil_SimpleDualBram_399_ena;
  wire       [13:0]   xil_SimpleDualBram_399_addrb;
  wire       [10:0]   xil_SimpleDualBram_400_addra;
  wire                xil_SimpleDualBram_400_ena;
  wire       [13:0]   xil_SimpleDualBram_400_addrb;
  wire       [10:0]   xil_SimpleDualBram_401_addra;
  wire                xil_SimpleDualBram_401_ena;
  wire       [13:0]   xil_SimpleDualBram_401_addrb;
  wire       [10:0]   xil_SimpleDualBram_402_addra;
  wire                xil_SimpleDualBram_402_ena;
  wire       [13:0]   xil_SimpleDualBram_402_addrb;
  wire       [10:0]   xil_SimpleDualBram_403_addra;
  wire                xil_SimpleDualBram_403_ena;
  wire       [13:0]   xil_SimpleDualBram_403_addrb;
  wire       [10:0]   xil_SimpleDualBram_404_addra;
  wire                xil_SimpleDualBram_404_ena;
  wire       [13:0]   xil_SimpleDualBram_404_addrb;
  wire       [10:0]   xil_SimpleDualBram_405_addra;
  wire                xil_SimpleDualBram_405_ena;
  wire       [13:0]   xil_SimpleDualBram_405_addrb;
  wire       [10:0]   xil_SimpleDualBram_406_addra;
  wire                xil_SimpleDualBram_406_ena;
  wire       [13:0]   xil_SimpleDualBram_406_addrb;
  wire       [10:0]   xil_SimpleDualBram_407_addra;
  wire                xil_SimpleDualBram_407_ena;
  wire       [13:0]   xil_SimpleDualBram_407_addrb;
  wire       [10:0]   xil_SimpleDualBram_408_addra;
  wire                xil_SimpleDualBram_408_ena;
  wire       [13:0]   xil_SimpleDualBram_408_addrb;
  wire       [10:0]   xil_SimpleDualBram_409_addra;
  wire                xil_SimpleDualBram_409_ena;
  wire       [13:0]   xil_SimpleDualBram_409_addrb;
  wire       [10:0]   xil_SimpleDualBram_410_addra;
  wire                xil_SimpleDualBram_410_ena;
  wire       [13:0]   xil_SimpleDualBram_410_addrb;
  wire       [10:0]   xil_SimpleDualBram_411_addra;
  wire                xil_SimpleDualBram_411_ena;
  wire       [13:0]   xil_SimpleDualBram_411_addrb;
  wire       [10:0]   xil_SimpleDualBram_412_addra;
  wire                xil_SimpleDualBram_412_ena;
  wire       [13:0]   xil_SimpleDualBram_412_addrb;
  wire       [10:0]   xil_SimpleDualBram_413_addra;
  wire                xil_SimpleDualBram_413_ena;
  wire       [13:0]   xil_SimpleDualBram_413_addrb;
  wire       [10:0]   xil_SimpleDualBram_414_addra;
  wire                xil_SimpleDualBram_414_ena;
  wire       [13:0]   xil_SimpleDualBram_414_addrb;
  wire       [10:0]   xil_SimpleDualBram_415_addra;
  wire                xil_SimpleDualBram_415_ena;
  wire       [13:0]   xil_SimpleDualBram_415_addrb;
  wire       [10:0]   xil_SimpleDualBram_416_addra;
  wire                xil_SimpleDualBram_416_ena;
  wire       [13:0]   xil_SimpleDualBram_416_addrb;
  wire       [10:0]   xil_SimpleDualBram_417_addra;
  wire                xil_SimpleDualBram_417_ena;
  wire       [13:0]   xil_SimpleDualBram_417_addrb;
  wire       [10:0]   xil_SimpleDualBram_418_addra;
  wire                xil_SimpleDualBram_418_ena;
  wire       [13:0]   xil_SimpleDualBram_418_addrb;
  wire       [10:0]   xil_SimpleDualBram_419_addra;
  wire                xil_SimpleDualBram_419_ena;
  wire       [13:0]   xil_SimpleDualBram_419_addrb;
  wire       [10:0]   xil_SimpleDualBram_420_addra;
  wire                xil_SimpleDualBram_420_ena;
  wire       [13:0]   xil_SimpleDualBram_420_addrb;
  wire       [10:0]   xil_SimpleDualBram_421_addra;
  wire                xil_SimpleDualBram_421_ena;
  wire       [13:0]   xil_SimpleDualBram_421_addrb;
  wire       [10:0]   xil_SimpleDualBram_422_addra;
  wire                xil_SimpleDualBram_422_ena;
  wire       [13:0]   xil_SimpleDualBram_422_addrb;
  wire       [10:0]   xil_SimpleDualBram_423_addra;
  wire                xil_SimpleDualBram_423_ena;
  wire       [13:0]   xil_SimpleDualBram_423_addrb;
  wire       [10:0]   xil_SimpleDualBram_424_addra;
  wire                xil_SimpleDualBram_424_ena;
  wire       [13:0]   xil_SimpleDualBram_424_addrb;
  wire       [10:0]   xil_SimpleDualBram_425_addra;
  wire                xil_SimpleDualBram_425_ena;
  wire       [13:0]   xil_SimpleDualBram_425_addrb;
  wire       [10:0]   xil_SimpleDualBram_426_addra;
  wire                xil_SimpleDualBram_426_ena;
  wire       [13:0]   xil_SimpleDualBram_426_addrb;
  wire       [10:0]   xil_SimpleDualBram_427_addra;
  wire                xil_SimpleDualBram_427_ena;
  wire       [13:0]   xil_SimpleDualBram_427_addrb;
  wire       [10:0]   xil_SimpleDualBram_428_addra;
  wire                xil_SimpleDualBram_428_ena;
  wire       [13:0]   xil_SimpleDualBram_428_addrb;
  wire       [10:0]   xil_SimpleDualBram_429_addra;
  wire                xil_SimpleDualBram_429_ena;
  wire       [13:0]   xil_SimpleDualBram_429_addrb;
  wire       [10:0]   xil_SimpleDualBram_430_addra;
  wire                xil_SimpleDualBram_430_ena;
  wire       [13:0]   xil_SimpleDualBram_430_addrb;
  wire       [10:0]   xil_SimpleDualBram_431_addra;
  wire                xil_SimpleDualBram_431_ena;
  wire       [13:0]   xil_SimpleDualBram_431_addrb;
  wire       [10:0]   xil_SimpleDualBram_432_addra;
  wire                xil_SimpleDualBram_432_ena;
  wire       [13:0]   xil_SimpleDualBram_432_addrb;
  wire       [10:0]   xil_SimpleDualBram_433_addra;
  wire                xil_SimpleDualBram_433_ena;
  wire       [13:0]   xil_SimpleDualBram_433_addrb;
  wire       [10:0]   xil_SimpleDualBram_434_addra;
  wire                xil_SimpleDualBram_434_ena;
  wire       [13:0]   xil_SimpleDualBram_434_addrb;
  wire       [10:0]   xil_SimpleDualBram_435_addra;
  wire                xil_SimpleDualBram_435_ena;
  wire       [13:0]   xil_SimpleDualBram_435_addrb;
  wire       [10:0]   xil_SimpleDualBram_436_addra;
  wire                xil_SimpleDualBram_436_ena;
  wire       [13:0]   xil_SimpleDualBram_436_addrb;
  wire       [10:0]   xil_SimpleDualBram_437_addra;
  wire                xil_SimpleDualBram_437_ena;
  wire       [13:0]   xil_SimpleDualBram_437_addrb;
  wire       [10:0]   xil_SimpleDualBram_438_addra;
  wire                xil_SimpleDualBram_438_ena;
  wire       [13:0]   xil_SimpleDualBram_438_addrb;
  wire       [10:0]   xil_SimpleDualBram_439_addra;
  wire                xil_SimpleDualBram_439_ena;
  wire       [13:0]   xil_SimpleDualBram_439_addrb;
  wire       [10:0]   xil_SimpleDualBram_440_addra;
  wire                xil_SimpleDualBram_440_ena;
  wire       [13:0]   xil_SimpleDualBram_440_addrb;
  wire       [10:0]   xil_SimpleDualBram_441_addra;
  wire                xil_SimpleDualBram_441_ena;
  wire       [13:0]   xil_SimpleDualBram_441_addrb;
  wire       [10:0]   xil_SimpleDualBram_442_addra;
  wire                xil_SimpleDualBram_442_ena;
  wire       [13:0]   xil_SimpleDualBram_442_addrb;
  wire       [10:0]   xil_SimpleDualBram_443_addra;
  wire                xil_SimpleDualBram_443_ena;
  wire       [13:0]   xil_SimpleDualBram_443_addrb;
  wire       [10:0]   xil_SimpleDualBram_444_addra;
  wire                xil_SimpleDualBram_444_ena;
  wire       [13:0]   xil_SimpleDualBram_444_addrb;
  wire       [10:0]   xil_SimpleDualBram_445_addra;
  wire                xil_SimpleDualBram_445_ena;
  wire       [13:0]   xil_SimpleDualBram_445_addrb;
  wire       [10:0]   xil_SimpleDualBram_446_addra;
  wire                xil_SimpleDualBram_446_ena;
  wire       [13:0]   xil_SimpleDualBram_446_addrb;
  wire       [10:0]   xil_SimpleDualBram_447_addra;
  wire                xil_SimpleDualBram_447_ena;
  wire       [13:0]   xil_SimpleDualBram_447_addrb;
  wire       [10:0]   xil_SimpleDualBram_448_addra;
  wire                xil_SimpleDualBram_448_ena;
  wire       [13:0]   xil_SimpleDualBram_448_addrb;
  wire       [10:0]   xil_SimpleDualBram_449_addra;
  wire                xil_SimpleDualBram_449_ena;
  wire       [13:0]   xil_SimpleDualBram_449_addrb;
  wire       [10:0]   xil_SimpleDualBram_450_addra;
  wire                xil_SimpleDualBram_450_ena;
  wire       [13:0]   xil_SimpleDualBram_450_addrb;
  wire       [10:0]   xil_SimpleDualBram_451_addra;
  wire                xil_SimpleDualBram_451_ena;
  wire       [13:0]   xil_SimpleDualBram_451_addrb;
  wire       [10:0]   xil_SimpleDualBram_452_addra;
  wire                xil_SimpleDualBram_452_ena;
  wire       [13:0]   xil_SimpleDualBram_452_addrb;
  wire       [10:0]   xil_SimpleDualBram_453_addra;
  wire                xil_SimpleDualBram_453_ena;
  wire       [13:0]   xil_SimpleDualBram_453_addrb;
  wire       [10:0]   xil_SimpleDualBram_454_addra;
  wire                xil_SimpleDualBram_454_ena;
  wire       [13:0]   xil_SimpleDualBram_454_addrb;
  wire       [10:0]   xil_SimpleDualBram_455_addra;
  wire                xil_SimpleDualBram_455_ena;
  wire       [13:0]   xil_SimpleDualBram_455_addrb;
  wire       [10:0]   xil_SimpleDualBram_456_addra;
  wire                xil_SimpleDualBram_456_ena;
  wire       [13:0]   xil_SimpleDualBram_456_addrb;
  wire       [10:0]   xil_SimpleDualBram_457_addra;
  wire                xil_SimpleDualBram_457_ena;
  wire       [13:0]   xil_SimpleDualBram_457_addrb;
  wire       [10:0]   xil_SimpleDualBram_458_addra;
  wire                xil_SimpleDualBram_458_ena;
  wire       [13:0]   xil_SimpleDualBram_458_addrb;
  wire       [10:0]   xil_SimpleDualBram_459_addra;
  wire                xil_SimpleDualBram_459_ena;
  wire       [13:0]   xil_SimpleDualBram_459_addrb;
  wire       [10:0]   xil_SimpleDualBram_460_addra;
  wire                xil_SimpleDualBram_460_ena;
  wire       [13:0]   xil_SimpleDualBram_460_addrb;
  wire       [10:0]   xil_SimpleDualBram_461_addra;
  wire                xil_SimpleDualBram_461_ena;
  wire       [13:0]   xil_SimpleDualBram_461_addrb;
  wire       [10:0]   xil_SimpleDualBram_462_addra;
  wire                xil_SimpleDualBram_462_ena;
  wire       [13:0]   xil_SimpleDualBram_462_addrb;
  wire       [10:0]   xil_SimpleDualBram_463_addra;
  wire                xil_SimpleDualBram_463_ena;
  wire       [13:0]   xil_SimpleDualBram_463_addrb;
  wire       [10:0]   xil_SimpleDualBram_464_addra;
  wire                xil_SimpleDualBram_464_ena;
  wire       [13:0]   xil_SimpleDualBram_464_addrb;
  wire       [10:0]   xil_SimpleDualBram_465_addra;
  wire                xil_SimpleDualBram_465_ena;
  wire       [13:0]   xil_SimpleDualBram_465_addrb;
  wire       [10:0]   xil_SimpleDualBram_466_addra;
  wire                xil_SimpleDualBram_466_ena;
  wire       [13:0]   xil_SimpleDualBram_466_addrb;
  wire       [10:0]   xil_SimpleDualBram_467_addra;
  wire                xil_SimpleDualBram_467_ena;
  wire       [13:0]   xil_SimpleDualBram_467_addrb;
  wire       [10:0]   xil_SimpleDualBram_468_addra;
  wire                xil_SimpleDualBram_468_ena;
  wire       [13:0]   xil_SimpleDualBram_468_addrb;
  wire       [10:0]   xil_SimpleDualBram_469_addra;
  wire                xil_SimpleDualBram_469_ena;
  wire       [13:0]   xil_SimpleDualBram_469_addrb;
  wire       [10:0]   xil_SimpleDualBram_470_addra;
  wire                xil_SimpleDualBram_470_ena;
  wire       [13:0]   xil_SimpleDualBram_470_addrb;
  wire       [10:0]   xil_SimpleDualBram_471_addra;
  wire                xil_SimpleDualBram_471_ena;
  wire       [13:0]   xil_SimpleDualBram_471_addrb;
  wire       [10:0]   xil_SimpleDualBram_472_addra;
  wire                xil_SimpleDualBram_472_ena;
  wire       [13:0]   xil_SimpleDualBram_472_addrb;
  wire       [10:0]   xil_SimpleDualBram_473_addra;
  wire                xil_SimpleDualBram_473_ena;
  wire       [13:0]   xil_SimpleDualBram_473_addrb;
  wire       [10:0]   xil_SimpleDualBram_474_addra;
  wire                xil_SimpleDualBram_474_ena;
  wire       [13:0]   xil_SimpleDualBram_474_addrb;
  wire       [10:0]   xil_SimpleDualBram_475_addra;
  wire                xil_SimpleDualBram_475_ena;
  wire       [13:0]   xil_SimpleDualBram_475_addrb;
  wire       [10:0]   xil_SimpleDualBram_476_addra;
  wire                xil_SimpleDualBram_476_ena;
  wire       [13:0]   xil_SimpleDualBram_476_addrb;
  wire       [10:0]   xil_SimpleDualBram_477_addra;
  wire                xil_SimpleDualBram_477_ena;
  wire       [13:0]   xil_SimpleDualBram_477_addrb;
  wire       [10:0]   xil_SimpleDualBram_478_addra;
  wire                xil_SimpleDualBram_478_ena;
  wire       [13:0]   xil_SimpleDualBram_478_addrb;
  wire       [10:0]   xil_SimpleDualBram_479_addra;
  wire                xil_SimpleDualBram_479_ena;
  wire       [13:0]   xil_SimpleDualBram_479_addrb;
  wire       [10:0]   xil_SimpleDualBram_480_addra;
  wire                xil_SimpleDualBram_480_ena;
  wire       [13:0]   xil_SimpleDualBram_480_addrb;
  wire       [10:0]   xil_SimpleDualBram_481_addra;
  wire                xil_SimpleDualBram_481_ena;
  wire       [13:0]   xil_SimpleDualBram_481_addrb;
  wire       [10:0]   xil_SimpleDualBram_482_addra;
  wire                xil_SimpleDualBram_482_ena;
  wire       [13:0]   xil_SimpleDualBram_482_addrb;
  wire       [10:0]   xil_SimpleDualBram_483_addra;
  wire                xil_SimpleDualBram_483_ena;
  wire       [13:0]   xil_SimpleDualBram_483_addrb;
  wire       [10:0]   xil_SimpleDualBram_484_addra;
  wire                xil_SimpleDualBram_484_ena;
  wire       [13:0]   xil_SimpleDualBram_484_addrb;
  wire       [10:0]   xil_SimpleDualBram_485_addra;
  wire                xil_SimpleDualBram_485_ena;
  wire       [13:0]   xil_SimpleDualBram_485_addrb;
  wire       [10:0]   xil_SimpleDualBram_486_addra;
  wire                xil_SimpleDualBram_486_ena;
  wire       [13:0]   xil_SimpleDualBram_486_addrb;
  wire       [10:0]   xil_SimpleDualBram_487_addra;
  wire                xil_SimpleDualBram_487_ena;
  wire       [13:0]   xil_SimpleDualBram_487_addrb;
  wire       [10:0]   xil_SimpleDualBram_488_addra;
  wire                xil_SimpleDualBram_488_ena;
  wire       [13:0]   xil_SimpleDualBram_488_addrb;
  wire       [10:0]   xil_SimpleDualBram_489_addra;
  wire                xil_SimpleDualBram_489_ena;
  wire       [13:0]   xil_SimpleDualBram_489_addrb;
  wire       [10:0]   xil_SimpleDualBram_490_addra;
  wire                xil_SimpleDualBram_490_ena;
  wire       [13:0]   xil_SimpleDualBram_490_addrb;
  wire       [10:0]   xil_SimpleDualBram_491_addra;
  wire                xil_SimpleDualBram_491_ena;
  wire       [13:0]   xil_SimpleDualBram_491_addrb;
  wire       [10:0]   xil_SimpleDualBram_492_addra;
  wire                xil_SimpleDualBram_492_ena;
  wire       [13:0]   xil_SimpleDualBram_492_addrb;
  wire       [10:0]   xil_SimpleDualBram_493_addra;
  wire                xil_SimpleDualBram_493_ena;
  wire       [13:0]   xil_SimpleDualBram_493_addrb;
  wire       [10:0]   xil_SimpleDualBram_494_addra;
  wire                xil_SimpleDualBram_494_ena;
  wire       [13:0]   xil_SimpleDualBram_494_addrb;
  wire       [10:0]   xil_SimpleDualBram_495_addra;
  wire                xil_SimpleDualBram_495_ena;
  wire       [13:0]   xil_SimpleDualBram_495_addrb;
  wire       [10:0]   xil_SimpleDualBram_496_addra;
  wire                xil_SimpleDualBram_496_ena;
  wire       [13:0]   xil_SimpleDualBram_496_addrb;
  wire       [10:0]   xil_SimpleDualBram_497_addra;
  wire                xil_SimpleDualBram_497_ena;
  wire       [13:0]   xil_SimpleDualBram_497_addrb;
  wire       [10:0]   xil_SimpleDualBram_498_addra;
  wire                xil_SimpleDualBram_498_ena;
  wire       [13:0]   xil_SimpleDualBram_498_addrb;
  wire       [10:0]   xil_SimpleDualBram_499_addra;
  wire                xil_SimpleDualBram_499_ena;
  wire       [13:0]   xil_SimpleDualBram_499_addrb;
  wire       [10:0]   xil_SimpleDualBram_500_addra;
  wire                xil_SimpleDualBram_500_ena;
  wire       [13:0]   xil_SimpleDualBram_500_addrb;
  wire       [10:0]   xil_SimpleDualBram_501_addra;
  wire                xil_SimpleDualBram_501_ena;
  wire       [13:0]   xil_SimpleDualBram_501_addrb;
  wire       [10:0]   xil_SimpleDualBram_502_addra;
  wire                xil_SimpleDualBram_502_ena;
  wire       [13:0]   xil_SimpleDualBram_502_addrb;
  wire       [10:0]   xil_SimpleDualBram_503_addra;
  wire                xil_SimpleDualBram_503_ena;
  wire       [13:0]   xil_SimpleDualBram_503_addrb;
  wire       [10:0]   xil_SimpleDualBram_504_addra;
  wire                xil_SimpleDualBram_504_ena;
  wire       [13:0]   xil_SimpleDualBram_504_addrb;
  wire       [10:0]   xil_SimpleDualBram_505_addra;
  wire                xil_SimpleDualBram_505_ena;
  wire       [13:0]   xil_SimpleDualBram_505_addrb;
  wire       [10:0]   xil_SimpleDualBram_506_addra;
  wire                xil_SimpleDualBram_506_ena;
  wire       [13:0]   xil_SimpleDualBram_506_addrb;
  wire       [10:0]   xil_SimpleDualBram_507_addra;
  wire                xil_SimpleDualBram_507_ena;
  wire       [13:0]   xil_SimpleDualBram_507_addrb;
  wire       [10:0]   xil_SimpleDualBram_508_addra;
  wire                xil_SimpleDualBram_508_ena;
  wire       [13:0]   xil_SimpleDualBram_508_addrb;
  wire       [10:0]   xil_SimpleDualBram_509_addra;
  wire                xil_SimpleDualBram_509_ena;
  wire       [13:0]   xil_SimpleDualBram_509_addrb;
  wire       [10:0]   xil_SimpleDualBram_510_addra;
  wire                xil_SimpleDualBram_510_ena;
  wire       [13:0]   xil_SimpleDualBram_510_addrb;
  wire       [10:0]   xil_SimpleDualBram_511_addra;
  wire                xil_SimpleDualBram_511_ena;
  wire       [13:0]   xil_SimpleDualBram_511_addrb;
  wire       [7:0]    xil_SimpleDualBram_doutb;
  wire       [7:0]    xil_SimpleDualBram_1_doutb;
  wire       [7:0]    xil_SimpleDualBram_2_doutb;
  wire       [7:0]    xil_SimpleDualBram_3_doutb;
  wire       [7:0]    xil_SimpleDualBram_4_doutb;
  wire       [7:0]    xil_SimpleDualBram_5_doutb;
  wire       [7:0]    xil_SimpleDualBram_6_doutb;
  wire       [7:0]    xil_SimpleDualBram_7_doutb;
  wire       [7:0]    xil_SimpleDualBram_8_doutb;
  wire       [7:0]    xil_SimpleDualBram_9_doutb;
  wire       [7:0]    xil_SimpleDualBram_10_doutb;
  wire       [7:0]    xil_SimpleDualBram_11_doutb;
  wire       [7:0]    xil_SimpleDualBram_12_doutb;
  wire       [7:0]    xil_SimpleDualBram_13_doutb;
  wire       [7:0]    xil_SimpleDualBram_14_doutb;
  wire       [7:0]    xil_SimpleDualBram_15_doutb;
  wire       [7:0]    xil_SimpleDualBram_16_doutb;
  wire       [7:0]    xil_SimpleDualBram_17_doutb;
  wire       [7:0]    xil_SimpleDualBram_18_doutb;
  wire       [7:0]    xil_SimpleDualBram_19_doutb;
  wire       [7:0]    xil_SimpleDualBram_20_doutb;
  wire       [7:0]    xil_SimpleDualBram_21_doutb;
  wire       [7:0]    xil_SimpleDualBram_22_doutb;
  wire       [7:0]    xil_SimpleDualBram_23_doutb;
  wire       [7:0]    xil_SimpleDualBram_24_doutb;
  wire       [7:0]    xil_SimpleDualBram_25_doutb;
  wire       [7:0]    xil_SimpleDualBram_26_doutb;
  wire       [7:0]    xil_SimpleDualBram_27_doutb;
  wire       [7:0]    xil_SimpleDualBram_28_doutb;
  wire       [7:0]    xil_SimpleDualBram_29_doutb;
  wire       [7:0]    xil_SimpleDualBram_30_doutb;
  wire       [7:0]    xil_SimpleDualBram_31_doutb;
  wire       [7:0]    xil_SimpleDualBram_32_doutb;
  wire       [7:0]    xil_SimpleDualBram_33_doutb;
  wire       [7:0]    xil_SimpleDualBram_34_doutb;
  wire       [7:0]    xil_SimpleDualBram_35_doutb;
  wire       [7:0]    xil_SimpleDualBram_36_doutb;
  wire       [7:0]    xil_SimpleDualBram_37_doutb;
  wire       [7:0]    xil_SimpleDualBram_38_doutb;
  wire       [7:0]    xil_SimpleDualBram_39_doutb;
  wire       [7:0]    xil_SimpleDualBram_40_doutb;
  wire       [7:0]    xil_SimpleDualBram_41_doutb;
  wire       [7:0]    xil_SimpleDualBram_42_doutb;
  wire       [7:0]    xil_SimpleDualBram_43_doutb;
  wire       [7:0]    xil_SimpleDualBram_44_doutb;
  wire       [7:0]    xil_SimpleDualBram_45_doutb;
  wire       [7:0]    xil_SimpleDualBram_46_doutb;
  wire       [7:0]    xil_SimpleDualBram_47_doutb;
  wire       [7:0]    xil_SimpleDualBram_48_doutb;
  wire       [7:0]    xil_SimpleDualBram_49_doutb;
  wire       [7:0]    xil_SimpleDualBram_50_doutb;
  wire       [7:0]    xil_SimpleDualBram_51_doutb;
  wire       [7:0]    xil_SimpleDualBram_52_doutb;
  wire       [7:0]    xil_SimpleDualBram_53_doutb;
  wire       [7:0]    xil_SimpleDualBram_54_doutb;
  wire       [7:0]    xil_SimpleDualBram_55_doutb;
  wire       [7:0]    xil_SimpleDualBram_56_doutb;
  wire       [7:0]    xil_SimpleDualBram_57_doutb;
  wire       [7:0]    xil_SimpleDualBram_58_doutb;
  wire       [7:0]    xil_SimpleDualBram_59_doutb;
  wire       [7:0]    xil_SimpleDualBram_60_doutb;
  wire       [7:0]    xil_SimpleDualBram_61_doutb;
  wire       [7:0]    xil_SimpleDualBram_62_doutb;
  wire       [7:0]    xil_SimpleDualBram_63_doutb;
  wire       [7:0]    xil_SimpleDualBram_64_doutb;
  wire       [7:0]    xil_SimpleDualBram_65_doutb;
  wire       [7:0]    xil_SimpleDualBram_66_doutb;
  wire       [7:0]    xil_SimpleDualBram_67_doutb;
  wire       [7:0]    xil_SimpleDualBram_68_doutb;
  wire       [7:0]    xil_SimpleDualBram_69_doutb;
  wire       [7:0]    xil_SimpleDualBram_70_doutb;
  wire       [7:0]    xil_SimpleDualBram_71_doutb;
  wire       [7:0]    xil_SimpleDualBram_72_doutb;
  wire       [7:0]    xil_SimpleDualBram_73_doutb;
  wire       [7:0]    xil_SimpleDualBram_74_doutb;
  wire       [7:0]    xil_SimpleDualBram_75_doutb;
  wire       [7:0]    xil_SimpleDualBram_76_doutb;
  wire       [7:0]    xil_SimpleDualBram_77_doutb;
  wire       [7:0]    xil_SimpleDualBram_78_doutb;
  wire       [7:0]    xil_SimpleDualBram_79_doutb;
  wire       [7:0]    xil_SimpleDualBram_80_doutb;
  wire       [7:0]    xil_SimpleDualBram_81_doutb;
  wire       [7:0]    xil_SimpleDualBram_82_doutb;
  wire       [7:0]    xil_SimpleDualBram_83_doutb;
  wire       [7:0]    xil_SimpleDualBram_84_doutb;
  wire       [7:0]    xil_SimpleDualBram_85_doutb;
  wire       [7:0]    xil_SimpleDualBram_86_doutb;
  wire       [7:0]    xil_SimpleDualBram_87_doutb;
  wire       [7:0]    xil_SimpleDualBram_88_doutb;
  wire       [7:0]    xil_SimpleDualBram_89_doutb;
  wire       [7:0]    xil_SimpleDualBram_90_doutb;
  wire       [7:0]    xil_SimpleDualBram_91_doutb;
  wire       [7:0]    xil_SimpleDualBram_92_doutb;
  wire       [7:0]    xil_SimpleDualBram_93_doutb;
  wire       [7:0]    xil_SimpleDualBram_94_doutb;
  wire       [7:0]    xil_SimpleDualBram_95_doutb;
  wire       [7:0]    xil_SimpleDualBram_96_doutb;
  wire       [7:0]    xil_SimpleDualBram_97_doutb;
  wire       [7:0]    xil_SimpleDualBram_98_doutb;
  wire       [7:0]    xil_SimpleDualBram_99_doutb;
  wire       [7:0]    xil_SimpleDualBram_100_doutb;
  wire       [7:0]    xil_SimpleDualBram_101_doutb;
  wire       [7:0]    xil_SimpleDualBram_102_doutb;
  wire       [7:0]    xil_SimpleDualBram_103_doutb;
  wire       [7:0]    xil_SimpleDualBram_104_doutb;
  wire       [7:0]    xil_SimpleDualBram_105_doutb;
  wire       [7:0]    xil_SimpleDualBram_106_doutb;
  wire       [7:0]    xil_SimpleDualBram_107_doutb;
  wire       [7:0]    xil_SimpleDualBram_108_doutb;
  wire       [7:0]    xil_SimpleDualBram_109_doutb;
  wire       [7:0]    xil_SimpleDualBram_110_doutb;
  wire       [7:0]    xil_SimpleDualBram_111_doutb;
  wire       [7:0]    xil_SimpleDualBram_112_doutb;
  wire       [7:0]    xil_SimpleDualBram_113_doutb;
  wire       [7:0]    xil_SimpleDualBram_114_doutb;
  wire       [7:0]    xil_SimpleDualBram_115_doutb;
  wire       [7:0]    xil_SimpleDualBram_116_doutb;
  wire       [7:0]    xil_SimpleDualBram_117_doutb;
  wire       [7:0]    xil_SimpleDualBram_118_doutb;
  wire       [7:0]    xil_SimpleDualBram_119_doutb;
  wire       [7:0]    xil_SimpleDualBram_120_doutb;
  wire       [7:0]    xil_SimpleDualBram_121_doutb;
  wire       [7:0]    xil_SimpleDualBram_122_doutb;
  wire       [7:0]    xil_SimpleDualBram_123_doutb;
  wire       [7:0]    xil_SimpleDualBram_124_doutb;
  wire       [7:0]    xil_SimpleDualBram_125_doutb;
  wire       [7:0]    xil_SimpleDualBram_126_doutb;
  wire       [7:0]    xil_SimpleDualBram_127_doutb;
  wire       [7:0]    xil_SimpleDualBram_128_doutb;
  wire       [7:0]    xil_SimpleDualBram_129_doutb;
  wire       [7:0]    xil_SimpleDualBram_130_doutb;
  wire       [7:0]    xil_SimpleDualBram_131_doutb;
  wire       [7:0]    xil_SimpleDualBram_132_doutb;
  wire       [7:0]    xil_SimpleDualBram_133_doutb;
  wire       [7:0]    xil_SimpleDualBram_134_doutb;
  wire       [7:0]    xil_SimpleDualBram_135_doutb;
  wire       [7:0]    xil_SimpleDualBram_136_doutb;
  wire       [7:0]    xil_SimpleDualBram_137_doutb;
  wire       [7:0]    xil_SimpleDualBram_138_doutb;
  wire       [7:0]    xil_SimpleDualBram_139_doutb;
  wire       [7:0]    xil_SimpleDualBram_140_doutb;
  wire       [7:0]    xil_SimpleDualBram_141_doutb;
  wire       [7:0]    xil_SimpleDualBram_142_doutb;
  wire       [7:0]    xil_SimpleDualBram_143_doutb;
  wire       [7:0]    xil_SimpleDualBram_144_doutb;
  wire       [7:0]    xil_SimpleDualBram_145_doutb;
  wire       [7:0]    xil_SimpleDualBram_146_doutb;
  wire       [7:0]    xil_SimpleDualBram_147_doutb;
  wire       [7:0]    xil_SimpleDualBram_148_doutb;
  wire       [7:0]    xil_SimpleDualBram_149_doutb;
  wire       [7:0]    xil_SimpleDualBram_150_doutb;
  wire       [7:0]    xil_SimpleDualBram_151_doutb;
  wire       [7:0]    xil_SimpleDualBram_152_doutb;
  wire       [7:0]    xil_SimpleDualBram_153_doutb;
  wire       [7:0]    xil_SimpleDualBram_154_doutb;
  wire       [7:0]    xil_SimpleDualBram_155_doutb;
  wire       [7:0]    xil_SimpleDualBram_156_doutb;
  wire       [7:0]    xil_SimpleDualBram_157_doutb;
  wire       [7:0]    xil_SimpleDualBram_158_doutb;
  wire       [7:0]    xil_SimpleDualBram_159_doutb;
  wire       [7:0]    xil_SimpleDualBram_160_doutb;
  wire       [7:0]    xil_SimpleDualBram_161_doutb;
  wire       [7:0]    xil_SimpleDualBram_162_doutb;
  wire       [7:0]    xil_SimpleDualBram_163_doutb;
  wire       [7:0]    xil_SimpleDualBram_164_doutb;
  wire       [7:0]    xil_SimpleDualBram_165_doutb;
  wire       [7:0]    xil_SimpleDualBram_166_doutb;
  wire       [7:0]    xil_SimpleDualBram_167_doutb;
  wire       [7:0]    xil_SimpleDualBram_168_doutb;
  wire       [7:0]    xil_SimpleDualBram_169_doutb;
  wire       [7:0]    xil_SimpleDualBram_170_doutb;
  wire       [7:0]    xil_SimpleDualBram_171_doutb;
  wire       [7:0]    xil_SimpleDualBram_172_doutb;
  wire       [7:0]    xil_SimpleDualBram_173_doutb;
  wire       [7:0]    xil_SimpleDualBram_174_doutb;
  wire       [7:0]    xil_SimpleDualBram_175_doutb;
  wire       [7:0]    xil_SimpleDualBram_176_doutb;
  wire       [7:0]    xil_SimpleDualBram_177_doutb;
  wire       [7:0]    xil_SimpleDualBram_178_doutb;
  wire       [7:0]    xil_SimpleDualBram_179_doutb;
  wire       [7:0]    xil_SimpleDualBram_180_doutb;
  wire       [7:0]    xil_SimpleDualBram_181_doutb;
  wire       [7:0]    xil_SimpleDualBram_182_doutb;
  wire       [7:0]    xil_SimpleDualBram_183_doutb;
  wire       [7:0]    xil_SimpleDualBram_184_doutb;
  wire       [7:0]    xil_SimpleDualBram_185_doutb;
  wire       [7:0]    xil_SimpleDualBram_186_doutb;
  wire       [7:0]    xil_SimpleDualBram_187_doutb;
  wire       [7:0]    xil_SimpleDualBram_188_doutb;
  wire       [7:0]    xil_SimpleDualBram_189_doutb;
  wire       [7:0]    xil_SimpleDualBram_190_doutb;
  wire       [7:0]    xil_SimpleDualBram_191_doutb;
  wire       [7:0]    xil_SimpleDualBram_192_doutb;
  wire       [7:0]    xil_SimpleDualBram_193_doutb;
  wire       [7:0]    xil_SimpleDualBram_194_doutb;
  wire       [7:0]    xil_SimpleDualBram_195_doutb;
  wire       [7:0]    xil_SimpleDualBram_196_doutb;
  wire       [7:0]    xil_SimpleDualBram_197_doutb;
  wire       [7:0]    xil_SimpleDualBram_198_doutb;
  wire       [7:0]    xil_SimpleDualBram_199_doutb;
  wire       [7:0]    xil_SimpleDualBram_200_doutb;
  wire       [7:0]    xil_SimpleDualBram_201_doutb;
  wire       [7:0]    xil_SimpleDualBram_202_doutb;
  wire       [7:0]    xil_SimpleDualBram_203_doutb;
  wire       [7:0]    xil_SimpleDualBram_204_doutb;
  wire       [7:0]    xil_SimpleDualBram_205_doutb;
  wire       [7:0]    xil_SimpleDualBram_206_doutb;
  wire       [7:0]    xil_SimpleDualBram_207_doutb;
  wire       [7:0]    xil_SimpleDualBram_208_doutb;
  wire       [7:0]    xil_SimpleDualBram_209_doutb;
  wire       [7:0]    xil_SimpleDualBram_210_doutb;
  wire       [7:0]    xil_SimpleDualBram_211_doutb;
  wire       [7:0]    xil_SimpleDualBram_212_doutb;
  wire       [7:0]    xil_SimpleDualBram_213_doutb;
  wire       [7:0]    xil_SimpleDualBram_214_doutb;
  wire       [7:0]    xil_SimpleDualBram_215_doutb;
  wire       [7:0]    xil_SimpleDualBram_216_doutb;
  wire       [7:0]    xil_SimpleDualBram_217_doutb;
  wire       [7:0]    xil_SimpleDualBram_218_doutb;
  wire       [7:0]    xil_SimpleDualBram_219_doutb;
  wire       [7:0]    xil_SimpleDualBram_220_doutb;
  wire       [7:0]    xil_SimpleDualBram_221_doutb;
  wire       [7:0]    xil_SimpleDualBram_222_doutb;
  wire       [7:0]    xil_SimpleDualBram_223_doutb;
  wire       [7:0]    xil_SimpleDualBram_224_doutb;
  wire       [7:0]    xil_SimpleDualBram_225_doutb;
  wire       [7:0]    xil_SimpleDualBram_226_doutb;
  wire       [7:0]    xil_SimpleDualBram_227_doutb;
  wire       [7:0]    xil_SimpleDualBram_228_doutb;
  wire       [7:0]    xil_SimpleDualBram_229_doutb;
  wire       [7:0]    xil_SimpleDualBram_230_doutb;
  wire       [7:0]    xil_SimpleDualBram_231_doutb;
  wire       [7:0]    xil_SimpleDualBram_232_doutb;
  wire       [7:0]    xil_SimpleDualBram_233_doutb;
  wire       [7:0]    xil_SimpleDualBram_234_doutb;
  wire       [7:0]    xil_SimpleDualBram_235_doutb;
  wire       [7:0]    xil_SimpleDualBram_236_doutb;
  wire       [7:0]    xil_SimpleDualBram_237_doutb;
  wire       [7:0]    xil_SimpleDualBram_238_doutb;
  wire       [7:0]    xil_SimpleDualBram_239_doutb;
  wire       [7:0]    xil_SimpleDualBram_240_doutb;
  wire       [7:0]    xil_SimpleDualBram_241_doutb;
  wire       [7:0]    xil_SimpleDualBram_242_doutb;
  wire       [7:0]    xil_SimpleDualBram_243_doutb;
  wire       [7:0]    xil_SimpleDualBram_244_doutb;
  wire       [7:0]    xil_SimpleDualBram_245_doutb;
  wire       [7:0]    xil_SimpleDualBram_246_doutb;
  wire       [7:0]    xil_SimpleDualBram_247_doutb;
  wire       [7:0]    xil_SimpleDualBram_248_doutb;
  wire       [7:0]    xil_SimpleDualBram_249_doutb;
  wire       [7:0]    xil_SimpleDualBram_250_doutb;
  wire       [7:0]    xil_SimpleDualBram_251_doutb;
  wire       [7:0]    xil_SimpleDualBram_252_doutb;
  wire       [7:0]    xil_SimpleDualBram_253_doutb;
  wire       [7:0]    xil_SimpleDualBram_254_doutb;
  wire       [7:0]    xil_SimpleDualBram_255_doutb;
  wire       [7:0]    xil_SimpleDualBram_256_doutb;
  wire       [7:0]    xil_SimpleDualBram_257_doutb;
  wire       [7:0]    xil_SimpleDualBram_258_doutb;
  wire       [7:0]    xil_SimpleDualBram_259_doutb;
  wire       [7:0]    xil_SimpleDualBram_260_doutb;
  wire       [7:0]    xil_SimpleDualBram_261_doutb;
  wire       [7:0]    xil_SimpleDualBram_262_doutb;
  wire       [7:0]    xil_SimpleDualBram_263_doutb;
  wire       [7:0]    xil_SimpleDualBram_264_doutb;
  wire       [7:0]    xil_SimpleDualBram_265_doutb;
  wire       [7:0]    xil_SimpleDualBram_266_doutb;
  wire       [7:0]    xil_SimpleDualBram_267_doutb;
  wire       [7:0]    xil_SimpleDualBram_268_doutb;
  wire       [7:0]    xil_SimpleDualBram_269_doutb;
  wire       [7:0]    xil_SimpleDualBram_270_doutb;
  wire       [7:0]    xil_SimpleDualBram_271_doutb;
  wire       [7:0]    xil_SimpleDualBram_272_doutb;
  wire       [7:0]    xil_SimpleDualBram_273_doutb;
  wire       [7:0]    xil_SimpleDualBram_274_doutb;
  wire       [7:0]    xil_SimpleDualBram_275_doutb;
  wire       [7:0]    xil_SimpleDualBram_276_doutb;
  wire       [7:0]    xil_SimpleDualBram_277_doutb;
  wire       [7:0]    xil_SimpleDualBram_278_doutb;
  wire       [7:0]    xil_SimpleDualBram_279_doutb;
  wire       [7:0]    xil_SimpleDualBram_280_doutb;
  wire       [7:0]    xil_SimpleDualBram_281_doutb;
  wire       [7:0]    xil_SimpleDualBram_282_doutb;
  wire       [7:0]    xil_SimpleDualBram_283_doutb;
  wire       [7:0]    xil_SimpleDualBram_284_doutb;
  wire       [7:0]    xil_SimpleDualBram_285_doutb;
  wire       [7:0]    xil_SimpleDualBram_286_doutb;
  wire       [7:0]    xil_SimpleDualBram_287_doutb;
  wire       [7:0]    xil_SimpleDualBram_288_doutb;
  wire       [7:0]    xil_SimpleDualBram_289_doutb;
  wire       [7:0]    xil_SimpleDualBram_290_doutb;
  wire       [7:0]    xil_SimpleDualBram_291_doutb;
  wire       [7:0]    xil_SimpleDualBram_292_doutb;
  wire       [7:0]    xil_SimpleDualBram_293_doutb;
  wire       [7:0]    xil_SimpleDualBram_294_doutb;
  wire       [7:0]    xil_SimpleDualBram_295_doutb;
  wire       [7:0]    xil_SimpleDualBram_296_doutb;
  wire       [7:0]    xil_SimpleDualBram_297_doutb;
  wire       [7:0]    xil_SimpleDualBram_298_doutb;
  wire       [7:0]    xil_SimpleDualBram_299_doutb;
  wire       [7:0]    xil_SimpleDualBram_300_doutb;
  wire       [7:0]    xil_SimpleDualBram_301_doutb;
  wire       [7:0]    xil_SimpleDualBram_302_doutb;
  wire       [7:0]    xil_SimpleDualBram_303_doutb;
  wire       [7:0]    xil_SimpleDualBram_304_doutb;
  wire       [7:0]    xil_SimpleDualBram_305_doutb;
  wire       [7:0]    xil_SimpleDualBram_306_doutb;
  wire       [7:0]    xil_SimpleDualBram_307_doutb;
  wire       [7:0]    xil_SimpleDualBram_308_doutb;
  wire       [7:0]    xil_SimpleDualBram_309_doutb;
  wire       [7:0]    xil_SimpleDualBram_310_doutb;
  wire       [7:0]    xil_SimpleDualBram_311_doutb;
  wire       [7:0]    xil_SimpleDualBram_312_doutb;
  wire       [7:0]    xil_SimpleDualBram_313_doutb;
  wire       [7:0]    xil_SimpleDualBram_314_doutb;
  wire       [7:0]    xil_SimpleDualBram_315_doutb;
  wire       [7:0]    xil_SimpleDualBram_316_doutb;
  wire       [7:0]    xil_SimpleDualBram_317_doutb;
  wire       [7:0]    xil_SimpleDualBram_318_doutb;
  wire       [7:0]    xil_SimpleDualBram_319_doutb;
  wire       [7:0]    xil_SimpleDualBram_320_doutb;
  wire       [7:0]    xil_SimpleDualBram_321_doutb;
  wire       [7:0]    xil_SimpleDualBram_322_doutb;
  wire       [7:0]    xil_SimpleDualBram_323_doutb;
  wire       [7:0]    xil_SimpleDualBram_324_doutb;
  wire       [7:0]    xil_SimpleDualBram_325_doutb;
  wire       [7:0]    xil_SimpleDualBram_326_doutb;
  wire       [7:0]    xil_SimpleDualBram_327_doutb;
  wire       [7:0]    xil_SimpleDualBram_328_doutb;
  wire       [7:0]    xil_SimpleDualBram_329_doutb;
  wire       [7:0]    xil_SimpleDualBram_330_doutb;
  wire       [7:0]    xil_SimpleDualBram_331_doutb;
  wire       [7:0]    xil_SimpleDualBram_332_doutb;
  wire       [7:0]    xil_SimpleDualBram_333_doutb;
  wire       [7:0]    xil_SimpleDualBram_334_doutb;
  wire       [7:0]    xil_SimpleDualBram_335_doutb;
  wire       [7:0]    xil_SimpleDualBram_336_doutb;
  wire       [7:0]    xil_SimpleDualBram_337_doutb;
  wire       [7:0]    xil_SimpleDualBram_338_doutb;
  wire       [7:0]    xil_SimpleDualBram_339_doutb;
  wire       [7:0]    xil_SimpleDualBram_340_doutb;
  wire       [7:0]    xil_SimpleDualBram_341_doutb;
  wire       [7:0]    xil_SimpleDualBram_342_doutb;
  wire       [7:0]    xil_SimpleDualBram_343_doutb;
  wire       [7:0]    xil_SimpleDualBram_344_doutb;
  wire       [7:0]    xil_SimpleDualBram_345_doutb;
  wire       [7:0]    xil_SimpleDualBram_346_doutb;
  wire       [7:0]    xil_SimpleDualBram_347_doutb;
  wire       [7:0]    xil_SimpleDualBram_348_doutb;
  wire       [7:0]    xil_SimpleDualBram_349_doutb;
  wire       [7:0]    xil_SimpleDualBram_350_doutb;
  wire       [7:0]    xil_SimpleDualBram_351_doutb;
  wire       [7:0]    xil_SimpleDualBram_352_doutb;
  wire       [7:0]    xil_SimpleDualBram_353_doutb;
  wire       [7:0]    xil_SimpleDualBram_354_doutb;
  wire       [7:0]    xil_SimpleDualBram_355_doutb;
  wire       [7:0]    xil_SimpleDualBram_356_doutb;
  wire       [7:0]    xil_SimpleDualBram_357_doutb;
  wire       [7:0]    xil_SimpleDualBram_358_doutb;
  wire       [7:0]    xil_SimpleDualBram_359_doutb;
  wire       [7:0]    xil_SimpleDualBram_360_doutb;
  wire       [7:0]    xil_SimpleDualBram_361_doutb;
  wire       [7:0]    xil_SimpleDualBram_362_doutb;
  wire       [7:0]    xil_SimpleDualBram_363_doutb;
  wire       [7:0]    xil_SimpleDualBram_364_doutb;
  wire       [7:0]    xil_SimpleDualBram_365_doutb;
  wire       [7:0]    xil_SimpleDualBram_366_doutb;
  wire       [7:0]    xil_SimpleDualBram_367_doutb;
  wire       [7:0]    xil_SimpleDualBram_368_doutb;
  wire       [7:0]    xil_SimpleDualBram_369_doutb;
  wire       [7:0]    xil_SimpleDualBram_370_doutb;
  wire       [7:0]    xil_SimpleDualBram_371_doutb;
  wire       [7:0]    xil_SimpleDualBram_372_doutb;
  wire       [7:0]    xil_SimpleDualBram_373_doutb;
  wire       [7:0]    xil_SimpleDualBram_374_doutb;
  wire       [7:0]    xil_SimpleDualBram_375_doutb;
  wire       [7:0]    xil_SimpleDualBram_376_doutb;
  wire       [7:0]    xil_SimpleDualBram_377_doutb;
  wire       [7:0]    xil_SimpleDualBram_378_doutb;
  wire       [7:0]    xil_SimpleDualBram_379_doutb;
  wire       [7:0]    xil_SimpleDualBram_380_doutb;
  wire       [7:0]    xil_SimpleDualBram_381_doutb;
  wire       [7:0]    xil_SimpleDualBram_382_doutb;
  wire       [7:0]    xil_SimpleDualBram_383_doutb;
  wire       [7:0]    xil_SimpleDualBram_384_doutb;
  wire       [7:0]    xil_SimpleDualBram_385_doutb;
  wire       [7:0]    xil_SimpleDualBram_386_doutb;
  wire       [7:0]    xil_SimpleDualBram_387_doutb;
  wire       [7:0]    xil_SimpleDualBram_388_doutb;
  wire       [7:0]    xil_SimpleDualBram_389_doutb;
  wire       [7:0]    xil_SimpleDualBram_390_doutb;
  wire       [7:0]    xil_SimpleDualBram_391_doutb;
  wire       [7:0]    xil_SimpleDualBram_392_doutb;
  wire       [7:0]    xil_SimpleDualBram_393_doutb;
  wire       [7:0]    xil_SimpleDualBram_394_doutb;
  wire       [7:0]    xil_SimpleDualBram_395_doutb;
  wire       [7:0]    xil_SimpleDualBram_396_doutb;
  wire       [7:0]    xil_SimpleDualBram_397_doutb;
  wire       [7:0]    xil_SimpleDualBram_398_doutb;
  wire       [7:0]    xil_SimpleDualBram_399_doutb;
  wire       [7:0]    xil_SimpleDualBram_400_doutb;
  wire       [7:0]    xil_SimpleDualBram_401_doutb;
  wire       [7:0]    xil_SimpleDualBram_402_doutb;
  wire       [7:0]    xil_SimpleDualBram_403_doutb;
  wire       [7:0]    xil_SimpleDualBram_404_doutb;
  wire       [7:0]    xil_SimpleDualBram_405_doutb;
  wire       [7:0]    xil_SimpleDualBram_406_doutb;
  wire       [7:0]    xil_SimpleDualBram_407_doutb;
  wire       [7:0]    xil_SimpleDualBram_408_doutb;
  wire       [7:0]    xil_SimpleDualBram_409_doutb;
  wire       [7:0]    xil_SimpleDualBram_410_doutb;
  wire       [7:0]    xil_SimpleDualBram_411_doutb;
  wire       [7:0]    xil_SimpleDualBram_412_doutb;
  wire       [7:0]    xil_SimpleDualBram_413_doutb;
  wire       [7:0]    xil_SimpleDualBram_414_doutb;
  wire       [7:0]    xil_SimpleDualBram_415_doutb;
  wire       [7:0]    xil_SimpleDualBram_416_doutb;
  wire       [7:0]    xil_SimpleDualBram_417_doutb;
  wire       [7:0]    xil_SimpleDualBram_418_doutb;
  wire       [7:0]    xil_SimpleDualBram_419_doutb;
  wire       [7:0]    xil_SimpleDualBram_420_doutb;
  wire       [7:0]    xil_SimpleDualBram_421_doutb;
  wire       [7:0]    xil_SimpleDualBram_422_doutb;
  wire       [7:0]    xil_SimpleDualBram_423_doutb;
  wire       [7:0]    xil_SimpleDualBram_424_doutb;
  wire       [7:0]    xil_SimpleDualBram_425_doutb;
  wire       [7:0]    xil_SimpleDualBram_426_doutb;
  wire       [7:0]    xil_SimpleDualBram_427_doutb;
  wire       [7:0]    xil_SimpleDualBram_428_doutb;
  wire       [7:0]    xil_SimpleDualBram_429_doutb;
  wire       [7:0]    xil_SimpleDualBram_430_doutb;
  wire       [7:0]    xil_SimpleDualBram_431_doutb;
  wire       [7:0]    xil_SimpleDualBram_432_doutb;
  wire       [7:0]    xil_SimpleDualBram_433_doutb;
  wire       [7:0]    xil_SimpleDualBram_434_doutb;
  wire       [7:0]    xil_SimpleDualBram_435_doutb;
  wire       [7:0]    xil_SimpleDualBram_436_doutb;
  wire       [7:0]    xil_SimpleDualBram_437_doutb;
  wire       [7:0]    xil_SimpleDualBram_438_doutb;
  wire       [7:0]    xil_SimpleDualBram_439_doutb;
  wire       [7:0]    xil_SimpleDualBram_440_doutb;
  wire       [7:0]    xil_SimpleDualBram_441_doutb;
  wire       [7:0]    xil_SimpleDualBram_442_doutb;
  wire       [7:0]    xil_SimpleDualBram_443_doutb;
  wire       [7:0]    xil_SimpleDualBram_444_doutb;
  wire       [7:0]    xil_SimpleDualBram_445_doutb;
  wire       [7:0]    xil_SimpleDualBram_446_doutb;
  wire       [7:0]    xil_SimpleDualBram_447_doutb;
  wire       [7:0]    xil_SimpleDualBram_448_doutb;
  wire       [7:0]    xil_SimpleDualBram_449_doutb;
  wire       [7:0]    xil_SimpleDualBram_450_doutb;
  wire       [7:0]    xil_SimpleDualBram_451_doutb;
  wire       [7:0]    xil_SimpleDualBram_452_doutb;
  wire       [7:0]    xil_SimpleDualBram_453_doutb;
  wire       [7:0]    xil_SimpleDualBram_454_doutb;
  wire       [7:0]    xil_SimpleDualBram_455_doutb;
  wire       [7:0]    xil_SimpleDualBram_456_doutb;
  wire       [7:0]    xil_SimpleDualBram_457_doutb;
  wire       [7:0]    xil_SimpleDualBram_458_doutb;
  wire       [7:0]    xil_SimpleDualBram_459_doutb;
  wire       [7:0]    xil_SimpleDualBram_460_doutb;
  wire       [7:0]    xil_SimpleDualBram_461_doutb;
  wire       [7:0]    xil_SimpleDualBram_462_doutb;
  wire       [7:0]    xil_SimpleDualBram_463_doutb;
  wire       [7:0]    xil_SimpleDualBram_464_doutb;
  wire       [7:0]    xil_SimpleDualBram_465_doutb;
  wire       [7:0]    xil_SimpleDualBram_466_doutb;
  wire       [7:0]    xil_SimpleDualBram_467_doutb;
  wire       [7:0]    xil_SimpleDualBram_468_doutb;
  wire       [7:0]    xil_SimpleDualBram_469_doutb;
  wire       [7:0]    xil_SimpleDualBram_470_doutb;
  wire       [7:0]    xil_SimpleDualBram_471_doutb;
  wire       [7:0]    xil_SimpleDualBram_472_doutb;
  wire       [7:0]    xil_SimpleDualBram_473_doutb;
  wire       [7:0]    xil_SimpleDualBram_474_doutb;
  wire       [7:0]    xil_SimpleDualBram_475_doutb;
  wire       [7:0]    xil_SimpleDualBram_476_doutb;
  wire       [7:0]    xil_SimpleDualBram_477_doutb;
  wire       [7:0]    xil_SimpleDualBram_478_doutb;
  wire       [7:0]    xil_SimpleDualBram_479_doutb;
  wire       [7:0]    xil_SimpleDualBram_480_doutb;
  wire       [7:0]    xil_SimpleDualBram_481_doutb;
  wire       [7:0]    xil_SimpleDualBram_482_doutb;
  wire       [7:0]    xil_SimpleDualBram_483_doutb;
  wire       [7:0]    xil_SimpleDualBram_484_doutb;
  wire       [7:0]    xil_SimpleDualBram_485_doutb;
  wire       [7:0]    xil_SimpleDualBram_486_doutb;
  wire       [7:0]    xil_SimpleDualBram_487_doutb;
  wire       [7:0]    xil_SimpleDualBram_488_doutb;
  wire       [7:0]    xil_SimpleDualBram_489_doutb;
  wire       [7:0]    xil_SimpleDualBram_490_doutb;
  wire       [7:0]    xil_SimpleDualBram_491_doutb;
  wire       [7:0]    xil_SimpleDualBram_492_doutb;
  wire       [7:0]    xil_SimpleDualBram_493_doutb;
  wire       [7:0]    xil_SimpleDualBram_494_doutb;
  wire       [7:0]    xil_SimpleDualBram_495_doutb;
  wire       [7:0]    xil_SimpleDualBram_496_doutb;
  wire       [7:0]    xil_SimpleDualBram_497_doutb;
  wire       [7:0]    xil_SimpleDualBram_498_doutb;
  wire       [7:0]    xil_SimpleDualBram_499_doutb;
  wire       [7:0]    xil_SimpleDualBram_500_doutb;
  wire       [7:0]    xil_SimpleDualBram_501_doutb;
  wire       [7:0]    xil_SimpleDualBram_502_doutb;
  wire       [7:0]    xil_SimpleDualBram_503_doutb;
  wire       [7:0]    xil_SimpleDualBram_504_doutb;
  wire       [7:0]    xil_SimpleDualBram_505_doutb;
  wire       [7:0]    xil_SimpleDualBram_506_doutb;
  wire       [7:0]    xil_SimpleDualBram_507_doutb;
  wire       [7:0]    xil_SimpleDualBram_508_doutb;
  wire       [7:0]    xil_SimpleDualBram_509_doutb;
  wire       [7:0]    xil_SimpleDualBram_510_doutb;
  wire       [7:0]    xil_SimpleDualBram_511_doutb;
  wire       [15:0]   _zz_In_Row_Cnt_valid;
  wire       [12:0]   _zz_In_Row_Cnt_valid_1;
  wire       [15:0]   _zz_In_Col_Cnt_valid;
  wire       [15:0]   _zz_OutRow_Cnt_valid;
  wire       [15:0]   _zz_OutCol_Cnt_valid;
  wire       [15:0]   _zz_OutCol_Cnt_count_1;
  wire       [15:0]   _zz_Write_Row_Base_Addr;
  wire       [15:0]   _zz_addra;
  wire       [15:0]   _zz_addrb;
  wire       [0:0]    _zz_ena;
  wire       [15:0]   _zz_addra_1;
  wire       [15:0]   _zz_addrb_1;
  wire       [0:0]    _zz_ena_1;
  wire       [15:0]   _zz_addra_2;
  wire       [15:0]   _zz_addrb_2;
  wire       [0:0]    _zz_ena_2;
  wire       [15:0]   _zz_addra_3;
  wire       [15:0]   _zz_addrb_3;
  wire       [0:0]    _zz_ena_3;
  wire       [15:0]   _zz_addra_4;
  wire       [15:0]   _zz_addrb_4;
  wire       [0:0]    _zz_ena_4;
  wire       [15:0]   _zz_addra_5;
  wire       [15:0]   _zz_addrb_5;
  wire       [0:0]    _zz_ena_5;
  wire       [15:0]   _zz_addra_6;
  wire       [15:0]   _zz_addrb_6;
  wire       [0:0]    _zz_ena_6;
  wire       [15:0]   _zz_addra_7;
  wire       [15:0]   _zz_addrb_7;
  wire       [0:0]    _zz_ena_7;
  wire       [15:0]   _zz_addra_8;
  wire       [15:0]   _zz_addrb_8;
  wire       [0:0]    _zz_ena_8;
  wire       [15:0]   _zz_addra_9;
  wire       [15:0]   _zz_addrb_9;
  wire       [0:0]    _zz_ena_9;
  wire       [15:0]   _zz_addra_10;
  wire       [15:0]   _zz_addrb_10;
  wire       [0:0]    _zz_ena_10;
  wire       [15:0]   _zz_addra_11;
  wire       [15:0]   _zz_addrb_11;
  wire       [0:0]    _zz_ena_11;
  wire       [15:0]   _zz_addra_12;
  wire       [15:0]   _zz_addrb_12;
  wire       [0:0]    _zz_ena_12;
  wire       [15:0]   _zz_addra_13;
  wire       [15:0]   _zz_addrb_13;
  wire       [0:0]    _zz_ena_13;
  wire       [15:0]   _zz_addra_14;
  wire       [15:0]   _zz_addrb_14;
  wire       [0:0]    _zz_ena_14;
  wire       [15:0]   _zz_addra_15;
  wire       [15:0]   _zz_addrb_15;
  wire       [0:0]    _zz_ena_15;
  wire       [15:0]   _zz_addra_16;
  wire       [15:0]   _zz_addrb_16;
  wire       [0:0]    _zz_ena_16;
  wire       [15:0]   _zz_addra_17;
  wire       [15:0]   _zz_addrb_17;
  wire       [0:0]    _zz_ena_17;
  wire       [15:0]   _zz_addra_18;
  wire       [15:0]   _zz_addrb_18;
  wire       [0:0]    _zz_ena_18;
  wire       [15:0]   _zz_addra_19;
  wire       [15:0]   _zz_addrb_19;
  wire       [0:0]    _zz_ena_19;
  wire       [15:0]   _zz_addra_20;
  wire       [15:0]   _zz_addrb_20;
  wire       [0:0]    _zz_ena_20;
  wire       [15:0]   _zz_addra_21;
  wire       [15:0]   _zz_addrb_21;
  wire       [0:0]    _zz_ena_21;
  wire       [15:0]   _zz_addra_22;
  wire       [15:0]   _zz_addrb_22;
  wire       [0:0]    _zz_ena_22;
  wire       [15:0]   _zz_addra_23;
  wire       [15:0]   _zz_addrb_23;
  wire       [0:0]    _zz_ena_23;
  wire       [15:0]   _zz_addra_24;
  wire       [15:0]   _zz_addrb_24;
  wire       [0:0]    _zz_ena_24;
  wire       [15:0]   _zz_addra_25;
  wire       [15:0]   _zz_addrb_25;
  wire       [0:0]    _zz_ena_25;
  wire       [15:0]   _zz_addra_26;
  wire       [15:0]   _zz_addrb_26;
  wire       [0:0]    _zz_ena_26;
  wire       [15:0]   _zz_addra_27;
  wire       [15:0]   _zz_addrb_27;
  wire       [0:0]    _zz_ena_27;
  wire       [15:0]   _zz_addra_28;
  wire       [15:0]   _zz_addrb_28;
  wire       [0:0]    _zz_ena_28;
  wire       [15:0]   _zz_addra_29;
  wire       [15:0]   _zz_addrb_29;
  wire       [0:0]    _zz_ena_29;
  wire       [15:0]   _zz_addra_30;
  wire       [15:0]   _zz_addrb_30;
  wire       [0:0]    _zz_ena_30;
  wire       [15:0]   _zz_addra_31;
  wire       [15:0]   _zz_addrb_31;
  wire       [0:0]    _zz_ena_31;
  wire       [15:0]   _zz_addra_32;
  wire       [15:0]   _zz_addrb_32;
  wire       [0:0]    _zz_ena_32;
  wire       [15:0]   _zz_addra_33;
  wire       [15:0]   _zz_addrb_33;
  wire       [0:0]    _zz_ena_33;
  wire       [15:0]   _zz_addra_34;
  wire       [15:0]   _zz_addrb_34;
  wire       [0:0]    _zz_ena_34;
  wire       [15:0]   _zz_addra_35;
  wire       [15:0]   _zz_addrb_35;
  wire       [0:0]    _zz_ena_35;
  wire       [15:0]   _zz_addra_36;
  wire       [15:0]   _zz_addrb_36;
  wire       [0:0]    _zz_ena_36;
  wire       [15:0]   _zz_addra_37;
  wire       [15:0]   _zz_addrb_37;
  wire       [0:0]    _zz_ena_37;
  wire       [15:0]   _zz_addra_38;
  wire       [15:0]   _zz_addrb_38;
  wire       [0:0]    _zz_ena_38;
  wire       [15:0]   _zz_addra_39;
  wire       [15:0]   _zz_addrb_39;
  wire       [0:0]    _zz_ena_39;
  wire       [15:0]   _zz_addra_40;
  wire       [15:0]   _zz_addrb_40;
  wire       [0:0]    _zz_ena_40;
  wire       [15:0]   _zz_addra_41;
  wire       [15:0]   _zz_addrb_41;
  wire       [0:0]    _zz_ena_41;
  wire       [15:0]   _zz_addra_42;
  wire       [15:0]   _zz_addrb_42;
  wire       [0:0]    _zz_ena_42;
  wire       [15:0]   _zz_addra_43;
  wire       [15:0]   _zz_addrb_43;
  wire       [0:0]    _zz_ena_43;
  wire       [15:0]   _zz_addra_44;
  wire       [15:0]   _zz_addrb_44;
  wire       [0:0]    _zz_ena_44;
  wire       [15:0]   _zz_addra_45;
  wire       [15:0]   _zz_addrb_45;
  wire       [0:0]    _zz_ena_45;
  wire       [15:0]   _zz_addra_46;
  wire       [15:0]   _zz_addrb_46;
  wire       [0:0]    _zz_ena_46;
  wire       [15:0]   _zz_addra_47;
  wire       [15:0]   _zz_addrb_47;
  wire       [0:0]    _zz_ena_47;
  wire       [15:0]   _zz_addra_48;
  wire       [15:0]   _zz_addrb_48;
  wire       [0:0]    _zz_ena_48;
  wire       [15:0]   _zz_addra_49;
  wire       [15:0]   _zz_addrb_49;
  wire       [0:0]    _zz_ena_49;
  wire       [15:0]   _zz_addra_50;
  wire       [15:0]   _zz_addrb_50;
  wire       [0:0]    _zz_ena_50;
  wire       [15:0]   _zz_addra_51;
  wire       [15:0]   _zz_addrb_51;
  wire       [0:0]    _zz_ena_51;
  wire       [15:0]   _zz_addra_52;
  wire       [15:0]   _zz_addrb_52;
  wire       [0:0]    _zz_ena_52;
  wire       [15:0]   _zz_addra_53;
  wire       [15:0]   _zz_addrb_53;
  wire       [0:0]    _zz_ena_53;
  wire       [15:0]   _zz_addra_54;
  wire       [15:0]   _zz_addrb_54;
  wire       [0:0]    _zz_ena_54;
  wire       [15:0]   _zz_addra_55;
  wire       [15:0]   _zz_addrb_55;
  wire       [0:0]    _zz_ena_55;
  wire       [15:0]   _zz_addra_56;
  wire       [15:0]   _zz_addrb_56;
  wire       [0:0]    _zz_ena_56;
  wire       [15:0]   _zz_addra_57;
  wire       [15:0]   _zz_addrb_57;
  wire       [0:0]    _zz_ena_57;
  wire       [15:0]   _zz_addra_58;
  wire       [15:0]   _zz_addrb_58;
  wire       [0:0]    _zz_ena_58;
  wire       [15:0]   _zz_addra_59;
  wire       [15:0]   _zz_addrb_59;
  wire       [0:0]    _zz_ena_59;
  wire       [15:0]   _zz_addra_60;
  wire       [15:0]   _zz_addrb_60;
  wire       [0:0]    _zz_ena_60;
  wire       [15:0]   _zz_addra_61;
  wire       [15:0]   _zz_addrb_61;
  wire       [0:0]    _zz_ena_61;
  wire       [15:0]   _zz_addra_62;
  wire       [15:0]   _zz_addrb_62;
  wire       [0:0]    _zz_ena_62;
  wire       [15:0]   _zz_addra_63;
  wire       [15:0]   _zz_addrb_63;
  wire       [0:0]    _zz_ena_63;
  wire       [15:0]   _zz_addra_64;
  wire       [15:0]   _zz_addrb_64;
  wire       [0:0]    _zz_ena_64;
  wire       [15:0]   _zz_addra_65;
  wire       [15:0]   _zz_addrb_65;
  wire       [0:0]    _zz_ena_65;
  wire       [15:0]   _zz_addra_66;
  wire       [15:0]   _zz_addrb_66;
  wire       [0:0]    _zz_ena_66;
  wire       [15:0]   _zz_addra_67;
  wire       [15:0]   _zz_addrb_67;
  wire       [0:0]    _zz_ena_67;
  wire       [15:0]   _zz_addra_68;
  wire       [15:0]   _zz_addrb_68;
  wire       [0:0]    _zz_ena_68;
  wire       [15:0]   _zz_addra_69;
  wire       [15:0]   _zz_addrb_69;
  wire       [0:0]    _zz_ena_69;
  wire       [15:0]   _zz_addra_70;
  wire       [15:0]   _zz_addrb_70;
  wire       [0:0]    _zz_ena_70;
  wire       [15:0]   _zz_addra_71;
  wire       [15:0]   _zz_addrb_71;
  wire       [0:0]    _zz_ena_71;
  wire       [15:0]   _zz_addra_72;
  wire       [15:0]   _zz_addrb_72;
  wire       [0:0]    _zz_ena_72;
  wire       [15:0]   _zz_addra_73;
  wire       [15:0]   _zz_addrb_73;
  wire       [0:0]    _zz_ena_73;
  wire       [15:0]   _zz_addra_74;
  wire       [15:0]   _zz_addrb_74;
  wire       [0:0]    _zz_ena_74;
  wire       [15:0]   _zz_addra_75;
  wire       [15:0]   _zz_addrb_75;
  wire       [0:0]    _zz_ena_75;
  wire       [15:0]   _zz_addra_76;
  wire       [15:0]   _zz_addrb_76;
  wire       [0:0]    _zz_ena_76;
  wire       [15:0]   _zz_addra_77;
  wire       [15:0]   _zz_addrb_77;
  wire       [0:0]    _zz_ena_77;
  wire       [15:0]   _zz_addra_78;
  wire       [15:0]   _zz_addrb_78;
  wire       [0:0]    _zz_ena_78;
  wire       [15:0]   _zz_addra_79;
  wire       [15:0]   _zz_addrb_79;
  wire       [0:0]    _zz_ena_79;
  wire       [15:0]   _zz_addra_80;
  wire       [15:0]   _zz_addrb_80;
  wire       [0:0]    _zz_ena_80;
  wire       [15:0]   _zz_addra_81;
  wire       [15:0]   _zz_addrb_81;
  wire       [0:0]    _zz_ena_81;
  wire       [15:0]   _zz_addra_82;
  wire       [15:0]   _zz_addrb_82;
  wire       [0:0]    _zz_ena_82;
  wire       [15:0]   _zz_addra_83;
  wire       [15:0]   _zz_addrb_83;
  wire       [0:0]    _zz_ena_83;
  wire       [15:0]   _zz_addra_84;
  wire       [15:0]   _zz_addrb_84;
  wire       [0:0]    _zz_ena_84;
  wire       [15:0]   _zz_addra_85;
  wire       [15:0]   _zz_addrb_85;
  wire       [0:0]    _zz_ena_85;
  wire       [15:0]   _zz_addra_86;
  wire       [15:0]   _zz_addrb_86;
  wire       [0:0]    _zz_ena_86;
  wire       [15:0]   _zz_addra_87;
  wire       [15:0]   _zz_addrb_87;
  wire       [0:0]    _zz_ena_87;
  wire       [15:0]   _zz_addra_88;
  wire       [15:0]   _zz_addrb_88;
  wire       [0:0]    _zz_ena_88;
  wire       [15:0]   _zz_addra_89;
  wire       [15:0]   _zz_addrb_89;
  wire       [0:0]    _zz_ena_89;
  wire       [15:0]   _zz_addra_90;
  wire       [15:0]   _zz_addrb_90;
  wire       [0:0]    _zz_ena_90;
  wire       [15:0]   _zz_addra_91;
  wire       [15:0]   _zz_addrb_91;
  wire       [0:0]    _zz_ena_91;
  wire       [15:0]   _zz_addra_92;
  wire       [15:0]   _zz_addrb_92;
  wire       [0:0]    _zz_ena_92;
  wire       [15:0]   _zz_addra_93;
  wire       [15:0]   _zz_addrb_93;
  wire       [0:0]    _zz_ena_93;
  wire       [15:0]   _zz_addra_94;
  wire       [15:0]   _zz_addrb_94;
  wire       [0:0]    _zz_ena_94;
  wire       [15:0]   _zz_addra_95;
  wire       [15:0]   _zz_addrb_95;
  wire       [0:0]    _zz_ena_95;
  wire       [15:0]   _zz_addra_96;
  wire       [15:0]   _zz_addrb_96;
  wire       [0:0]    _zz_ena_96;
  wire       [15:0]   _zz_addra_97;
  wire       [15:0]   _zz_addrb_97;
  wire       [0:0]    _zz_ena_97;
  wire       [15:0]   _zz_addra_98;
  wire       [15:0]   _zz_addrb_98;
  wire       [0:0]    _zz_ena_98;
  wire       [15:0]   _zz_addra_99;
  wire       [15:0]   _zz_addrb_99;
  wire       [0:0]    _zz_ena_99;
  wire       [15:0]   _zz_addra_100;
  wire       [15:0]   _zz_addrb_100;
  wire       [0:0]    _zz_ena_100;
  wire       [15:0]   _zz_addra_101;
  wire       [15:0]   _zz_addrb_101;
  wire       [0:0]    _zz_ena_101;
  wire       [15:0]   _zz_addra_102;
  wire       [15:0]   _zz_addrb_102;
  wire       [0:0]    _zz_ena_102;
  wire       [15:0]   _zz_addra_103;
  wire       [15:0]   _zz_addrb_103;
  wire       [0:0]    _zz_ena_103;
  wire       [15:0]   _zz_addra_104;
  wire       [15:0]   _zz_addrb_104;
  wire       [0:0]    _zz_ena_104;
  wire       [15:0]   _zz_addra_105;
  wire       [15:0]   _zz_addrb_105;
  wire       [0:0]    _zz_ena_105;
  wire       [15:0]   _zz_addra_106;
  wire       [15:0]   _zz_addrb_106;
  wire       [0:0]    _zz_ena_106;
  wire       [15:0]   _zz_addra_107;
  wire       [15:0]   _zz_addrb_107;
  wire       [0:0]    _zz_ena_107;
  wire       [15:0]   _zz_addra_108;
  wire       [15:0]   _zz_addrb_108;
  wire       [0:0]    _zz_ena_108;
  wire       [15:0]   _zz_addra_109;
  wire       [15:0]   _zz_addrb_109;
  wire       [0:0]    _zz_ena_109;
  wire       [15:0]   _zz_addra_110;
  wire       [15:0]   _zz_addrb_110;
  wire       [0:0]    _zz_ena_110;
  wire       [15:0]   _zz_addra_111;
  wire       [15:0]   _zz_addrb_111;
  wire       [0:0]    _zz_ena_111;
  wire       [15:0]   _zz_addra_112;
  wire       [15:0]   _zz_addrb_112;
  wire       [0:0]    _zz_ena_112;
  wire       [15:0]   _zz_addra_113;
  wire       [15:0]   _zz_addrb_113;
  wire       [0:0]    _zz_ena_113;
  wire       [15:0]   _zz_addra_114;
  wire       [15:0]   _zz_addrb_114;
  wire       [0:0]    _zz_ena_114;
  wire       [15:0]   _zz_addra_115;
  wire       [15:0]   _zz_addrb_115;
  wire       [0:0]    _zz_ena_115;
  wire       [15:0]   _zz_addra_116;
  wire       [15:0]   _zz_addrb_116;
  wire       [0:0]    _zz_ena_116;
  wire       [15:0]   _zz_addra_117;
  wire       [15:0]   _zz_addrb_117;
  wire       [0:0]    _zz_ena_117;
  wire       [15:0]   _zz_addra_118;
  wire       [15:0]   _zz_addrb_118;
  wire       [0:0]    _zz_ena_118;
  wire       [15:0]   _zz_addra_119;
  wire       [15:0]   _zz_addrb_119;
  wire       [0:0]    _zz_ena_119;
  wire       [15:0]   _zz_addra_120;
  wire       [15:0]   _zz_addrb_120;
  wire       [0:0]    _zz_ena_120;
  wire       [15:0]   _zz_addra_121;
  wire       [15:0]   _zz_addrb_121;
  wire       [0:0]    _zz_ena_121;
  wire       [15:0]   _zz_addra_122;
  wire       [15:0]   _zz_addrb_122;
  wire       [0:0]    _zz_ena_122;
  wire       [15:0]   _zz_addra_123;
  wire       [15:0]   _zz_addrb_123;
  wire       [0:0]    _zz_ena_123;
  wire       [15:0]   _zz_addra_124;
  wire       [15:0]   _zz_addrb_124;
  wire       [0:0]    _zz_ena_124;
  wire       [15:0]   _zz_addra_125;
  wire       [15:0]   _zz_addrb_125;
  wire       [0:0]    _zz_ena_125;
  wire       [15:0]   _zz_addra_126;
  wire       [15:0]   _zz_addrb_126;
  wire       [0:0]    _zz_ena_126;
  wire       [15:0]   _zz_addra_127;
  wire       [15:0]   _zz_addrb_127;
  wire       [0:0]    _zz_ena_127;
  wire       [15:0]   _zz_addra_128;
  wire       [15:0]   _zz_addrb_128;
  wire       [0:0]    _zz_ena_128;
  wire       [15:0]   _zz_addra_129;
  wire       [15:0]   _zz_addrb_129;
  wire       [0:0]    _zz_ena_129;
  wire       [15:0]   _zz_addra_130;
  wire       [15:0]   _zz_addrb_130;
  wire       [0:0]    _zz_ena_130;
  wire       [15:0]   _zz_addra_131;
  wire       [15:0]   _zz_addrb_131;
  wire       [0:0]    _zz_ena_131;
  wire       [15:0]   _zz_addra_132;
  wire       [15:0]   _zz_addrb_132;
  wire       [0:0]    _zz_ena_132;
  wire       [15:0]   _zz_addra_133;
  wire       [15:0]   _zz_addrb_133;
  wire       [0:0]    _zz_ena_133;
  wire       [15:0]   _zz_addra_134;
  wire       [15:0]   _zz_addrb_134;
  wire       [0:0]    _zz_ena_134;
  wire       [15:0]   _zz_addra_135;
  wire       [15:0]   _zz_addrb_135;
  wire       [0:0]    _zz_ena_135;
  wire       [15:0]   _zz_addra_136;
  wire       [15:0]   _zz_addrb_136;
  wire       [0:0]    _zz_ena_136;
  wire       [15:0]   _zz_addra_137;
  wire       [15:0]   _zz_addrb_137;
  wire       [0:0]    _zz_ena_137;
  wire       [15:0]   _zz_addra_138;
  wire       [15:0]   _zz_addrb_138;
  wire       [0:0]    _zz_ena_138;
  wire       [15:0]   _zz_addra_139;
  wire       [15:0]   _zz_addrb_139;
  wire       [0:0]    _zz_ena_139;
  wire       [15:0]   _zz_addra_140;
  wire       [15:0]   _zz_addrb_140;
  wire       [0:0]    _zz_ena_140;
  wire       [15:0]   _zz_addra_141;
  wire       [15:0]   _zz_addrb_141;
  wire       [0:0]    _zz_ena_141;
  wire       [15:0]   _zz_addra_142;
  wire       [15:0]   _zz_addrb_142;
  wire       [0:0]    _zz_ena_142;
  wire       [15:0]   _zz_addra_143;
  wire       [15:0]   _zz_addrb_143;
  wire       [0:0]    _zz_ena_143;
  wire       [15:0]   _zz_addra_144;
  wire       [15:0]   _zz_addrb_144;
  wire       [0:0]    _zz_ena_144;
  wire       [15:0]   _zz_addra_145;
  wire       [15:0]   _zz_addrb_145;
  wire       [0:0]    _zz_ena_145;
  wire       [15:0]   _zz_addra_146;
  wire       [15:0]   _zz_addrb_146;
  wire       [0:0]    _zz_ena_146;
  wire       [15:0]   _zz_addra_147;
  wire       [15:0]   _zz_addrb_147;
  wire       [0:0]    _zz_ena_147;
  wire       [15:0]   _zz_addra_148;
  wire       [15:0]   _zz_addrb_148;
  wire       [0:0]    _zz_ena_148;
  wire       [15:0]   _zz_addra_149;
  wire       [15:0]   _zz_addrb_149;
  wire       [0:0]    _zz_ena_149;
  wire       [15:0]   _zz_addra_150;
  wire       [15:0]   _zz_addrb_150;
  wire       [0:0]    _zz_ena_150;
  wire       [15:0]   _zz_addra_151;
  wire       [15:0]   _zz_addrb_151;
  wire       [0:0]    _zz_ena_151;
  wire       [15:0]   _zz_addra_152;
  wire       [15:0]   _zz_addrb_152;
  wire       [0:0]    _zz_ena_152;
  wire       [15:0]   _zz_addra_153;
  wire       [15:0]   _zz_addrb_153;
  wire       [0:0]    _zz_ena_153;
  wire       [15:0]   _zz_addra_154;
  wire       [15:0]   _zz_addrb_154;
  wire       [0:0]    _zz_ena_154;
  wire       [15:0]   _zz_addra_155;
  wire       [15:0]   _zz_addrb_155;
  wire       [0:0]    _zz_ena_155;
  wire       [15:0]   _zz_addra_156;
  wire       [15:0]   _zz_addrb_156;
  wire       [0:0]    _zz_ena_156;
  wire       [15:0]   _zz_addra_157;
  wire       [15:0]   _zz_addrb_157;
  wire       [0:0]    _zz_ena_157;
  wire       [15:0]   _zz_addra_158;
  wire       [15:0]   _zz_addrb_158;
  wire       [0:0]    _zz_ena_158;
  wire       [15:0]   _zz_addra_159;
  wire       [15:0]   _zz_addrb_159;
  wire       [0:0]    _zz_ena_159;
  wire       [15:0]   _zz_addra_160;
  wire       [15:0]   _zz_addrb_160;
  wire       [0:0]    _zz_ena_160;
  wire       [15:0]   _zz_addra_161;
  wire       [15:0]   _zz_addrb_161;
  wire       [0:0]    _zz_ena_161;
  wire       [15:0]   _zz_addra_162;
  wire       [15:0]   _zz_addrb_162;
  wire       [0:0]    _zz_ena_162;
  wire       [15:0]   _zz_addra_163;
  wire       [15:0]   _zz_addrb_163;
  wire       [0:0]    _zz_ena_163;
  wire       [15:0]   _zz_addra_164;
  wire       [15:0]   _zz_addrb_164;
  wire       [0:0]    _zz_ena_164;
  wire       [15:0]   _zz_addra_165;
  wire       [15:0]   _zz_addrb_165;
  wire       [0:0]    _zz_ena_165;
  wire       [15:0]   _zz_addra_166;
  wire       [15:0]   _zz_addrb_166;
  wire       [0:0]    _zz_ena_166;
  wire       [15:0]   _zz_addra_167;
  wire       [15:0]   _zz_addrb_167;
  wire       [0:0]    _zz_ena_167;
  wire       [15:0]   _zz_addra_168;
  wire       [15:0]   _zz_addrb_168;
  wire       [0:0]    _zz_ena_168;
  wire       [15:0]   _zz_addra_169;
  wire       [15:0]   _zz_addrb_169;
  wire       [0:0]    _zz_ena_169;
  wire       [15:0]   _zz_addra_170;
  wire       [15:0]   _zz_addrb_170;
  wire       [0:0]    _zz_ena_170;
  wire       [15:0]   _zz_addra_171;
  wire       [15:0]   _zz_addrb_171;
  wire       [0:0]    _zz_ena_171;
  wire       [15:0]   _zz_addra_172;
  wire       [15:0]   _zz_addrb_172;
  wire       [0:0]    _zz_ena_172;
  wire       [15:0]   _zz_addra_173;
  wire       [15:0]   _zz_addrb_173;
  wire       [0:0]    _zz_ena_173;
  wire       [15:0]   _zz_addra_174;
  wire       [15:0]   _zz_addrb_174;
  wire       [0:0]    _zz_ena_174;
  wire       [15:0]   _zz_addra_175;
  wire       [15:0]   _zz_addrb_175;
  wire       [0:0]    _zz_ena_175;
  wire       [15:0]   _zz_addra_176;
  wire       [15:0]   _zz_addrb_176;
  wire       [0:0]    _zz_ena_176;
  wire       [15:0]   _zz_addra_177;
  wire       [15:0]   _zz_addrb_177;
  wire       [0:0]    _zz_ena_177;
  wire       [15:0]   _zz_addra_178;
  wire       [15:0]   _zz_addrb_178;
  wire       [0:0]    _zz_ena_178;
  wire       [15:0]   _zz_addra_179;
  wire       [15:0]   _zz_addrb_179;
  wire       [0:0]    _zz_ena_179;
  wire       [15:0]   _zz_addra_180;
  wire       [15:0]   _zz_addrb_180;
  wire       [0:0]    _zz_ena_180;
  wire       [15:0]   _zz_addra_181;
  wire       [15:0]   _zz_addrb_181;
  wire       [0:0]    _zz_ena_181;
  wire       [15:0]   _zz_addra_182;
  wire       [15:0]   _zz_addrb_182;
  wire       [0:0]    _zz_ena_182;
  wire       [15:0]   _zz_addra_183;
  wire       [15:0]   _zz_addrb_183;
  wire       [0:0]    _zz_ena_183;
  wire       [15:0]   _zz_addra_184;
  wire       [15:0]   _zz_addrb_184;
  wire       [0:0]    _zz_ena_184;
  wire       [15:0]   _zz_addra_185;
  wire       [15:0]   _zz_addrb_185;
  wire       [0:0]    _zz_ena_185;
  wire       [15:0]   _zz_addra_186;
  wire       [15:0]   _zz_addrb_186;
  wire       [0:0]    _zz_ena_186;
  wire       [15:0]   _zz_addra_187;
  wire       [15:0]   _zz_addrb_187;
  wire       [0:0]    _zz_ena_187;
  wire       [15:0]   _zz_addra_188;
  wire       [15:0]   _zz_addrb_188;
  wire       [0:0]    _zz_ena_188;
  wire       [15:0]   _zz_addra_189;
  wire       [15:0]   _zz_addrb_189;
  wire       [0:0]    _zz_ena_189;
  wire       [15:0]   _zz_addra_190;
  wire       [15:0]   _zz_addrb_190;
  wire       [0:0]    _zz_ena_190;
  wire       [15:0]   _zz_addra_191;
  wire       [15:0]   _zz_addrb_191;
  wire       [0:0]    _zz_ena_191;
  wire       [15:0]   _zz_addra_192;
  wire       [15:0]   _zz_addrb_192;
  wire       [0:0]    _zz_ena_192;
  wire       [15:0]   _zz_addra_193;
  wire       [15:0]   _zz_addrb_193;
  wire       [0:0]    _zz_ena_193;
  wire       [15:0]   _zz_addra_194;
  wire       [15:0]   _zz_addrb_194;
  wire       [0:0]    _zz_ena_194;
  wire       [15:0]   _zz_addra_195;
  wire       [15:0]   _zz_addrb_195;
  wire       [0:0]    _zz_ena_195;
  wire       [15:0]   _zz_addra_196;
  wire       [15:0]   _zz_addrb_196;
  wire       [0:0]    _zz_ena_196;
  wire       [15:0]   _zz_addra_197;
  wire       [15:0]   _zz_addrb_197;
  wire       [0:0]    _zz_ena_197;
  wire       [15:0]   _zz_addra_198;
  wire       [15:0]   _zz_addrb_198;
  wire       [0:0]    _zz_ena_198;
  wire       [15:0]   _zz_addra_199;
  wire       [15:0]   _zz_addrb_199;
  wire       [0:0]    _zz_ena_199;
  wire       [15:0]   _zz_addra_200;
  wire       [15:0]   _zz_addrb_200;
  wire       [0:0]    _zz_ena_200;
  wire       [15:0]   _zz_addra_201;
  wire       [15:0]   _zz_addrb_201;
  wire       [0:0]    _zz_ena_201;
  wire       [15:0]   _zz_addra_202;
  wire       [15:0]   _zz_addrb_202;
  wire       [0:0]    _zz_ena_202;
  wire       [15:0]   _zz_addra_203;
  wire       [15:0]   _zz_addrb_203;
  wire       [0:0]    _zz_ena_203;
  wire       [15:0]   _zz_addra_204;
  wire       [15:0]   _zz_addrb_204;
  wire       [0:0]    _zz_ena_204;
  wire       [15:0]   _zz_addra_205;
  wire       [15:0]   _zz_addrb_205;
  wire       [0:0]    _zz_ena_205;
  wire       [15:0]   _zz_addra_206;
  wire       [15:0]   _zz_addrb_206;
  wire       [0:0]    _zz_ena_206;
  wire       [15:0]   _zz_addra_207;
  wire       [15:0]   _zz_addrb_207;
  wire       [0:0]    _zz_ena_207;
  wire       [15:0]   _zz_addra_208;
  wire       [15:0]   _zz_addrb_208;
  wire       [0:0]    _zz_ena_208;
  wire       [15:0]   _zz_addra_209;
  wire       [15:0]   _zz_addrb_209;
  wire       [0:0]    _zz_ena_209;
  wire       [15:0]   _zz_addra_210;
  wire       [15:0]   _zz_addrb_210;
  wire       [0:0]    _zz_ena_210;
  wire       [15:0]   _zz_addra_211;
  wire       [15:0]   _zz_addrb_211;
  wire       [0:0]    _zz_ena_211;
  wire       [15:0]   _zz_addra_212;
  wire       [15:0]   _zz_addrb_212;
  wire       [0:0]    _zz_ena_212;
  wire       [15:0]   _zz_addra_213;
  wire       [15:0]   _zz_addrb_213;
  wire       [0:0]    _zz_ena_213;
  wire       [15:0]   _zz_addra_214;
  wire       [15:0]   _zz_addrb_214;
  wire       [0:0]    _zz_ena_214;
  wire       [15:0]   _zz_addra_215;
  wire       [15:0]   _zz_addrb_215;
  wire       [0:0]    _zz_ena_215;
  wire       [15:0]   _zz_addra_216;
  wire       [15:0]   _zz_addrb_216;
  wire       [0:0]    _zz_ena_216;
  wire       [15:0]   _zz_addra_217;
  wire       [15:0]   _zz_addrb_217;
  wire       [0:0]    _zz_ena_217;
  wire       [15:0]   _zz_addra_218;
  wire       [15:0]   _zz_addrb_218;
  wire       [0:0]    _zz_ena_218;
  wire       [15:0]   _zz_addra_219;
  wire       [15:0]   _zz_addrb_219;
  wire       [0:0]    _zz_ena_219;
  wire       [15:0]   _zz_addra_220;
  wire       [15:0]   _zz_addrb_220;
  wire       [0:0]    _zz_ena_220;
  wire       [15:0]   _zz_addra_221;
  wire       [15:0]   _zz_addrb_221;
  wire       [0:0]    _zz_ena_221;
  wire       [15:0]   _zz_addra_222;
  wire       [15:0]   _zz_addrb_222;
  wire       [0:0]    _zz_ena_222;
  wire       [15:0]   _zz_addra_223;
  wire       [15:0]   _zz_addrb_223;
  wire       [0:0]    _zz_ena_223;
  wire       [15:0]   _zz_addra_224;
  wire       [15:0]   _zz_addrb_224;
  wire       [0:0]    _zz_ena_224;
  wire       [15:0]   _zz_addra_225;
  wire       [15:0]   _zz_addrb_225;
  wire       [0:0]    _zz_ena_225;
  wire       [15:0]   _zz_addra_226;
  wire       [15:0]   _zz_addrb_226;
  wire       [0:0]    _zz_ena_226;
  wire       [15:0]   _zz_addra_227;
  wire       [15:0]   _zz_addrb_227;
  wire       [0:0]    _zz_ena_227;
  wire       [15:0]   _zz_addra_228;
  wire       [15:0]   _zz_addrb_228;
  wire       [0:0]    _zz_ena_228;
  wire       [15:0]   _zz_addra_229;
  wire       [15:0]   _zz_addrb_229;
  wire       [0:0]    _zz_ena_229;
  wire       [15:0]   _zz_addra_230;
  wire       [15:0]   _zz_addrb_230;
  wire       [0:0]    _zz_ena_230;
  wire       [15:0]   _zz_addra_231;
  wire       [15:0]   _zz_addrb_231;
  wire       [0:0]    _zz_ena_231;
  wire       [15:0]   _zz_addra_232;
  wire       [15:0]   _zz_addrb_232;
  wire       [0:0]    _zz_ena_232;
  wire       [15:0]   _zz_addra_233;
  wire       [15:0]   _zz_addrb_233;
  wire       [0:0]    _zz_ena_233;
  wire       [15:0]   _zz_addra_234;
  wire       [15:0]   _zz_addrb_234;
  wire       [0:0]    _zz_ena_234;
  wire       [15:0]   _zz_addra_235;
  wire       [15:0]   _zz_addrb_235;
  wire       [0:0]    _zz_ena_235;
  wire       [15:0]   _zz_addra_236;
  wire       [15:0]   _zz_addrb_236;
  wire       [0:0]    _zz_ena_236;
  wire       [15:0]   _zz_addra_237;
  wire       [15:0]   _zz_addrb_237;
  wire       [0:0]    _zz_ena_237;
  wire       [15:0]   _zz_addra_238;
  wire       [15:0]   _zz_addrb_238;
  wire       [0:0]    _zz_ena_238;
  wire       [15:0]   _zz_addra_239;
  wire       [15:0]   _zz_addrb_239;
  wire       [0:0]    _zz_ena_239;
  wire       [15:0]   _zz_addra_240;
  wire       [15:0]   _zz_addrb_240;
  wire       [0:0]    _zz_ena_240;
  wire       [15:0]   _zz_addra_241;
  wire       [15:0]   _zz_addrb_241;
  wire       [0:0]    _zz_ena_241;
  wire       [15:0]   _zz_addra_242;
  wire       [15:0]   _zz_addrb_242;
  wire       [0:0]    _zz_ena_242;
  wire       [15:0]   _zz_addra_243;
  wire       [15:0]   _zz_addrb_243;
  wire       [0:0]    _zz_ena_243;
  wire       [15:0]   _zz_addra_244;
  wire       [15:0]   _zz_addrb_244;
  wire       [0:0]    _zz_ena_244;
  wire       [15:0]   _zz_addra_245;
  wire       [15:0]   _zz_addrb_245;
  wire       [0:0]    _zz_ena_245;
  wire       [15:0]   _zz_addra_246;
  wire       [15:0]   _zz_addrb_246;
  wire       [0:0]    _zz_ena_246;
  wire       [15:0]   _zz_addra_247;
  wire       [15:0]   _zz_addrb_247;
  wire       [0:0]    _zz_ena_247;
  wire       [15:0]   _zz_addra_248;
  wire       [15:0]   _zz_addrb_248;
  wire       [0:0]    _zz_ena_248;
  wire       [15:0]   _zz_addra_249;
  wire       [15:0]   _zz_addrb_249;
  wire       [0:0]    _zz_ena_249;
  wire       [15:0]   _zz_addra_250;
  wire       [15:0]   _zz_addrb_250;
  wire       [0:0]    _zz_ena_250;
  wire       [15:0]   _zz_addra_251;
  wire       [15:0]   _zz_addrb_251;
  wire       [0:0]    _zz_ena_251;
  wire       [15:0]   _zz_addra_252;
  wire       [15:0]   _zz_addrb_252;
  wire       [0:0]    _zz_ena_252;
  wire       [15:0]   _zz_addra_253;
  wire       [15:0]   _zz_addrb_253;
  wire       [0:0]    _zz_ena_253;
  wire       [15:0]   _zz_addra_254;
  wire       [15:0]   _zz_addrb_254;
  wire       [0:0]    _zz_ena_254;
  wire       [15:0]   _zz_addra_255;
  wire       [15:0]   _zz_addrb_255;
  wire       [0:0]    _zz_ena_255;
  wire       [15:0]   _zz_addra_256;
  wire       [15:0]   _zz_addrb_256;
  wire       [0:0]    _zz_ena_256;
  wire       [15:0]   _zz_addra_257;
  wire       [15:0]   _zz_addrb_257;
  wire       [0:0]    _zz_ena_257;
  wire       [15:0]   _zz_addra_258;
  wire       [15:0]   _zz_addrb_258;
  wire       [0:0]    _zz_ena_258;
  wire       [15:0]   _zz_addra_259;
  wire       [15:0]   _zz_addrb_259;
  wire       [0:0]    _zz_ena_259;
  wire       [15:0]   _zz_addra_260;
  wire       [15:0]   _zz_addrb_260;
  wire       [0:0]    _zz_ena_260;
  wire       [15:0]   _zz_addra_261;
  wire       [15:0]   _zz_addrb_261;
  wire       [0:0]    _zz_ena_261;
  wire       [15:0]   _zz_addra_262;
  wire       [15:0]   _zz_addrb_262;
  wire       [0:0]    _zz_ena_262;
  wire       [15:0]   _zz_addra_263;
  wire       [15:0]   _zz_addrb_263;
  wire       [0:0]    _zz_ena_263;
  wire       [15:0]   _zz_addra_264;
  wire       [15:0]   _zz_addrb_264;
  wire       [0:0]    _zz_ena_264;
  wire       [15:0]   _zz_addra_265;
  wire       [15:0]   _zz_addrb_265;
  wire       [0:0]    _zz_ena_265;
  wire       [15:0]   _zz_addra_266;
  wire       [15:0]   _zz_addrb_266;
  wire       [0:0]    _zz_ena_266;
  wire       [15:0]   _zz_addra_267;
  wire       [15:0]   _zz_addrb_267;
  wire       [0:0]    _zz_ena_267;
  wire       [15:0]   _zz_addra_268;
  wire       [15:0]   _zz_addrb_268;
  wire       [0:0]    _zz_ena_268;
  wire       [15:0]   _zz_addra_269;
  wire       [15:0]   _zz_addrb_269;
  wire       [0:0]    _zz_ena_269;
  wire       [15:0]   _zz_addra_270;
  wire       [15:0]   _zz_addrb_270;
  wire       [0:0]    _zz_ena_270;
  wire       [15:0]   _zz_addra_271;
  wire       [15:0]   _zz_addrb_271;
  wire       [0:0]    _zz_ena_271;
  wire       [15:0]   _zz_addra_272;
  wire       [15:0]   _zz_addrb_272;
  wire       [0:0]    _zz_ena_272;
  wire       [15:0]   _zz_addra_273;
  wire       [15:0]   _zz_addrb_273;
  wire       [0:0]    _zz_ena_273;
  wire       [15:0]   _zz_addra_274;
  wire       [15:0]   _zz_addrb_274;
  wire       [0:0]    _zz_ena_274;
  wire       [15:0]   _zz_addra_275;
  wire       [15:0]   _zz_addrb_275;
  wire       [0:0]    _zz_ena_275;
  wire       [15:0]   _zz_addra_276;
  wire       [15:0]   _zz_addrb_276;
  wire       [0:0]    _zz_ena_276;
  wire       [15:0]   _zz_addra_277;
  wire       [15:0]   _zz_addrb_277;
  wire       [0:0]    _zz_ena_277;
  wire       [15:0]   _zz_addra_278;
  wire       [15:0]   _zz_addrb_278;
  wire       [0:0]    _zz_ena_278;
  wire       [15:0]   _zz_addra_279;
  wire       [15:0]   _zz_addrb_279;
  wire       [0:0]    _zz_ena_279;
  wire       [15:0]   _zz_addra_280;
  wire       [15:0]   _zz_addrb_280;
  wire       [0:0]    _zz_ena_280;
  wire       [15:0]   _zz_addra_281;
  wire       [15:0]   _zz_addrb_281;
  wire       [0:0]    _zz_ena_281;
  wire       [15:0]   _zz_addra_282;
  wire       [15:0]   _zz_addrb_282;
  wire       [0:0]    _zz_ena_282;
  wire       [15:0]   _zz_addra_283;
  wire       [15:0]   _zz_addrb_283;
  wire       [0:0]    _zz_ena_283;
  wire       [15:0]   _zz_addra_284;
  wire       [15:0]   _zz_addrb_284;
  wire       [0:0]    _zz_ena_284;
  wire       [15:0]   _zz_addra_285;
  wire       [15:0]   _zz_addrb_285;
  wire       [0:0]    _zz_ena_285;
  wire       [15:0]   _zz_addra_286;
  wire       [15:0]   _zz_addrb_286;
  wire       [0:0]    _zz_ena_286;
  wire       [15:0]   _zz_addra_287;
  wire       [15:0]   _zz_addrb_287;
  wire       [0:0]    _zz_ena_287;
  wire       [15:0]   _zz_addra_288;
  wire       [15:0]   _zz_addrb_288;
  wire       [0:0]    _zz_ena_288;
  wire       [15:0]   _zz_addra_289;
  wire       [15:0]   _zz_addrb_289;
  wire       [0:0]    _zz_ena_289;
  wire       [15:0]   _zz_addra_290;
  wire       [15:0]   _zz_addrb_290;
  wire       [0:0]    _zz_ena_290;
  wire       [15:0]   _zz_addra_291;
  wire       [15:0]   _zz_addrb_291;
  wire       [0:0]    _zz_ena_291;
  wire       [15:0]   _zz_addra_292;
  wire       [15:0]   _zz_addrb_292;
  wire       [0:0]    _zz_ena_292;
  wire       [15:0]   _zz_addra_293;
  wire       [15:0]   _zz_addrb_293;
  wire       [0:0]    _zz_ena_293;
  wire       [15:0]   _zz_addra_294;
  wire       [15:0]   _zz_addrb_294;
  wire       [0:0]    _zz_ena_294;
  wire       [15:0]   _zz_addra_295;
  wire       [15:0]   _zz_addrb_295;
  wire       [0:0]    _zz_ena_295;
  wire       [15:0]   _zz_addra_296;
  wire       [15:0]   _zz_addrb_296;
  wire       [0:0]    _zz_ena_296;
  wire       [15:0]   _zz_addra_297;
  wire       [15:0]   _zz_addrb_297;
  wire       [0:0]    _zz_ena_297;
  wire       [15:0]   _zz_addra_298;
  wire       [15:0]   _zz_addrb_298;
  wire       [0:0]    _zz_ena_298;
  wire       [15:0]   _zz_addra_299;
  wire       [15:0]   _zz_addrb_299;
  wire       [0:0]    _zz_ena_299;
  wire       [15:0]   _zz_addra_300;
  wire       [15:0]   _zz_addrb_300;
  wire       [0:0]    _zz_ena_300;
  wire       [15:0]   _zz_addra_301;
  wire       [15:0]   _zz_addrb_301;
  wire       [0:0]    _zz_ena_301;
  wire       [15:0]   _zz_addra_302;
  wire       [15:0]   _zz_addrb_302;
  wire       [0:0]    _zz_ena_302;
  wire       [15:0]   _zz_addra_303;
  wire       [15:0]   _zz_addrb_303;
  wire       [0:0]    _zz_ena_303;
  wire       [15:0]   _zz_addra_304;
  wire       [15:0]   _zz_addrb_304;
  wire       [0:0]    _zz_ena_304;
  wire       [15:0]   _zz_addra_305;
  wire       [15:0]   _zz_addrb_305;
  wire       [0:0]    _zz_ena_305;
  wire       [15:0]   _zz_addra_306;
  wire       [15:0]   _zz_addrb_306;
  wire       [0:0]    _zz_ena_306;
  wire       [15:0]   _zz_addra_307;
  wire       [15:0]   _zz_addrb_307;
  wire       [0:0]    _zz_ena_307;
  wire       [15:0]   _zz_addra_308;
  wire       [15:0]   _zz_addrb_308;
  wire       [0:0]    _zz_ena_308;
  wire       [15:0]   _zz_addra_309;
  wire       [15:0]   _zz_addrb_309;
  wire       [0:0]    _zz_ena_309;
  wire       [15:0]   _zz_addra_310;
  wire       [15:0]   _zz_addrb_310;
  wire       [0:0]    _zz_ena_310;
  wire       [15:0]   _zz_addra_311;
  wire       [15:0]   _zz_addrb_311;
  wire       [0:0]    _zz_ena_311;
  wire       [15:0]   _zz_addra_312;
  wire       [15:0]   _zz_addrb_312;
  wire       [0:0]    _zz_ena_312;
  wire       [15:0]   _zz_addra_313;
  wire       [15:0]   _zz_addrb_313;
  wire       [0:0]    _zz_ena_313;
  wire       [15:0]   _zz_addra_314;
  wire       [15:0]   _zz_addrb_314;
  wire       [0:0]    _zz_ena_314;
  wire       [15:0]   _zz_addra_315;
  wire       [15:0]   _zz_addrb_315;
  wire       [0:0]    _zz_ena_315;
  wire       [15:0]   _zz_addra_316;
  wire       [15:0]   _zz_addrb_316;
  wire       [0:0]    _zz_ena_316;
  wire       [15:0]   _zz_addra_317;
  wire       [15:0]   _zz_addrb_317;
  wire       [0:0]    _zz_ena_317;
  wire       [15:0]   _zz_addra_318;
  wire       [15:0]   _zz_addrb_318;
  wire       [0:0]    _zz_ena_318;
  wire       [15:0]   _zz_addra_319;
  wire       [15:0]   _zz_addrb_319;
  wire       [0:0]    _zz_ena_319;
  wire       [15:0]   _zz_addra_320;
  wire       [15:0]   _zz_addrb_320;
  wire       [0:0]    _zz_ena_320;
  wire       [15:0]   _zz_addra_321;
  wire       [15:0]   _zz_addrb_321;
  wire       [0:0]    _zz_ena_321;
  wire       [15:0]   _zz_addra_322;
  wire       [15:0]   _zz_addrb_322;
  wire       [0:0]    _zz_ena_322;
  wire       [15:0]   _zz_addra_323;
  wire       [15:0]   _zz_addrb_323;
  wire       [0:0]    _zz_ena_323;
  wire       [15:0]   _zz_addra_324;
  wire       [15:0]   _zz_addrb_324;
  wire       [0:0]    _zz_ena_324;
  wire       [15:0]   _zz_addra_325;
  wire       [15:0]   _zz_addrb_325;
  wire       [0:0]    _zz_ena_325;
  wire       [15:0]   _zz_addra_326;
  wire       [15:0]   _zz_addrb_326;
  wire       [0:0]    _zz_ena_326;
  wire       [15:0]   _zz_addra_327;
  wire       [15:0]   _zz_addrb_327;
  wire       [0:0]    _zz_ena_327;
  wire       [15:0]   _zz_addra_328;
  wire       [15:0]   _zz_addrb_328;
  wire       [0:0]    _zz_ena_328;
  wire       [15:0]   _zz_addra_329;
  wire       [15:0]   _zz_addrb_329;
  wire       [0:0]    _zz_ena_329;
  wire       [15:0]   _zz_addra_330;
  wire       [15:0]   _zz_addrb_330;
  wire       [0:0]    _zz_ena_330;
  wire       [15:0]   _zz_addra_331;
  wire       [15:0]   _zz_addrb_331;
  wire       [0:0]    _zz_ena_331;
  wire       [15:0]   _zz_addra_332;
  wire       [15:0]   _zz_addrb_332;
  wire       [0:0]    _zz_ena_332;
  wire       [15:0]   _zz_addra_333;
  wire       [15:0]   _zz_addrb_333;
  wire       [0:0]    _zz_ena_333;
  wire       [15:0]   _zz_addra_334;
  wire       [15:0]   _zz_addrb_334;
  wire       [0:0]    _zz_ena_334;
  wire       [15:0]   _zz_addra_335;
  wire       [15:0]   _zz_addrb_335;
  wire       [0:0]    _zz_ena_335;
  wire       [15:0]   _zz_addra_336;
  wire       [15:0]   _zz_addrb_336;
  wire       [0:0]    _zz_ena_336;
  wire       [15:0]   _zz_addra_337;
  wire       [15:0]   _zz_addrb_337;
  wire       [0:0]    _zz_ena_337;
  wire       [15:0]   _zz_addra_338;
  wire       [15:0]   _zz_addrb_338;
  wire       [0:0]    _zz_ena_338;
  wire       [15:0]   _zz_addra_339;
  wire       [15:0]   _zz_addrb_339;
  wire       [0:0]    _zz_ena_339;
  wire       [15:0]   _zz_addra_340;
  wire       [15:0]   _zz_addrb_340;
  wire       [0:0]    _zz_ena_340;
  wire       [15:0]   _zz_addra_341;
  wire       [15:0]   _zz_addrb_341;
  wire       [0:0]    _zz_ena_341;
  wire       [15:0]   _zz_addra_342;
  wire       [15:0]   _zz_addrb_342;
  wire       [0:0]    _zz_ena_342;
  wire       [15:0]   _zz_addra_343;
  wire       [15:0]   _zz_addrb_343;
  wire       [0:0]    _zz_ena_343;
  wire       [15:0]   _zz_addra_344;
  wire       [15:0]   _zz_addrb_344;
  wire       [0:0]    _zz_ena_344;
  wire       [15:0]   _zz_addra_345;
  wire       [15:0]   _zz_addrb_345;
  wire       [0:0]    _zz_ena_345;
  wire       [15:0]   _zz_addra_346;
  wire       [15:0]   _zz_addrb_346;
  wire       [0:0]    _zz_ena_346;
  wire       [15:0]   _zz_addra_347;
  wire       [15:0]   _zz_addrb_347;
  wire       [0:0]    _zz_ena_347;
  wire       [15:0]   _zz_addra_348;
  wire       [15:0]   _zz_addrb_348;
  wire       [0:0]    _zz_ena_348;
  wire       [15:0]   _zz_addra_349;
  wire       [15:0]   _zz_addrb_349;
  wire       [0:0]    _zz_ena_349;
  wire       [15:0]   _zz_addra_350;
  wire       [15:0]   _zz_addrb_350;
  wire       [0:0]    _zz_ena_350;
  wire       [15:0]   _zz_addra_351;
  wire       [15:0]   _zz_addrb_351;
  wire       [0:0]    _zz_ena_351;
  wire       [15:0]   _zz_addra_352;
  wire       [15:0]   _zz_addrb_352;
  wire       [0:0]    _zz_ena_352;
  wire       [15:0]   _zz_addra_353;
  wire       [15:0]   _zz_addrb_353;
  wire       [0:0]    _zz_ena_353;
  wire       [15:0]   _zz_addra_354;
  wire       [15:0]   _zz_addrb_354;
  wire       [0:0]    _zz_ena_354;
  wire       [15:0]   _zz_addra_355;
  wire       [15:0]   _zz_addrb_355;
  wire       [0:0]    _zz_ena_355;
  wire       [15:0]   _zz_addra_356;
  wire       [15:0]   _zz_addrb_356;
  wire       [0:0]    _zz_ena_356;
  wire       [15:0]   _zz_addra_357;
  wire       [15:0]   _zz_addrb_357;
  wire       [0:0]    _zz_ena_357;
  wire       [15:0]   _zz_addra_358;
  wire       [15:0]   _zz_addrb_358;
  wire       [0:0]    _zz_ena_358;
  wire       [15:0]   _zz_addra_359;
  wire       [15:0]   _zz_addrb_359;
  wire       [0:0]    _zz_ena_359;
  wire       [15:0]   _zz_addra_360;
  wire       [15:0]   _zz_addrb_360;
  wire       [0:0]    _zz_ena_360;
  wire       [15:0]   _zz_addra_361;
  wire       [15:0]   _zz_addrb_361;
  wire       [0:0]    _zz_ena_361;
  wire       [15:0]   _zz_addra_362;
  wire       [15:0]   _zz_addrb_362;
  wire       [0:0]    _zz_ena_362;
  wire       [15:0]   _zz_addra_363;
  wire       [15:0]   _zz_addrb_363;
  wire       [0:0]    _zz_ena_363;
  wire       [15:0]   _zz_addra_364;
  wire       [15:0]   _zz_addrb_364;
  wire       [0:0]    _zz_ena_364;
  wire       [15:0]   _zz_addra_365;
  wire       [15:0]   _zz_addrb_365;
  wire       [0:0]    _zz_ena_365;
  wire       [15:0]   _zz_addra_366;
  wire       [15:0]   _zz_addrb_366;
  wire       [0:0]    _zz_ena_366;
  wire       [15:0]   _zz_addra_367;
  wire       [15:0]   _zz_addrb_367;
  wire       [0:0]    _zz_ena_367;
  wire       [15:0]   _zz_addra_368;
  wire       [15:0]   _zz_addrb_368;
  wire       [0:0]    _zz_ena_368;
  wire       [15:0]   _zz_addra_369;
  wire       [15:0]   _zz_addrb_369;
  wire       [0:0]    _zz_ena_369;
  wire       [15:0]   _zz_addra_370;
  wire       [15:0]   _zz_addrb_370;
  wire       [0:0]    _zz_ena_370;
  wire       [15:0]   _zz_addra_371;
  wire       [15:0]   _zz_addrb_371;
  wire       [0:0]    _zz_ena_371;
  wire       [15:0]   _zz_addra_372;
  wire       [15:0]   _zz_addrb_372;
  wire       [0:0]    _zz_ena_372;
  wire       [15:0]   _zz_addra_373;
  wire       [15:0]   _zz_addrb_373;
  wire       [0:0]    _zz_ena_373;
  wire       [15:0]   _zz_addra_374;
  wire       [15:0]   _zz_addrb_374;
  wire       [0:0]    _zz_ena_374;
  wire       [15:0]   _zz_addra_375;
  wire       [15:0]   _zz_addrb_375;
  wire       [0:0]    _zz_ena_375;
  wire       [15:0]   _zz_addra_376;
  wire       [15:0]   _zz_addrb_376;
  wire       [0:0]    _zz_ena_376;
  wire       [15:0]   _zz_addra_377;
  wire       [15:0]   _zz_addrb_377;
  wire       [0:0]    _zz_ena_377;
  wire       [15:0]   _zz_addra_378;
  wire       [15:0]   _zz_addrb_378;
  wire       [0:0]    _zz_ena_378;
  wire       [15:0]   _zz_addra_379;
  wire       [15:0]   _zz_addrb_379;
  wire       [0:0]    _zz_ena_379;
  wire       [15:0]   _zz_addra_380;
  wire       [15:0]   _zz_addrb_380;
  wire       [0:0]    _zz_ena_380;
  wire       [15:0]   _zz_addra_381;
  wire       [15:0]   _zz_addrb_381;
  wire       [0:0]    _zz_ena_381;
  wire       [15:0]   _zz_addra_382;
  wire       [15:0]   _zz_addrb_382;
  wire       [0:0]    _zz_ena_382;
  wire       [15:0]   _zz_addra_383;
  wire       [15:0]   _zz_addrb_383;
  wire       [0:0]    _zz_ena_383;
  wire       [15:0]   _zz_addra_384;
  wire       [15:0]   _zz_addrb_384;
  wire       [0:0]    _zz_ena_384;
  wire       [15:0]   _zz_addra_385;
  wire       [15:0]   _zz_addrb_385;
  wire       [0:0]    _zz_ena_385;
  wire       [15:0]   _zz_addra_386;
  wire       [15:0]   _zz_addrb_386;
  wire       [0:0]    _zz_ena_386;
  wire       [15:0]   _zz_addra_387;
  wire       [15:0]   _zz_addrb_387;
  wire       [0:0]    _zz_ena_387;
  wire       [15:0]   _zz_addra_388;
  wire       [15:0]   _zz_addrb_388;
  wire       [0:0]    _zz_ena_388;
  wire       [15:0]   _zz_addra_389;
  wire       [15:0]   _zz_addrb_389;
  wire       [0:0]    _zz_ena_389;
  wire       [15:0]   _zz_addra_390;
  wire       [15:0]   _zz_addrb_390;
  wire       [0:0]    _zz_ena_390;
  wire       [15:0]   _zz_addra_391;
  wire       [15:0]   _zz_addrb_391;
  wire       [0:0]    _zz_ena_391;
  wire       [15:0]   _zz_addra_392;
  wire       [15:0]   _zz_addrb_392;
  wire       [0:0]    _zz_ena_392;
  wire       [15:0]   _zz_addra_393;
  wire       [15:0]   _zz_addrb_393;
  wire       [0:0]    _zz_ena_393;
  wire       [15:0]   _zz_addra_394;
  wire       [15:0]   _zz_addrb_394;
  wire       [0:0]    _zz_ena_394;
  wire       [15:0]   _zz_addra_395;
  wire       [15:0]   _zz_addrb_395;
  wire       [0:0]    _zz_ena_395;
  wire       [15:0]   _zz_addra_396;
  wire       [15:0]   _zz_addrb_396;
  wire       [0:0]    _zz_ena_396;
  wire       [15:0]   _zz_addra_397;
  wire       [15:0]   _zz_addrb_397;
  wire       [0:0]    _zz_ena_397;
  wire       [15:0]   _zz_addra_398;
  wire       [15:0]   _zz_addrb_398;
  wire       [0:0]    _zz_ena_398;
  wire       [15:0]   _zz_addra_399;
  wire       [15:0]   _zz_addrb_399;
  wire       [0:0]    _zz_ena_399;
  wire       [15:0]   _zz_addra_400;
  wire       [15:0]   _zz_addrb_400;
  wire       [0:0]    _zz_ena_400;
  wire       [15:0]   _zz_addra_401;
  wire       [15:0]   _zz_addrb_401;
  wire       [0:0]    _zz_ena_401;
  wire       [15:0]   _zz_addra_402;
  wire       [15:0]   _zz_addrb_402;
  wire       [0:0]    _zz_ena_402;
  wire       [15:0]   _zz_addra_403;
  wire       [15:0]   _zz_addrb_403;
  wire       [0:0]    _zz_ena_403;
  wire       [15:0]   _zz_addra_404;
  wire       [15:0]   _zz_addrb_404;
  wire       [0:0]    _zz_ena_404;
  wire       [15:0]   _zz_addra_405;
  wire       [15:0]   _zz_addrb_405;
  wire       [0:0]    _zz_ena_405;
  wire       [15:0]   _zz_addra_406;
  wire       [15:0]   _zz_addrb_406;
  wire       [0:0]    _zz_ena_406;
  wire       [15:0]   _zz_addra_407;
  wire       [15:0]   _zz_addrb_407;
  wire       [0:0]    _zz_ena_407;
  wire       [15:0]   _zz_addra_408;
  wire       [15:0]   _zz_addrb_408;
  wire       [0:0]    _zz_ena_408;
  wire       [15:0]   _zz_addra_409;
  wire       [15:0]   _zz_addrb_409;
  wire       [0:0]    _zz_ena_409;
  wire       [15:0]   _zz_addra_410;
  wire       [15:0]   _zz_addrb_410;
  wire       [0:0]    _zz_ena_410;
  wire       [15:0]   _zz_addra_411;
  wire       [15:0]   _zz_addrb_411;
  wire       [0:0]    _zz_ena_411;
  wire       [15:0]   _zz_addra_412;
  wire       [15:0]   _zz_addrb_412;
  wire       [0:0]    _zz_ena_412;
  wire       [15:0]   _zz_addra_413;
  wire       [15:0]   _zz_addrb_413;
  wire       [0:0]    _zz_ena_413;
  wire       [15:0]   _zz_addra_414;
  wire       [15:0]   _zz_addrb_414;
  wire       [0:0]    _zz_ena_414;
  wire       [15:0]   _zz_addra_415;
  wire       [15:0]   _zz_addrb_415;
  wire       [0:0]    _zz_ena_415;
  wire       [15:0]   _zz_addra_416;
  wire       [15:0]   _zz_addrb_416;
  wire       [0:0]    _zz_ena_416;
  wire       [15:0]   _zz_addra_417;
  wire       [15:0]   _zz_addrb_417;
  wire       [0:0]    _zz_ena_417;
  wire       [15:0]   _zz_addra_418;
  wire       [15:0]   _zz_addrb_418;
  wire       [0:0]    _zz_ena_418;
  wire       [15:0]   _zz_addra_419;
  wire       [15:0]   _zz_addrb_419;
  wire       [0:0]    _zz_ena_419;
  wire       [15:0]   _zz_addra_420;
  wire       [15:0]   _zz_addrb_420;
  wire       [0:0]    _zz_ena_420;
  wire       [15:0]   _zz_addra_421;
  wire       [15:0]   _zz_addrb_421;
  wire       [0:0]    _zz_ena_421;
  wire       [15:0]   _zz_addra_422;
  wire       [15:0]   _zz_addrb_422;
  wire       [0:0]    _zz_ena_422;
  wire       [15:0]   _zz_addra_423;
  wire       [15:0]   _zz_addrb_423;
  wire       [0:0]    _zz_ena_423;
  wire       [15:0]   _zz_addra_424;
  wire       [15:0]   _zz_addrb_424;
  wire       [0:0]    _zz_ena_424;
  wire       [15:0]   _zz_addra_425;
  wire       [15:0]   _zz_addrb_425;
  wire       [0:0]    _zz_ena_425;
  wire       [15:0]   _zz_addra_426;
  wire       [15:0]   _zz_addrb_426;
  wire       [0:0]    _zz_ena_426;
  wire       [15:0]   _zz_addra_427;
  wire       [15:0]   _zz_addrb_427;
  wire       [0:0]    _zz_ena_427;
  wire       [15:0]   _zz_addra_428;
  wire       [15:0]   _zz_addrb_428;
  wire       [0:0]    _zz_ena_428;
  wire       [15:0]   _zz_addra_429;
  wire       [15:0]   _zz_addrb_429;
  wire       [0:0]    _zz_ena_429;
  wire       [15:0]   _zz_addra_430;
  wire       [15:0]   _zz_addrb_430;
  wire       [0:0]    _zz_ena_430;
  wire       [15:0]   _zz_addra_431;
  wire       [15:0]   _zz_addrb_431;
  wire       [0:0]    _zz_ena_431;
  wire       [15:0]   _zz_addra_432;
  wire       [15:0]   _zz_addrb_432;
  wire       [0:0]    _zz_ena_432;
  wire       [15:0]   _zz_addra_433;
  wire       [15:0]   _zz_addrb_433;
  wire       [0:0]    _zz_ena_433;
  wire       [15:0]   _zz_addra_434;
  wire       [15:0]   _zz_addrb_434;
  wire       [0:0]    _zz_ena_434;
  wire       [15:0]   _zz_addra_435;
  wire       [15:0]   _zz_addrb_435;
  wire       [0:0]    _zz_ena_435;
  wire       [15:0]   _zz_addra_436;
  wire       [15:0]   _zz_addrb_436;
  wire       [0:0]    _zz_ena_436;
  wire       [15:0]   _zz_addra_437;
  wire       [15:0]   _zz_addrb_437;
  wire       [0:0]    _zz_ena_437;
  wire       [15:0]   _zz_addra_438;
  wire       [15:0]   _zz_addrb_438;
  wire       [0:0]    _zz_ena_438;
  wire       [15:0]   _zz_addra_439;
  wire       [15:0]   _zz_addrb_439;
  wire       [0:0]    _zz_ena_439;
  wire       [15:0]   _zz_addra_440;
  wire       [15:0]   _zz_addrb_440;
  wire       [0:0]    _zz_ena_440;
  wire       [15:0]   _zz_addra_441;
  wire       [15:0]   _zz_addrb_441;
  wire       [0:0]    _zz_ena_441;
  wire       [15:0]   _zz_addra_442;
  wire       [15:0]   _zz_addrb_442;
  wire       [0:0]    _zz_ena_442;
  wire       [15:0]   _zz_addra_443;
  wire       [15:0]   _zz_addrb_443;
  wire       [0:0]    _zz_ena_443;
  wire       [15:0]   _zz_addra_444;
  wire       [15:0]   _zz_addrb_444;
  wire       [0:0]    _zz_ena_444;
  wire       [15:0]   _zz_addra_445;
  wire       [15:0]   _zz_addrb_445;
  wire       [0:0]    _zz_ena_445;
  wire       [15:0]   _zz_addra_446;
  wire       [15:0]   _zz_addrb_446;
  wire       [0:0]    _zz_ena_446;
  wire       [15:0]   _zz_addra_447;
  wire       [15:0]   _zz_addrb_447;
  wire       [0:0]    _zz_ena_447;
  wire       [15:0]   _zz_addra_448;
  wire       [15:0]   _zz_addrb_448;
  wire       [0:0]    _zz_ena_448;
  wire       [15:0]   _zz_addra_449;
  wire       [15:0]   _zz_addrb_449;
  wire       [0:0]    _zz_ena_449;
  wire       [15:0]   _zz_addra_450;
  wire       [15:0]   _zz_addrb_450;
  wire       [0:0]    _zz_ena_450;
  wire       [15:0]   _zz_addra_451;
  wire       [15:0]   _zz_addrb_451;
  wire       [0:0]    _zz_ena_451;
  wire       [15:0]   _zz_addra_452;
  wire       [15:0]   _zz_addrb_452;
  wire       [0:0]    _zz_ena_452;
  wire       [15:0]   _zz_addra_453;
  wire       [15:0]   _zz_addrb_453;
  wire       [0:0]    _zz_ena_453;
  wire       [15:0]   _zz_addra_454;
  wire       [15:0]   _zz_addrb_454;
  wire       [0:0]    _zz_ena_454;
  wire       [15:0]   _zz_addra_455;
  wire       [15:0]   _zz_addrb_455;
  wire       [0:0]    _zz_ena_455;
  wire       [15:0]   _zz_addra_456;
  wire       [15:0]   _zz_addrb_456;
  wire       [0:0]    _zz_ena_456;
  wire       [15:0]   _zz_addra_457;
  wire       [15:0]   _zz_addrb_457;
  wire       [0:0]    _zz_ena_457;
  wire       [15:0]   _zz_addra_458;
  wire       [15:0]   _zz_addrb_458;
  wire       [0:0]    _zz_ena_458;
  wire       [15:0]   _zz_addra_459;
  wire       [15:0]   _zz_addrb_459;
  wire       [0:0]    _zz_ena_459;
  wire       [15:0]   _zz_addra_460;
  wire       [15:0]   _zz_addrb_460;
  wire       [0:0]    _zz_ena_460;
  wire       [15:0]   _zz_addra_461;
  wire       [15:0]   _zz_addrb_461;
  wire       [0:0]    _zz_ena_461;
  wire       [15:0]   _zz_addra_462;
  wire       [15:0]   _zz_addrb_462;
  wire       [0:0]    _zz_ena_462;
  wire       [15:0]   _zz_addra_463;
  wire       [15:0]   _zz_addrb_463;
  wire       [0:0]    _zz_ena_463;
  wire       [15:0]   _zz_addra_464;
  wire       [15:0]   _zz_addrb_464;
  wire       [0:0]    _zz_ena_464;
  wire       [15:0]   _zz_addra_465;
  wire       [15:0]   _zz_addrb_465;
  wire       [0:0]    _zz_ena_465;
  wire       [15:0]   _zz_addra_466;
  wire       [15:0]   _zz_addrb_466;
  wire       [0:0]    _zz_ena_466;
  wire       [15:0]   _zz_addra_467;
  wire       [15:0]   _zz_addrb_467;
  wire       [0:0]    _zz_ena_467;
  wire       [15:0]   _zz_addra_468;
  wire       [15:0]   _zz_addrb_468;
  wire       [0:0]    _zz_ena_468;
  wire       [15:0]   _zz_addra_469;
  wire       [15:0]   _zz_addrb_469;
  wire       [0:0]    _zz_ena_469;
  wire       [15:0]   _zz_addra_470;
  wire       [15:0]   _zz_addrb_470;
  wire       [0:0]    _zz_ena_470;
  wire       [15:0]   _zz_addra_471;
  wire       [15:0]   _zz_addrb_471;
  wire       [0:0]    _zz_ena_471;
  wire       [15:0]   _zz_addra_472;
  wire       [15:0]   _zz_addrb_472;
  wire       [0:0]    _zz_ena_472;
  wire       [15:0]   _zz_addra_473;
  wire       [15:0]   _zz_addrb_473;
  wire       [0:0]    _zz_ena_473;
  wire       [15:0]   _zz_addra_474;
  wire       [15:0]   _zz_addrb_474;
  wire       [0:0]    _zz_ena_474;
  wire       [15:0]   _zz_addra_475;
  wire       [15:0]   _zz_addrb_475;
  wire       [0:0]    _zz_ena_475;
  wire       [15:0]   _zz_addra_476;
  wire       [15:0]   _zz_addrb_476;
  wire       [0:0]    _zz_ena_476;
  wire       [15:0]   _zz_addra_477;
  wire       [15:0]   _zz_addrb_477;
  wire       [0:0]    _zz_ena_477;
  wire       [15:0]   _zz_addra_478;
  wire       [15:0]   _zz_addrb_478;
  wire       [0:0]    _zz_ena_478;
  wire       [15:0]   _zz_addra_479;
  wire       [15:0]   _zz_addrb_479;
  wire       [0:0]    _zz_ena_479;
  wire       [15:0]   _zz_addra_480;
  wire       [15:0]   _zz_addrb_480;
  wire       [0:0]    _zz_ena_480;
  wire       [15:0]   _zz_addra_481;
  wire       [15:0]   _zz_addrb_481;
  wire       [0:0]    _zz_ena_481;
  wire       [15:0]   _zz_addra_482;
  wire       [15:0]   _zz_addrb_482;
  wire       [0:0]    _zz_ena_482;
  wire       [15:0]   _zz_addra_483;
  wire       [15:0]   _zz_addrb_483;
  wire       [0:0]    _zz_ena_483;
  wire       [15:0]   _zz_addra_484;
  wire       [15:0]   _zz_addrb_484;
  wire       [0:0]    _zz_ena_484;
  wire       [15:0]   _zz_addra_485;
  wire       [15:0]   _zz_addrb_485;
  wire       [0:0]    _zz_ena_485;
  wire       [15:0]   _zz_addra_486;
  wire       [15:0]   _zz_addrb_486;
  wire       [0:0]    _zz_ena_486;
  wire       [15:0]   _zz_addra_487;
  wire       [15:0]   _zz_addrb_487;
  wire       [0:0]    _zz_ena_487;
  wire       [15:0]   _zz_addra_488;
  wire       [15:0]   _zz_addrb_488;
  wire       [0:0]    _zz_ena_488;
  wire       [15:0]   _zz_addra_489;
  wire       [15:0]   _zz_addrb_489;
  wire       [0:0]    _zz_ena_489;
  wire       [15:0]   _zz_addra_490;
  wire       [15:0]   _zz_addrb_490;
  wire       [0:0]    _zz_ena_490;
  wire       [15:0]   _zz_addra_491;
  wire       [15:0]   _zz_addrb_491;
  wire       [0:0]    _zz_ena_491;
  wire       [15:0]   _zz_addra_492;
  wire       [15:0]   _zz_addrb_492;
  wire       [0:0]    _zz_ena_492;
  wire       [15:0]   _zz_addra_493;
  wire       [15:0]   _zz_addrb_493;
  wire       [0:0]    _zz_ena_493;
  wire       [15:0]   _zz_addra_494;
  wire       [15:0]   _zz_addrb_494;
  wire       [0:0]    _zz_ena_494;
  wire       [15:0]   _zz_addra_495;
  wire       [15:0]   _zz_addrb_495;
  wire       [0:0]    _zz_ena_495;
  wire       [15:0]   _zz_addra_496;
  wire       [15:0]   _zz_addrb_496;
  wire       [0:0]    _zz_ena_496;
  wire       [15:0]   _zz_addra_497;
  wire       [15:0]   _zz_addrb_497;
  wire       [0:0]    _zz_ena_497;
  wire       [15:0]   _zz_addra_498;
  wire       [15:0]   _zz_addrb_498;
  wire       [0:0]    _zz_ena_498;
  wire       [15:0]   _zz_addra_499;
  wire       [15:0]   _zz_addrb_499;
  wire       [0:0]    _zz_ena_499;
  wire       [15:0]   _zz_addra_500;
  wire       [15:0]   _zz_addrb_500;
  wire       [0:0]    _zz_ena_500;
  wire       [15:0]   _zz_addra_501;
  wire       [15:0]   _zz_addrb_501;
  wire       [0:0]    _zz_ena_501;
  wire       [15:0]   _zz_addra_502;
  wire       [15:0]   _zz_addrb_502;
  wire       [0:0]    _zz_ena_502;
  wire       [15:0]   _zz_addra_503;
  wire       [15:0]   _zz_addrb_503;
  wire       [0:0]    _zz_ena_503;
  wire       [15:0]   _zz_addra_504;
  wire       [15:0]   _zz_addrb_504;
  wire       [0:0]    _zz_ena_504;
  wire       [15:0]   _zz_addra_505;
  wire       [15:0]   _zz_addrb_505;
  wire       [0:0]    _zz_ena_505;
  wire       [15:0]   _zz_addra_506;
  wire       [15:0]   _zz_addrb_506;
  wire       [0:0]    _zz_ena_506;
  wire       [15:0]   _zz_addra_507;
  wire       [15:0]   _zz_addrb_507;
  wire       [0:0]    _zz_ena_507;
  wire       [15:0]   _zz_addra_508;
  wire       [15:0]   _zz_addrb_508;
  wire       [0:0]    _zz_ena_508;
  wire       [15:0]   _zz_addra_509;
  wire       [15:0]   _zz_addrb_509;
  wire       [0:0]    _zz_ena_509;
  wire       [15:0]   _zz_addra_510;
  wire       [15:0]   _zz_addrb_510;
  wire       [0:0]    _zz_ena_510;
  wire       [15:0]   _zz_addra_511;
  wire       [15:0]   _zz_addrb_511;
  wire       [0:0]    _zz_ena_511;
  reg                 start_regNext;
  wire                when_SA3D_WeightCache_l33;
  reg        [3:0]    Fsm_currentState;
  reg        [3:0]    Fsm_nextState;
  wire                Fsm_Init_End;
  wire                Fsm_Weight_All_Cached;
  wire                Fsm_SA_Computed;
  wire                when_WaCounter_l19;
  reg        [2:0]    Init_Count_count;
  reg                 Init_Count_valid;
  wire                when_WaCounter_l14;
  reg        [511:0]  InData_Switch;
  wire       [12:0]   Matrix_In_MaxCnt;
  wire                sData_fire;
  reg        [15:0]   In_Row_Cnt_count;
  wire                In_Row_Cnt_valid;
  reg        [15:0]   In_Col_Cnt_count;
  wire                In_Col_Cnt_valid;
  reg        [15:0]   Read_Row_Base_Addr;
  reg        [15:0]   Write_Row_Base_Addr;
  wire                when_WaCounter_l40;
  reg        [15:0]   OutRow_Cnt_count;
  wire                OutRow_Cnt_valid;
  wire       [3:0]    _zz_OutCol_Cnt_count;
  reg        [15:0]   OutCol_Cnt_count;
  reg                 OutCol_Cnt_valid;
  reg        [8:0]    Col_In_8_Cnt_count;
  reg                 Col_In_8_Cnt_valid;
  wire                when_SA3D_WeightCache_l129;
  wire                when_SA3D_WeightCache_l134;
  wire                sData_fire_1;
  wire                sData_fire_2;
  wire                sData_fire_3;
  wire                sData_fire_4;
  wire                sData_fire_5;
  wire                sData_fire_6;
  wire                sData_fire_7;
  wire                sData_fire_8;
  wire                sData_fire_9;
  wire                sData_fire_10;
  wire                sData_fire_11;
  wire                sData_fire_12;
  wire                sData_fire_13;
  wire                sData_fire_14;
  wire                sData_fire_15;
  wire                sData_fire_16;
  wire                sData_fire_17;
  wire                sData_fire_18;
  wire                sData_fire_19;
  wire                sData_fire_20;
  wire                sData_fire_21;
  wire                sData_fire_22;
  wire                sData_fire_23;
  wire                sData_fire_24;
  wire                sData_fire_25;
  wire                sData_fire_26;
  wire                sData_fire_27;
  wire                sData_fire_28;
  wire                sData_fire_29;
  wire                sData_fire_30;
  wire                sData_fire_31;
  wire                sData_fire_32;
  wire                sData_fire_33;
  wire                sData_fire_34;
  wire                sData_fire_35;
  wire                sData_fire_36;
  wire                sData_fire_37;
  wire                sData_fire_38;
  wire                sData_fire_39;
  wire                sData_fire_40;
  wire                sData_fire_41;
  wire                sData_fire_42;
  wire                sData_fire_43;
  wire                sData_fire_44;
  wire                sData_fire_45;
  wire                sData_fire_46;
  wire                sData_fire_47;
  wire                sData_fire_48;
  wire                sData_fire_49;
  wire                sData_fire_50;
  wire                sData_fire_51;
  wire                sData_fire_52;
  wire                sData_fire_53;
  wire                sData_fire_54;
  wire                sData_fire_55;
  wire                sData_fire_56;
  wire                sData_fire_57;
  wire                sData_fire_58;
  wire                sData_fire_59;
  wire                sData_fire_60;
  wire                sData_fire_61;
  wire                sData_fire_62;
  wire                sData_fire_63;
  wire                sData_fire_64;
  wire                sData_fire_65;
  wire                sData_fire_66;
  wire                sData_fire_67;
  wire                sData_fire_68;
  wire                sData_fire_69;
  wire                sData_fire_70;
  wire                sData_fire_71;
  wire                sData_fire_72;
  wire                sData_fire_73;
  wire                sData_fire_74;
  wire                sData_fire_75;
  wire                sData_fire_76;
  wire                sData_fire_77;
  wire                sData_fire_78;
  wire                sData_fire_79;
  wire                sData_fire_80;
  wire                sData_fire_81;
  wire                sData_fire_82;
  wire                sData_fire_83;
  wire                sData_fire_84;
  wire                sData_fire_85;
  wire                sData_fire_86;
  wire                sData_fire_87;
  wire                sData_fire_88;
  wire                sData_fire_89;
  wire                sData_fire_90;
  wire                sData_fire_91;
  wire                sData_fire_92;
  wire                sData_fire_93;
  wire                sData_fire_94;
  wire                sData_fire_95;
  wire                sData_fire_96;
  wire                sData_fire_97;
  wire                sData_fire_98;
  wire                sData_fire_99;
  wire                sData_fire_100;
  wire                sData_fire_101;
  wire                sData_fire_102;
  wire                sData_fire_103;
  wire                sData_fire_104;
  wire                sData_fire_105;
  wire                sData_fire_106;
  wire                sData_fire_107;
  wire                sData_fire_108;
  wire                sData_fire_109;
  wire                sData_fire_110;
  wire                sData_fire_111;
  wire                sData_fire_112;
  wire                sData_fire_113;
  wire                sData_fire_114;
  wire                sData_fire_115;
  wire                sData_fire_116;
  wire                sData_fire_117;
  wire                sData_fire_118;
  wire                sData_fire_119;
  wire                sData_fire_120;
  wire                sData_fire_121;
  wire                sData_fire_122;
  wire                sData_fire_123;
  wire                sData_fire_124;
  wire                sData_fire_125;
  wire                sData_fire_126;
  wire                sData_fire_127;
  wire                sData_fire_128;
  wire                sData_fire_129;
  wire                sData_fire_130;
  wire                sData_fire_131;
  wire                sData_fire_132;
  wire                sData_fire_133;
  wire                sData_fire_134;
  wire                sData_fire_135;
  wire                sData_fire_136;
  wire                sData_fire_137;
  wire                sData_fire_138;
  wire                sData_fire_139;
  wire                sData_fire_140;
  wire                sData_fire_141;
  wire                sData_fire_142;
  wire                sData_fire_143;
  wire                sData_fire_144;
  wire                sData_fire_145;
  wire                sData_fire_146;
  wire                sData_fire_147;
  wire                sData_fire_148;
  wire                sData_fire_149;
  wire                sData_fire_150;
  wire                sData_fire_151;
  wire                sData_fire_152;
  wire                sData_fire_153;
  wire                sData_fire_154;
  wire                sData_fire_155;
  wire                sData_fire_156;
  wire                sData_fire_157;
  wire                sData_fire_158;
  wire                sData_fire_159;
  wire                sData_fire_160;
  wire                sData_fire_161;
  wire                sData_fire_162;
  wire                sData_fire_163;
  wire                sData_fire_164;
  wire                sData_fire_165;
  wire                sData_fire_166;
  wire                sData_fire_167;
  wire                sData_fire_168;
  wire                sData_fire_169;
  wire                sData_fire_170;
  wire                sData_fire_171;
  wire                sData_fire_172;
  wire                sData_fire_173;
  wire                sData_fire_174;
  wire                sData_fire_175;
  wire                sData_fire_176;
  wire                sData_fire_177;
  wire                sData_fire_178;
  wire                sData_fire_179;
  wire                sData_fire_180;
  wire                sData_fire_181;
  wire                sData_fire_182;
  wire                sData_fire_183;
  wire                sData_fire_184;
  wire                sData_fire_185;
  wire                sData_fire_186;
  wire                sData_fire_187;
  wire                sData_fire_188;
  wire                sData_fire_189;
  wire                sData_fire_190;
  wire                sData_fire_191;
  wire                sData_fire_192;
  wire                sData_fire_193;
  wire                sData_fire_194;
  wire                sData_fire_195;
  wire                sData_fire_196;
  wire                sData_fire_197;
  wire                sData_fire_198;
  wire                sData_fire_199;
  wire                sData_fire_200;
  wire                sData_fire_201;
  wire                sData_fire_202;
  wire                sData_fire_203;
  wire                sData_fire_204;
  wire                sData_fire_205;
  wire                sData_fire_206;
  wire                sData_fire_207;
  wire                sData_fire_208;
  wire                sData_fire_209;
  wire                sData_fire_210;
  wire                sData_fire_211;
  wire                sData_fire_212;
  wire                sData_fire_213;
  wire                sData_fire_214;
  wire                sData_fire_215;
  wire                sData_fire_216;
  wire                sData_fire_217;
  wire                sData_fire_218;
  wire                sData_fire_219;
  wire                sData_fire_220;
  wire                sData_fire_221;
  wire                sData_fire_222;
  wire                sData_fire_223;
  wire                sData_fire_224;
  wire                sData_fire_225;
  wire                sData_fire_226;
  wire                sData_fire_227;
  wire                sData_fire_228;
  wire                sData_fire_229;
  wire                sData_fire_230;
  wire                sData_fire_231;
  wire                sData_fire_232;
  wire                sData_fire_233;
  wire                sData_fire_234;
  wire                sData_fire_235;
  wire                sData_fire_236;
  wire                sData_fire_237;
  wire                sData_fire_238;
  wire                sData_fire_239;
  wire                sData_fire_240;
  wire                sData_fire_241;
  wire                sData_fire_242;
  wire                sData_fire_243;
  wire                sData_fire_244;
  wire                sData_fire_245;
  wire                sData_fire_246;
  wire                sData_fire_247;
  wire                sData_fire_248;
  wire                sData_fire_249;
  wire                sData_fire_250;
  wire                sData_fire_251;
  wire                sData_fire_252;
  wire                sData_fire_253;
  wire                sData_fire_254;
  wire                sData_fire_255;
  wire                sData_fire_256;
  wire                sData_fire_257;
  wire                sData_fire_258;
  wire                sData_fire_259;
  wire                sData_fire_260;
  wire                sData_fire_261;
  wire                sData_fire_262;
  wire                sData_fire_263;
  wire                sData_fire_264;
  wire                sData_fire_265;
  wire                sData_fire_266;
  wire                sData_fire_267;
  wire                sData_fire_268;
  wire                sData_fire_269;
  wire                sData_fire_270;
  wire                sData_fire_271;
  wire                sData_fire_272;
  wire                sData_fire_273;
  wire                sData_fire_274;
  wire                sData_fire_275;
  wire                sData_fire_276;
  wire                sData_fire_277;
  wire                sData_fire_278;
  wire                sData_fire_279;
  wire                sData_fire_280;
  wire                sData_fire_281;
  wire                sData_fire_282;
  wire                sData_fire_283;
  wire                sData_fire_284;
  wire                sData_fire_285;
  wire                sData_fire_286;
  wire                sData_fire_287;
  wire                sData_fire_288;
  wire                sData_fire_289;
  wire                sData_fire_290;
  wire                sData_fire_291;
  wire                sData_fire_292;
  wire                sData_fire_293;
  wire                sData_fire_294;
  wire                sData_fire_295;
  wire                sData_fire_296;
  wire                sData_fire_297;
  wire                sData_fire_298;
  wire                sData_fire_299;
  wire                sData_fire_300;
  wire                sData_fire_301;
  wire                sData_fire_302;
  wire                sData_fire_303;
  wire                sData_fire_304;
  wire                sData_fire_305;
  wire                sData_fire_306;
  wire                sData_fire_307;
  wire                sData_fire_308;
  wire                sData_fire_309;
  wire                sData_fire_310;
  wire                sData_fire_311;
  wire                sData_fire_312;
  wire                sData_fire_313;
  wire                sData_fire_314;
  wire                sData_fire_315;
  wire                sData_fire_316;
  wire                sData_fire_317;
  wire                sData_fire_318;
  wire                sData_fire_319;
  wire                sData_fire_320;
  wire                sData_fire_321;
  wire                sData_fire_322;
  wire                sData_fire_323;
  wire                sData_fire_324;
  wire                sData_fire_325;
  wire                sData_fire_326;
  wire                sData_fire_327;
  wire                sData_fire_328;
  wire                sData_fire_329;
  wire                sData_fire_330;
  wire                sData_fire_331;
  wire                sData_fire_332;
  wire                sData_fire_333;
  wire                sData_fire_334;
  wire                sData_fire_335;
  wire                sData_fire_336;
  wire                sData_fire_337;
  wire                sData_fire_338;
  wire                sData_fire_339;
  wire                sData_fire_340;
  wire                sData_fire_341;
  wire                sData_fire_342;
  wire                sData_fire_343;
  wire                sData_fire_344;
  wire                sData_fire_345;
  wire                sData_fire_346;
  wire                sData_fire_347;
  wire                sData_fire_348;
  wire                sData_fire_349;
  wire                sData_fire_350;
  wire                sData_fire_351;
  wire                sData_fire_352;
  wire                sData_fire_353;
  wire                sData_fire_354;
  wire                sData_fire_355;
  wire                sData_fire_356;
  wire                sData_fire_357;
  wire                sData_fire_358;
  wire                sData_fire_359;
  wire                sData_fire_360;
  wire                sData_fire_361;
  wire                sData_fire_362;
  wire                sData_fire_363;
  wire                sData_fire_364;
  wire                sData_fire_365;
  wire                sData_fire_366;
  wire                sData_fire_367;
  wire                sData_fire_368;
  wire                sData_fire_369;
  wire                sData_fire_370;
  wire                sData_fire_371;
  wire                sData_fire_372;
  wire                sData_fire_373;
  wire                sData_fire_374;
  wire                sData_fire_375;
  wire                sData_fire_376;
  wire                sData_fire_377;
  wire                sData_fire_378;
  wire                sData_fire_379;
  wire                sData_fire_380;
  wire                sData_fire_381;
  wire                sData_fire_382;
  wire                sData_fire_383;
  wire                sData_fire_384;
  wire                sData_fire_385;
  wire                sData_fire_386;
  wire                sData_fire_387;
  wire                sData_fire_388;
  wire                sData_fire_389;
  wire                sData_fire_390;
  wire                sData_fire_391;
  wire                sData_fire_392;
  wire                sData_fire_393;
  wire                sData_fire_394;
  wire                sData_fire_395;
  wire                sData_fire_396;
  wire                sData_fire_397;
  wire                sData_fire_398;
  wire                sData_fire_399;
  wire                sData_fire_400;
  wire                sData_fire_401;
  wire                sData_fire_402;
  wire                sData_fire_403;
  wire                sData_fire_404;
  wire                sData_fire_405;
  wire                sData_fire_406;
  wire                sData_fire_407;
  wire                sData_fire_408;
  wire                sData_fire_409;
  wire                sData_fire_410;
  wire                sData_fire_411;
  wire                sData_fire_412;
  wire                sData_fire_413;
  wire                sData_fire_414;
  wire                sData_fire_415;
  wire                sData_fire_416;
  wire                sData_fire_417;
  wire                sData_fire_418;
  wire                sData_fire_419;
  wire                sData_fire_420;
  wire                sData_fire_421;
  wire                sData_fire_422;
  wire                sData_fire_423;
  wire                sData_fire_424;
  wire                sData_fire_425;
  wire                sData_fire_426;
  wire                sData_fire_427;
  wire                sData_fire_428;
  wire                sData_fire_429;
  wire                sData_fire_430;
  wire                sData_fire_431;
  wire                sData_fire_432;
  wire                sData_fire_433;
  wire                sData_fire_434;
  wire                sData_fire_435;
  wire                sData_fire_436;
  wire                sData_fire_437;
  wire                sData_fire_438;
  wire                sData_fire_439;
  wire                sData_fire_440;
  wire                sData_fire_441;
  wire                sData_fire_442;
  wire                sData_fire_443;
  wire                sData_fire_444;
  wire                sData_fire_445;
  wire                sData_fire_446;
  wire                sData_fire_447;
  wire                sData_fire_448;
  wire                sData_fire_449;
  wire                sData_fire_450;
  wire                sData_fire_451;
  wire                sData_fire_452;
  wire                sData_fire_453;
  wire                sData_fire_454;
  wire                sData_fire_455;
  wire                sData_fire_456;
  wire                sData_fire_457;
  wire                sData_fire_458;
  wire                sData_fire_459;
  wire                sData_fire_460;
  wire                sData_fire_461;
  wire                sData_fire_462;
  wire                sData_fire_463;
  wire                sData_fire_464;
  wire                sData_fire_465;
  wire                sData_fire_466;
  wire                sData_fire_467;
  wire                sData_fire_468;
  wire                sData_fire_469;
  wire                sData_fire_470;
  wire                sData_fire_471;
  wire                sData_fire_472;
  wire                sData_fire_473;
  wire                sData_fire_474;
  wire                sData_fire_475;
  wire                sData_fire_476;
  wire                sData_fire_477;
  wire                sData_fire_478;
  wire                sData_fire_479;
  wire                sData_fire_480;
  wire                sData_fire_481;
  wire                sData_fire_482;
  wire                sData_fire_483;
  wire                sData_fire_484;
  wire                sData_fire_485;
  wire                sData_fire_486;
  wire                sData_fire_487;
  wire                sData_fire_488;
  wire                sData_fire_489;
  wire                sData_fire_490;
  wire                sData_fire_491;
  wire                sData_fire_492;
  wire                sData_fire_493;
  wire                sData_fire_494;
  wire                sData_fire_495;
  wire                sData_fire_496;
  wire                sData_fire_497;
  wire                sData_fire_498;
  wire                sData_fire_499;
  wire                sData_fire_500;
  wire                sData_fire_501;
  wire                sData_fire_502;
  wire                sData_fire_503;
  wire                sData_fire_504;
  wire                sData_fire_505;
  wire                sData_fire_506;
  wire                sData_fire_507;
  wire                sData_fire_508;
  wire                sData_fire_509;
  wire                sData_fire_510;
  wire                sData_fire_511;
  wire                sData_fire_512;
  reg        [7:0]    MatrixCol_Switch_1;
  reg        [7:0]    MatrixCol_Switch_1_regNext;
  `ifndef SYNTHESIS
  reg [95:0] Fsm_currentState_string;
  reg [95:0] Fsm_nextState_string;
  `endif


  assign _zz_In_Row_Cnt_valid_1 = (Matrix_In_MaxCnt - 13'h0001);
  assign _zz_In_Row_Cnt_valid = {3'd0, _zz_In_Row_Cnt_valid_1};
  assign _zz_In_Col_Cnt_valid = (Matrix_Col - 16'h0001);
  assign _zz_OutRow_Cnt_valid = (Matrix_Row - 16'h0001);
  assign _zz_OutCol_Cnt_valid = {12'd0, _zz_OutCol_Cnt_count};
  assign _zz_OutCol_Cnt_count_1 = {12'd0, _zz_OutCol_Cnt_count};
  assign _zz_Write_Row_Base_Addr = {3'd0, Matrix_In_MaxCnt};
  assign _zz_addra = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena = InData_Switch[0 : 0];
  assign _zz_addra_1 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_1 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_1 = InData_Switch[1 : 1];
  assign _zz_addra_2 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_2 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_2 = InData_Switch[2 : 2];
  assign _zz_addra_3 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_3 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_3 = InData_Switch[3 : 3];
  assign _zz_addra_4 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_4 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_4 = InData_Switch[4 : 4];
  assign _zz_addra_5 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_5 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_5 = InData_Switch[5 : 5];
  assign _zz_addra_6 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_6 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_6 = InData_Switch[6 : 6];
  assign _zz_addra_7 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_7 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_7 = InData_Switch[7 : 7];
  assign _zz_addra_8 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_8 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_8 = InData_Switch[8 : 8];
  assign _zz_addra_9 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_9 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_9 = InData_Switch[9 : 9];
  assign _zz_addra_10 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_10 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_10 = InData_Switch[10 : 10];
  assign _zz_addra_11 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_11 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_11 = InData_Switch[11 : 11];
  assign _zz_addra_12 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_12 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_12 = InData_Switch[12 : 12];
  assign _zz_addra_13 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_13 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_13 = InData_Switch[13 : 13];
  assign _zz_addra_14 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_14 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_14 = InData_Switch[14 : 14];
  assign _zz_addra_15 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_15 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_15 = InData_Switch[15 : 15];
  assign _zz_addra_16 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_16 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_16 = InData_Switch[16 : 16];
  assign _zz_addra_17 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_17 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_17 = InData_Switch[17 : 17];
  assign _zz_addra_18 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_18 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_18 = InData_Switch[18 : 18];
  assign _zz_addra_19 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_19 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_19 = InData_Switch[19 : 19];
  assign _zz_addra_20 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_20 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_20 = InData_Switch[20 : 20];
  assign _zz_addra_21 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_21 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_21 = InData_Switch[21 : 21];
  assign _zz_addra_22 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_22 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_22 = InData_Switch[22 : 22];
  assign _zz_addra_23 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_23 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_23 = InData_Switch[23 : 23];
  assign _zz_addra_24 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_24 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_24 = InData_Switch[24 : 24];
  assign _zz_addra_25 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_25 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_25 = InData_Switch[25 : 25];
  assign _zz_addra_26 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_26 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_26 = InData_Switch[26 : 26];
  assign _zz_addra_27 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_27 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_27 = InData_Switch[27 : 27];
  assign _zz_addra_28 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_28 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_28 = InData_Switch[28 : 28];
  assign _zz_addra_29 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_29 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_29 = InData_Switch[29 : 29];
  assign _zz_addra_30 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_30 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_30 = InData_Switch[30 : 30];
  assign _zz_addra_31 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_31 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_31 = InData_Switch[31 : 31];
  assign _zz_addra_32 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_32 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_32 = InData_Switch[32 : 32];
  assign _zz_addra_33 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_33 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_33 = InData_Switch[33 : 33];
  assign _zz_addra_34 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_34 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_34 = InData_Switch[34 : 34];
  assign _zz_addra_35 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_35 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_35 = InData_Switch[35 : 35];
  assign _zz_addra_36 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_36 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_36 = InData_Switch[36 : 36];
  assign _zz_addra_37 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_37 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_37 = InData_Switch[37 : 37];
  assign _zz_addra_38 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_38 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_38 = InData_Switch[38 : 38];
  assign _zz_addra_39 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_39 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_39 = InData_Switch[39 : 39];
  assign _zz_addra_40 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_40 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_40 = InData_Switch[40 : 40];
  assign _zz_addra_41 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_41 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_41 = InData_Switch[41 : 41];
  assign _zz_addra_42 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_42 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_42 = InData_Switch[42 : 42];
  assign _zz_addra_43 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_43 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_43 = InData_Switch[43 : 43];
  assign _zz_addra_44 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_44 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_44 = InData_Switch[44 : 44];
  assign _zz_addra_45 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_45 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_45 = InData_Switch[45 : 45];
  assign _zz_addra_46 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_46 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_46 = InData_Switch[46 : 46];
  assign _zz_addra_47 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_47 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_47 = InData_Switch[47 : 47];
  assign _zz_addra_48 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_48 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_48 = InData_Switch[48 : 48];
  assign _zz_addra_49 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_49 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_49 = InData_Switch[49 : 49];
  assign _zz_addra_50 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_50 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_50 = InData_Switch[50 : 50];
  assign _zz_addra_51 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_51 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_51 = InData_Switch[51 : 51];
  assign _zz_addra_52 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_52 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_52 = InData_Switch[52 : 52];
  assign _zz_addra_53 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_53 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_53 = InData_Switch[53 : 53];
  assign _zz_addra_54 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_54 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_54 = InData_Switch[54 : 54];
  assign _zz_addra_55 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_55 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_55 = InData_Switch[55 : 55];
  assign _zz_addra_56 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_56 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_56 = InData_Switch[56 : 56];
  assign _zz_addra_57 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_57 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_57 = InData_Switch[57 : 57];
  assign _zz_addra_58 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_58 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_58 = InData_Switch[58 : 58];
  assign _zz_addra_59 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_59 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_59 = InData_Switch[59 : 59];
  assign _zz_addra_60 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_60 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_60 = InData_Switch[60 : 60];
  assign _zz_addra_61 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_61 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_61 = InData_Switch[61 : 61];
  assign _zz_addra_62 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_62 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_62 = InData_Switch[62 : 62];
  assign _zz_addra_63 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_63 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_63 = InData_Switch[63 : 63];
  assign _zz_addra_64 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_64 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_64 = InData_Switch[64 : 64];
  assign _zz_addra_65 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_65 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_65 = InData_Switch[65 : 65];
  assign _zz_addra_66 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_66 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_66 = InData_Switch[66 : 66];
  assign _zz_addra_67 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_67 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_67 = InData_Switch[67 : 67];
  assign _zz_addra_68 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_68 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_68 = InData_Switch[68 : 68];
  assign _zz_addra_69 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_69 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_69 = InData_Switch[69 : 69];
  assign _zz_addra_70 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_70 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_70 = InData_Switch[70 : 70];
  assign _zz_addra_71 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_71 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_71 = InData_Switch[71 : 71];
  assign _zz_addra_72 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_72 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_72 = InData_Switch[72 : 72];
  assign _zz_addra_73 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_73 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_73 = InData_Switch[73 : 73];
  assign _zz_addra_74 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_74 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_74 = InData_Switch[74 : 74];
  assign _zz_addra_75 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_75 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_75 = InData_Switch[75 : 75];
  assign _zz_addra_76 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_76 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_76 = InData_Switch[76 : 76];
  assign _zz_addra_77 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_77 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_77 = InData_Switch[77 : 77];
  assign _zz_addra_78 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_78 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_78 = InData_Switch[78 : 78];
  assign _zz_addra_79 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_79 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_79 = InData_Switch[79 : 79];
  assign _zz_addra_80 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_80 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_80 = InData_Switch[80 : 80];
  assign _zz_addra_81 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_81 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_81 = InData_Switch[81 : 81];
  assign _zz_addra_82 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_82 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_82 = InData_Switch[82 : 82];
  assign _zz_addra_83 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_83 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_83 = InData_Switch[83 : 83];
  assign _zz_addra_84 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_84 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_84 = InData_Switch[84 : 84];
  assign _zz_addra_85 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_85 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_85 = InData_Switch[85 : 85];
  assign _zz_addra_86 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_86 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_86 = InData_Switch[86 : 86];
  assign _zz_addra_87 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_87 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_87 = InData_Switch[87 : 87];
  assign _zz_addra_88 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_88 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_88 = InData_Switch[88 : 88];
  assign _zz_addra_89 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_89 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_89 = InData_Switch[89 : 89];
  assign _zz_addra_90 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_90 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_90 = InData_Switch[90 : 90];
  assign _zz_addra_91 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_91 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_91 = InData_Switch[91 : 91];
  assign _zz_addra_92 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_92 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_92 = InData_Switch[92 : 92];
  assign _zz_addra_93 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_93 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_93 = InData_Switch[93 : 93];
  assign _zz_addra_94 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_94 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_94 = InData_Switch[94 : 94];
  assign _zz_addra_95 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_95 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_95 = InData_Switch[95 : 95];
  assign _zz_addra_96 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_96 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_96 = InData_Switch[96 : 96];
  assign _zz_addra_97 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_97 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_97 = InData_Switch[97 : 97];
  assign _zz_addra_98 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_98 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_98 = InData_Switch[98 : 98];
  assign _zz_addra_99 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_99 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_99 = InData_Switch[99 : 99];
  assign _zz_addra_100 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_100 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_100 = InData_Switch[100 : 100];
  assign _zz_addra_101 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_101 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_101 = InData_Switch[101 : 101];
  assign _zz_addra_102 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_102 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_102 = InData_Switch[102 : 102];
  assign _zz_addra_103 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_103 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_103 = InData_Switch[103 : 103];
  assign _zz_addra_104 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_104 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_104 = InData_Switch[104 : 104];
  assign _zz_addra_105 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_105 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_105 = InData_Switch[105 : 105];
  assign _zz_addra_106 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_106 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_106 = InData_Switch[106 : 106];
  assign _zz_addra_107 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_107 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_107 = InData_Switch[107 : 107];
  assign _zz_addra_108 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_108 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_108 = InData_Switch[108 : 108];
  assign _zz_addra_109 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_109 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_109 = InData_Switch[109 : 109];
  assign _zz_addra_110 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_110 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_110 = InData_Switch[110 : 110];
  assign _zz_addra_111 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_111 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_111 = InData_Switch[111 : 111];
  assign _zz_addra_112 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_112 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_112 = InData_Switch[112 : 112];
  assign _zz_addra_113 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_113 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_113 = InData_Switch[113 : 113];
  assign _zz_addra_114 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_114 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_114 = InData_Switch[114 : 114];
  assign _zz_addra_115 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_115 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_115 = InData_Switch[115 : 115];
  assign _zz_addra_116 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_116 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_116 = InData_Switch[116 : 116];
  assign _zz_addra_117 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_117 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_117 = InData_Switch[117 : 117];
  assign _zz_addra_118 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_118 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_118 = InData_Switch[118 : 118];
  assign _zz_addra_119 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_119 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_119 = InData_Switch[119 : 119];
  assign _zz_addra_120 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_120 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_120 = InData_Switch[120 : 120];
  assign _zz_addra_121 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_121 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_121 = InData_Switch[121 : 121];
  assign _zz_addra_122 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_122 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_122 = InData_Switch[122 : 122];
  assign _zz_addra_123 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_123 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_123 = InData_Switch[123 : 123];
  assign _zz_addra_124 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_124 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_124 = InData_Switch[124 : 124];
  assign _zz_addra_125 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_125 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_125 = InData_Switch[125 : 125];
  assign _zz_addra_126 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_126 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_126 = InData_Switch[126 : 126];
  assign _zz_addra_127 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_127 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_127 = InData_Switch[127 : 127];
  assign _zz_addra_128 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_128 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_128 = InData_Switch[128 : 128];
  assign _zz_addra_129 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_129 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_129 = InData_Switch[129 : 129];
  assign _zz_addra_130 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_130 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_130 = InData_Switch[130 : 130];
  assign _zz_addra_131 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_131 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_131 = InData_Switch[131 : 131];
  assign _zz_addra_132 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_132 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_132 = InData_Switch[132 : 132];
  assign _zz_addra_133 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_133 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_133 = InData_Switch[133 : 133];
  assign _zz_addra_134 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_134 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_134 = InData_Switch[134 : 134];
  assign _zz_addra_135 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_135 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_135 = InData_Switch[135 : 135];
  assign _zz_addra_136 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_136 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_136 = InData_Switch[136 : 136];
  assign _zz_addra_137 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_137 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_137 = InData_Switch[137 : 137];
  assign _zz_addra_138 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_138 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_138 = InData_Switch[138 : 138];
  assign _zz_addra_139 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_139 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_139 = InData_Switch[139 : 139];
  assign _zz_addra_140 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_140 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_140 = InData_Switch[140 : 140];
  assign _zz_addra_141 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_141 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_141 = InData_Switch[141 : 141];
  assign _zz_addra_142 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_142 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_142 = InData_Switch[142 : 142];
  assign _zz_addra_143 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_143 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_143 = InData_Switch[143 : 143];
  assign _zz_addra_144 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_144 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_144 = InData_Switch[144 : 144];
  assign _zz_addra_145 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_145 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_145 = InData_Switch[145 : 145];
  assign _zz_addra_146 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_146 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_146 = InData_Switch[146 : 146];
  assign _zz_addra_147 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_147 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_147 = InData_Switch[147 : 147];
  assign _zz_addra_148 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_148 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_148 = InData_Switch[148 : 148];
  assign _zz_addra_149 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_149 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_149 = InData_Switch[149 : 149];
  assign _zz_addra_150 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_150 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_150 = InData_Switch[150 : 150];
  assign _zz_addra_151 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_151 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_151 = InData_Switch[151 : 151];
  assign _zz_addra_152 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_152 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_152 = InData_Switch[152 : 152];
  assign _zz_addra_153 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_153 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_153 = InData_Switch[153 : 153];
  assign _zz_addra_154 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_154 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_154 = InData_Switch[154 : 154];
  assign _zz_addra_155 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_155 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_155 = InData_Switch[155 : 155];
  assign _zz_addra_156 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_156 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_156 = InData_Switch[156 : 156];
  assign _zz_addra_157 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_157 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_157 = InData_Switch[157 : 157];
  assign _zz_addra_158 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_158 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_158 = InData_Switch[158 : 158];
  assign _zz_addra_159 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_159 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_159 = InData_Switch[159 : 159];
  assign _zz_addra_160 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_160 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_160 = InData_Switch[160 : 160];
  assign _zz_addra_161 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_161 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_161 = InData_Switch[161 : 161];
  assign _zz_addra_162 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_162 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_162 = InData_Switch[162 : 162];
  assign _zz_addra_163 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_163 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_163 = InData_Switch[163 : 163];
  assign _zz_addra_164 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_164 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_164 = InData_Switch[164 : 164];
  assign _zz_addra_165 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_165 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_165 = InData_Switch[165 : 165];
  assign _zz_addra_166 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_166 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_166 = InData_Switch[166 : 166];
  assign _zz_addra_167 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_167 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_167 = InData_Switch[167 : 167];
  assign _zz_addra_168 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_168 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_168 = InData_Switch[168 : 168];
  assign _zz_addra_169 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_169 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_169 = InData_Switch[169 : 169];
  assign _zz_addra_170 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_170 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_170 = InData_Switch[170 : 170];
  assign _zz_addra_171 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_171 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_171 = InData_Switch[171 : 171];
  assign _zz_addra_172 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_172 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_172 = InData_Switch[172 : 172];
  assign _zz_addra_173 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_173 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_173 = InData_Switch[173 : 173];
  assign _zz_addra_174 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_174 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_174 = InData_Switch[174 : 174];
  assign _zz_addra_175 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_175 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_175 = InData_Switch[175 : 175];
  assign _zz_addra_176 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_176 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_176 = InData_Switch[176 : 176];
  assign _zz_addra_177 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_177 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_177 = InData_Switch[177 : 177];
  assign _zz_addra_178 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_178 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_178 = InData_Switch[178 : 178];
  assign _zz_addra_179 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_179 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_179 = InData_Switch[179 : 179];
  assign _zz_addra_180 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_180 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_180 = InData_Switch[180 : 180];
  assign _zz_addra_181 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_181 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_181 = InData_Switch[181 : 181];
  assign _zz_addra_182 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_182 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_182 = InData_Switch[182 : 182];
  assign _zz_addra_183 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_183 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_183 = InData_Switch[183 : 183];
  assign _zz_addra_184 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_184 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_184 = InData_Switch[184 : 184];
  assign _zz_addra_185 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_185 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_185 = InData_Switch[185 : 185];
  assign _zz_addra_186 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_186 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_186 = InData_Switch[186 : 186];
  assign _zz_addra_187 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_187 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_187 = InData_Switch[187 : 187];
  assign _zz_addra_188 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_188 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_188 = InData_Switch[188 : 188];
  assign _zz_addra_189 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_189 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_189 = InData_Switch[189 : 189];
  assign _zz_addra_190 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_190 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_190 = InData_Switch[190 : 190];
  assign _zz_addra_191 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_191 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_191 = InData_Switch[191 : 191];
  assign _zz_addra_192 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_192 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_192 = InData_Switch[192 : 192];
  assign _zz_addra_193 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_193 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_193 = InData_Switch[193 : 193];
  assign _zz_addra_194 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_194 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_194 = InData_Switch[194 : 194];
  assign _zz_addra_195 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_195 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_195 = InData_Switch[195 : 195];
  assign _zz_addra_196 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_196 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_196 = InData_Switch[196 : 196];
  assign _zz_addra_197 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_197 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_197 = InData_Switch[197 : 197];
  assign _zz_addra_198 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_198 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_198 = InData_Switch[198 : 198];
  assign _zz_addra_199 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_199 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_199 = InData_Switch[199 : 199];
  assign _zz_addra_200 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_200 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_200 = InData_Switch[200 : 200];
  assign _zz_addra_201 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_201 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_201 = InData_Switch[201 : 201];
  assign _zz_addra_202 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_202 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_202 = InData_Switch[202 : 202];
  assign _zz_addra_203 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_203 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_203 = InData_Switch[203 : 203];
  assign _zz_addra_204 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_204 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_204 = InData_Switch[204 : 204];
  assign _zz_addra_205 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_205 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_205 = InData_Switch[205 : 205];
  assign _zz_addra_206 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_206 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_206 = InData_Switch[206 : 206];
  assign _zz_addra_207 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_207 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_207 = InData_Switch[207 : 207];
  assign _zz_addra_208 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_208 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_208 = InData_Switch[208 : 208];
  assign _zz_addra_209 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_209 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_209 = InData_Switch[209 : 209];
  assign _zz_addra_210 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_210 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_210 = InData_Switch[210 : 210];
  assign _zz_addra_211 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_211 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_211 = InData_Switch[211 : 211];
  assign _zz_addra_212 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_212 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_212 = InData_Switch[212 : 212];
  assign _zz_addra_213 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_213 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_213 = InData_Switch[213 : 213];
  assign _zz_addra_214 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_214 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_214 = InData_Switch[214 : 214];
  assign _zz_addra_215 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_215 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_215 = InData_Switch[215 : 215];
  assign _zz_addra_216 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_216 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_216 = InData_Switch[216 : 216];
  assign _zz_addra_217 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_217 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_217 = InData_Switch[217 : 217];
  assign _zz_addra_218 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_218 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_218 = InData_Switch[218 : 218];
  assign _zz_addra_219 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_219 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_219 = InData_Switch[219 : 219];
  assign _zz_addra_220 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_220 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_220 = InData_Switch[220 : 220];
  assign _zz_addra_221 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_221 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_221 = InData_Switch[221 : 221];
  assign _zz_addra_222 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_222 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_222 = InData_Switch[222 : 222];
  assign _zz_addra_223 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_223 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_223 = InData_Switch[223 : 223];
  assign _zz_addra_224 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_224 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_224 = InData_Switch[224 : 224];
  assign _zz_addra_225 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_225 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_225 = InData_Switch[225 : 225];
  assign _zz_addra_226 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_226 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_226 = InData_Switch[226 : 226];
  assign _zz_addra_227 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_227 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_227 = InData_Switch[227 : 227];
  assign _zz_addra_228 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_228 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_228 = InData_Switch[228 : 228];
  assign _zz_addra_229 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_229 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_229 = InData_Switch[229 : 229];
  assign _zz_addra_230 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_230 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_230 = InData_Switch[230 : 230];
  assign _zz_addra_231 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_231 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_231 = InData_Switch[231 : 231];
  assign _zz_addra_232 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_232 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_232 = InData_Switch[232 : 232];
  assign _zz_addra_233 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_233 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_233 = InData_Switch[233 : 233];
  assign _zz_addra_234 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_234 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_234 = InData_Switch[234 : 234];
  assign _zz_addra_235 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_235 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_235 = InData_Switch[235 : 235];
  assign _zz_addra_236 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_236 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_236 = InData_Switch[236 : 236];
  assign _zz_addra_237 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_237 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_237 = InData_Switch[237 : 237];
  assign _zz_addra_238 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_238 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_238 = InData_Switch[238 : 238];
  assign _zz_addra_239 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_239 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_239 = InData_Switch[239 : 239];
  assign _zz_addra_240 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_240 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_240 = InData_Switch[240 : 240];
  assign _zz_addra_241 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_241 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_241 = InData_Switch[241 : 241];
  assign _zz_addra_242 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_242 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_242 = InData_Switch[242 : 242];
  assign _zz_addra_243 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_243 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_243 = InData_Switch[243 : 243];
  assign _zz_addra_244 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_244 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_244 = InData_Switch[244 : 244];
  assign _zz_addra_245 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_245 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_245 = InData_Switch[245 : 245];
  assign _zz_addra_246 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_246 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_246 = InData_Switch[246 : 246];
  assign _zz_addra_247 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_247 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_247 = InData_Switch[247 : 247];
  assign _zz_addra_248 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_248 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_248 = InData_Switch[248 : 248];
  assign _zz_addra_249 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_249 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_249 = InData_Switch[249 : 249];
  assign _zz_addra_250 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_250 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_250 = InData_Switch[250 : 250];
  assign _zz_addra_251 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_251 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_251 = InData_Switch[251 : 251];
  assign _zz_addra_252 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_252 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_252 = InData_Switch[252 : 252];
  assign _zz_addra_253 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_253 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_253 = InData_Switch[253 : 253];
  assign _zz_addra_254 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_254 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_254 = InData_Switch[254 : 254];
  assign _zz_addra_255 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_255 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_255 = InData_Switch[255 : 255];
  assign _zz_addra_256 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_256 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_256 = InData_Switch[256 : 256];
  assign _zz_addra_257 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_257 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_257 = InData_Switch[257 : 257];
  assign _zz_addra_258 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_258 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_258 = InData_Switch[258 : 258];
  assign _zz_addra_259 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_259 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_259 = InData_Switch[259 : 259];
  assign _zz_addra_260 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_260 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_260 = InData_Switch[260 : 260];
  assign _zz_addra_261 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_261 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_261 = InData_Switch[261 : 261];
  assign _zz_addra_262 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_262 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_262 = InData_Switch[262 : 262];
  assign _zz_addra_263 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_263 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_263 = InData_Switch[263 : 263];
  assign _zz_addra_264 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_264 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_264 = InData_Switch[264 : 264];
  assign _zz_addra_265 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_265 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_265 = InData_Switch[265 : 265];
  assign _zz_addra_266 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_266 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_266 = InData_Switch[266 : 266];
  assign _zz_addra_267 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_267 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_267 = InData_Switch[267 : 267];
  assign _zz_addra_268 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_268 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_268 = InData_Switch[268 : 268];
  assign _zz_addra_269 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_269 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_269 = InData_Switch[269 : 269];
  assign _zz_addra_270 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_270 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_270 = InData_Switch[270 : 270];
  assign _zz_addra_271 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_271 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_271 = InData_Switch[271 : 271];
  assign _zz_addra_272 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_272 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_272 = InData_Switch[272 : 272];
  assign _zz_addra_273 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_273 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_273 = InData_Switch[273 : 273];
  assign _zz_addra_274 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_274 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_274 = InData_Switch[274 : 274];
  assign _zz_addra_275 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_275 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_275 = InData_Switch[275 : 275];
  assign _zz_addra_276 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_276 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_276 = InData_Switch[276 : 276];
  assign _zz_addra_277 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_277 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_277 = InData_Switch[277 : 277];
  assign _zz_addra_278 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_278 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_278 = InData_Switch[278 : 278];
  assign _zz_addra_279 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_279 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_279 = InData_Switch[279 : 279];
  assign _zz_addra_280 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_280 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_280 = InData_Switch[280 : 280];
  assign _zz_addra_281 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_281 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_281 = InData_Switch[281 : 281];
  assign _zz_addra_282 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_282 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_282 = InData_Switch[282 : 282];
  assign _zz_addra_283 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_283 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_283 = InData_Switch[283 : 283];
  assign _zz_addra_284 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_284 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_284 = InData_Switch[284 : 284];
  assign _zz_addra_285 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_285 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_285 = InData_Switch[285 : 285];
  assign _zz_addra_286 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_286 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_286 = InData_Switch[286 : 286];
  assign _zz_addra_287 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_287 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_287 = InData_Switch[287 : 287];
  assign _zz_addra_288 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_288 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_288 = InData_Switch[288 : 288];
  assign _zz_addra_289 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_289 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_289 = InData_Switch[289 : 289];
  assign _zz_addra_290 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_290 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_290 = InData_Switch[290 : 290];
  assign _zz_addra_291 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_291 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_291 = InData_Switch[291 : 291];
  assign _zz_addra_292 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_292 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_292 = InData_Switch[292 : 292];
  assign _zz_addra_293 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_293 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_293 = InData_Switch[293 : 293];
  assign _zz_addra_294 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_294 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_294 = InData_Switch[294 : 294];
  assign _zz_addra_295 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_295 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_295 = InData_Switch[295 : 295];
  assign _zz_addra_296 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_296 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_296 = InData_Switch[296 : 296];
  assign _zz_addra_297 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_297 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_297 = InData_Switch[297 : 297];
  assign _zz_addra_298 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_298 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_298 = InData_Switch[298 : 298];
  assign _zz_addra_299 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_299 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_299 = InData_Switch[299 : 299];
  assign _zz_addra_300 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_300 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_300 = InData_Switch[300 : 300];
  assign _zz_addra_301 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_301 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_301 = InData_Switch[301 : 301];
  assign _zz_addra_302 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_302 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_302 = InData_Switch[302 : 302];
  assign _zz_addra_303 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_303 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_303 = InData_Switch[303 : 303];
  assign _zz_addra_304 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_304 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_304 = InData_Switch[304 : 304];
  assign _zz_addra_305 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_305 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_305 = InData_Switch[305 : 305];
  assign _zz_addra_306 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_306 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_306 = InData_Switch[306 : 306];
  assign _zz_addra_307 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_307 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_307 = InData_Switch[307 : 307];
  assign _zz_addra_308 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_308 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_308 = InData_Switch[308 : 308];
  assign _zz_addra_309 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_309 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_309 = InData_Switch[309 : 309];
  assign _zz_addra_310 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_310 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_310 = InData_Switch[310 : 310];
  assign _zz_addra_311 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_311 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_311 = InData_Switch[311 : 311];
  assign _zz_addra_312 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_312 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_312 = InData_Switch[312 : 312];
  assign _zz_addra_313 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_313 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_313 = InData_Switch[313 : 313];
  assign _zz_addra_314 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_314 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_314 = InData_Switch[314 : 314];
  assign _zz_addra_315 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_315 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_315 = InData_Switch[315 : 315];
  assign _zz_addra_316 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_316 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_316 = InData_Switch[316 : 316];
  assign _zz_addra_317 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_317 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_317 = InData_Switch[317 : 317];
  assign _zz_addra_318 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_318 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_318 = InData_Switch[318 : 318];
  assign _zz_addra_319 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_319 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_319 = InData_Switch[319 : 319];
  assign _zz_addra_320 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_320 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_320 = InData_Switch[320 : 320];
  assign _zz_addra_321 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_321 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_321 = InData_Switch[321 : 321];
  assign _zz_addra_322 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_322 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_322 = InData_Switch[322 : 322];
  assign _zz_addra_323 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_323 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_323 = InData_Switch[323 : 323];
  assign _zz_addra_324 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_324 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_324 = InData_Switch[324 : 324];
  assign _zz_addra_325 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_325 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_325 = InData_Switch[325 : 325];
  assign _zz_addra_326 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_326 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_326 = InData_Switch[326 : 326];
  assign _zz_addra_327 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_327 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_327 = InData_Switch[327 : 327];
  assign _zz_addra_328 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_328 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_328 = InData_Switch[328 : 328];
  assign _zz_addra_329 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_329 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_329 = InData_Switch[329 : 329];
  assign _zz_addra_330 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_330 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_330 = InData_Switch[330 : 330];
  assign _zz_addra_331 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_331 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_331 = InData_Switch[331 : 331];
  assign _zz_addra_332 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_332 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_332 = InData_Switch[332 : 332];
  assign _zz_addra_333 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_333 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_333 = InData_Switch[333 : 333];
  assign _zz_addra_334 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_334 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_334 = InData_Switch[334 : 334];
  assign _zz_addra_335 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_335 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_335 = InData_Switch[335 : 335];
  assign _zz_addra_336 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_336 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_336 = InData_Switch[336 : 336];
  assign _zz_addra_337 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_337 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_337 = InData_Switch[337 : 337];
  assign _zz_addra_338 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_338 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_338 = InData_Switch[338 : 338];
  assign _zz_addra_339 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_339 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_339 = InData_Switch[339 : 339];
  assign _zz_addra_340 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_340 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_340 = InData_Switch[340 : 340];
  assign _zz_addra_341 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_341 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_341 = InData_Switch[341 : 341];
  assign _zz_addra_342 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_342 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_342 = InData_Switch[342 : 342];
  assign _zz_addra_343 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_343 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_343 = InData_Switch[343 : 343];
  assign _zz_addra_344 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_344 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_344 = InData_Switch[344 : 344];
  assign _zz_addra_345 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_345 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_345 = InData_Switch[345 : 345];
  assign _zz_addra_346 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_346 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_346 = InData_Switch[346 : 346];
  assign _zz_addra_347 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_347 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_347 = InData_Switch[347 : 347];
  assign _zz_addra_348 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_348 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_348 = InData_Switch[348 : 348];
  assign _zz_addra_349 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_349 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_349 = InData_Switch[349 : 349];
  assign _zz_addra_350 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_350 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_350 = InData_Switch[350 : 350];
  assign _zz_addra_351 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_351 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_351 = InData_Switch[351 : 351];
  assign _zz_addra_352 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_352 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_352 = InData_Switch[352 : 352];
  assign _zz_addra_353 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_353 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_353 = InData_Switch[353 : 353];
  assign _zz_addra_354 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_354 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_354 = InData_Switch[354 : 354];
  assign _zz_addra_355 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_355 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_355 = InData_Switch[355 : 355];
  assign _zz_addra_356 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_356 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_356 = InData_Switch[356 : 356];
  assign _zz_addra_357 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_357 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_357 = InData_Switch[357 : 357];
  assign _zz_addra_358 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_358 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_358 = InData_Switch[358 : 358];
  assign _zz_addra_359 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_359 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_359 = InData_Switch[359 : 359];
  assign _zz_addra_360 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_360 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_360 = InData_Switch[360 : 360];
  assign _zz_addra_361 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_361 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_361 = InData_Switch[361 : 361];
  assign _zz_addra_362 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_362 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_362 = InData_Switch[362 : 362];
  assign _zz_addra_363 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_363 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_363 = InData_Switch[363 : 363];
  assign _zz_addra_364 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_364 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_364 = InData_Switch[364 : 364];
  assign _zz_addra_365 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_365 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_365 = InData_Switch[365 : 365];
  assign _zz_addra_366 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_366 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_366 = InData_Switch[366 : 366];
  assign _zz_addra_367 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_367 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_367 = InData_Switch[367 : 367];
  assign _zz_addra_368 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_368 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_368 = InData_Switch[368 : 368];
  assign _zz_addra_369 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_369 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_369 = InData_Switch[369 : 369];
  assign _zz_addra_370 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_370 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_370 = InData_Switch[370 : 370];
  assign _zz_addra_371 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_371 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_371 = InData_Switch[371 : 371];
  assign _zz_addra_372 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_372 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_372 = InData_Switch[372 : 372];
  assign _zz_addra_373 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_373 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_373 = InData_Switch[373 : 373];
  assign _zz_addra_374 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_374 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_374 = InData_Switch[374 : 374];
  assign _zz_addra_375 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_375 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_375 = InData_Switch[375 : 375];
  assign _zz_addra_376 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_376 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_376 = InData_Switch[376 : 376];
  assign _zz_addra_377 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_377 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_377 = InData_Switch[377 : 377];
  assign _zz_addra_378 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_378 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_378 = InData_Switch[378 : 378];
  assign _zz_addra_379 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_379 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_379 = InData_Switch[379 : 379];
  assign _zz_addra_380 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_380 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_380 = InData_Switch[380 : 380];
  assign _zz_addra_381 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_381 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_381 = InData_Switch[381 : 381];
  assign _zz_addra_382 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_382 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_382 = InData_Switch[382 : 382];
  assign _zz_addra_383 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_383 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_383 = InData_Switch[383 : 383];
  assign _zz_addra_384 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_384 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_384 = InData_Switch[384 : 384];
  assign _zz_addra_385 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_385 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_385 = InData_Switch[385 : 385];
  assign _zz_addra_386 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_386 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_386 = InData_Switch[386 : 386];
  assign _zz_addra_387 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_387 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_387 = InData_Switch[387 : 387];
  assign _zz_addra_388 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_388 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_388 = InData_Switch[388 : 388];
  assign _zz_addra_389 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_389 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_389 = InData_Switch[389 : 389];
  assign _zz_addra_390 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_390 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_390 = InData_Switch[390 : 390];
  assign _zz_addra_391 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_391 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_391 = InData_Switch[391 : 391];
  assign _zz_addra_392 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_392 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_392 = InData_Switch[392 : 392];
  assign _zz_addra_393 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_393 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_393 = InData_Switch[393 : 393];
  assign _zz_addra_394 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_394 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_394 = InData_Switch[394 : 394];
  assign _zz_addra_395 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_395 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_395 = InData_Switch[395 : 395];
  assign _zz_addra_396 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_396 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_396 = InData_Switch[396 : 396];
  assign _zz_addra_397 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_397 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_397 = InData_Switch[397 : 397];
  assign _zz_addra_398 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_398 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_398 = InData_Switch[398 : 398];
  assign _zz_addra_399 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_399 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_399 = InData_Switch[399 : 399];
  assign _zz_addra_400 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_400 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_400 = InData_Switch[400 : 400];
  assign _zz_addra_401 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_401 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_401 = InData_Switch[401 : 401];
  assign _zz_addra_402 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_402 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_402 = InData_Switch[402 : 402];
  assign _zz_addra_403 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_403 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_403 = InData_Switch[403 : 403];
  assign _zz_addra_404 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_404 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_404 = InData_Switch[404 : 404];
  assign _zz_addra_405 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_405 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_405 = InData_Switch[405 : 405];
  assign _zz_addra_406 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_406 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_406 = InData_Switch[406 : 406];
  assign _zz_addra_407 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_407 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_407 = InData_Switch[407 : 407];
  assign _zz_addra_408 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_408 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_408 = InData_Switch[408 : 408];
  assign _zz_addra_409 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_409 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_409 = InData_Switch[409 : 409];
  assign _zz_addra_410 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_410 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_410 = InData_Switch[410 : 410];
  assign _zz_addra_411 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_411 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_411 = InData_Switch[411 : 411];
  assign _zz_addra_412 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_412 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_412 = InData_Switch[412 : 412];
  assign _zz_addra_413 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_413 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_413 = InData_Switch[413 : 413];
  assign _zz_addra_414 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_414 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_414 = InData_Switch[414 : 414];
  assign _zz_addra_415 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_415 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_415 = InData_Switch[415 : 415];
  assign _zz_addra_416 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_416 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_416 = InData_Switch[416 : 416];
  assign _zz_addra_417 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_417 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_417 = InData_Switch[417 : 417];
  assign _zz_addra_418 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_418 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_418 = InData_Switch[418 : 418];
  assign _zz_addra_419 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_419 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_419 = InData_Switch[419 : 419];
  assign _zz_addra_420 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_420 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_420 = InData_Switch[420 : 420];
  assign _zz_addra_421 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_421 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_421 = InData_Switch[421 : 421];
  assign _zz_addra_422 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_422 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_422 = InData_Switch[422 : 422];
  assign _zz_addra_423 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_423 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_423 = InData_Switch[423 : 423];
  assign _zz_addra_424 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_424 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_424 = InData_Switch[424 : 424];
  assign _zz_addra_425 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_425 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_425 = InData_Switch[425 : 425];
  assign _zz_addra_426 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_426 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_426 = InData_Switch[426 : 426];
  assign _zz_addra_427 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_427 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_427 = InData_Switch[427 : 427];
  assign _zz_addra_428 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_428 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_428 = InData_Switch[428 : 428];
  assign _zz_addra_429 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_429 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_429 = InData_Switch[429 : 429];
  assign _zz_addra_430 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_430 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_430 = InData_Switch[430 : 430];
  assign _zz_addra_431 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_431 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_431 = InData_Switch[431 : 431];
  assign _zz_addra_432 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_432 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_432 = InData_Switch[432 : 432];
  assign _zz_addra_433 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_433 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_433 = InData_Switch[433 : 433];
  assign _zz_addra_434 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_434 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_434 = InData_Switch[434 : 434];
  assign _zz_addra_435 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_435 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_435 = InData_Switch[435 : 435];
  assign _zz_addra_436 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_436 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_436 = InData_Switch[436 : 436];
  assign _zz_addra_437 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_437 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_437 = InData_Switch[437 : 437];
  assign _zz_addra_438 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_438 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_438 = InData_Switch[438 : 438];
  assign _zz_addra_439 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_439 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_439 = InData_Switch[439 : 439];
  assign _zz_addra_440 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_440 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_440 = InData_Switch[440 : 440];
  assign _zz_addra_441 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_441 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_441 = InData_Switch[441 : 441];
  assign _zz_addra_442 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_442 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_442 = InData_Switch[442 : 442];
  assign _zz_addra_443 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_443 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_443 = InData_Switch[443 : 443];
  assign _zz_addra_444 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_444 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_444 = InData_Switch[444 : 444];
  assign _zz_addra_445 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_445 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_445 = InData_Switch[445 : 445];
  assign _zz_addra_446 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_446 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_446 = InData_Switch[446 : 446];
  assign _zz_addra_447 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_447 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_447 = InData_Switch[447 : 447];
  assign _zz_addra_448 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_448 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_448 = InData_Switch[448 : 448];
  assign _zz_addra_449 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_449 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_449 = InData_Switch[449 : 449];
  assign _zz_addra_450 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_450 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_450 = InData_Switch[450 : 450];
  assign _zz_addra_451 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_451 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_451 = InData_Switch[451 : 451];
  assign _zz_addra_452 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_452 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_452 = InData_Switch[452 : 452];
  assign _zz_addra_453 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_453 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_453 = InData_Switch[453 : 453];
  assign _zz_addra_454 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_454 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_454 = InData_Switch[454 : 454];
  assign _zz_addra_455 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_455 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_455 = InData_Switch[455 : 455];
  assign _zz_addra_456 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_456 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_456 = InData_Switch[456 : 456];
  assign _zz_addra_457 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_457 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_457 = InData_Switch[457 : 457];
  assign _zz_addra_458 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_458 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_458 = InData_Switch[458 : 458];
  assign _zz_addra_459 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_459 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_459 = InData_Switch[459 : 459];
  assign _zz_addra_460 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_460 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_460 = InData_Switch[460 : 460];
  assign _zz_addra_461 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_461 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_461 = InData_Switch[461 : 461];
  assign _zz_addra_462 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_462 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_462 = InData_Switch[462 : 462];
  assign _zz_addra_463 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_463 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_463 = InData_Switch[463 : 463];
  assign _zz_addra_464 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_464 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_464 = InData_Switch[464 : 464];
  assign _zz_addra_465 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_465 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_465 = InData_Switch[465 : 465];
  assign _zz_addra_466 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_466 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_466 = InData_Switch[466 : 466];
  assign _zz_addra_467 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_467 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_467 = InData_Switch[467 : 467];
  assign _zz_addra_468 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_468 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_468 = InData_Switch[468 : 468];
  assign _zz_addra_469 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_469 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_469 = InData_Switch[469 : 469];
  assign _zz_addra_470 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_470 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_470 = InData_Switch[470 : 470];
  assign _zz_addra_471 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_471 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_471 = InData_Switch[471 : 471];
  assign _zz_addra_472 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_472 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_472 = InData_Switch[472 : 472];
  assign _zz_addra_473 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_473 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_473 = InData_Switch[473 : 473];
  assign _zz_addra_474 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_474 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_474 = InData_Switch[474 : 474];
  assign _zz_addra_475 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_475 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_475 = InData_Switch[475 : 475];
  assign _zz_addra_476 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_476 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_476 = InData_Switch[476 : 476];
  assign _zz_addra_477 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_477 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_477 = InData_Switch[477 : 477];
  assign _zz_addra_478 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_478 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_478 = InData_Switch[478 : 478];
  assign _zz_addra_479 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_479 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_479 = InData_Switch[479 : 479];
  assign _zz_addra_480 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_480 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_480 = InData_Switch[480 : 480];
  assign _zz_addra_481 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_481 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_481 = InData_Switch[481 : 481];
  assign _zz_addra_482 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_482 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_482 = InData_Switch[482 : 482];
  assign _zz_addra_483 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_483 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_483 = InData_Switch[483 : 483];
  assign _zz_addra_484 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_484 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_484 = InData_Switch[484 : 484];
  assign _zz_addra_485 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_485 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_485 = InData_Switch[485 : 485];
  assign _zz_addra_486 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_486 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_486 = InData_Switch[486 : 486];
  assign _zz_addra_487 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_487 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_487 = InData_Switch[487 : 487];
  assign _zz_addra_488 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_488 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_488 = InData_Switch[488 : 488];
  assign _zz_addra_489 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_489 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_489 = InData_Switch[489 : 489];
  assign _zz_addra_490 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_490 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_490 = InData_Switch[490 : 490];
  assign _zz_addra_491 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_491 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_491 = InData_Switch[491 : 491];
  assign _zz_addra_492 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_492 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_492 = InData_Switch[492 : 492];
  assign _zz_addra_493 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_493 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_493 = InData_Switch[493 : 493];
  assign _zz_addra_494 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_494 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_494 = InData_Switch[494 : 494];
  assign _zz_addra_495 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_495 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_495 = InData_Switch[495 : 495];
  assign _zz_addra_496 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_496 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_496 = InData_Switch[496 : 496];
  assign _zz_addra_497 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_497 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_497 = InData_Switch[497 : 497];
  assign _zz_addra_498 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_498 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_498 = InData_Switch[498 : 498];
  assign _zz_addra_499 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_499 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_499 = InData_Switch[499 : 499];
  assign _zz_addra_500 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_500 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_500 = InData_Switch[500 : 500];
  assign _zz_addra_501 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_501 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_501 = InData_Switch[501 : 501];
  assign _zz_addra_502 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_502 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_502 = InData_Switch[502 : 502];
  assign _zz_addra_503 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_503 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_503 = InData_Switch[503 : 503];
  assign _zz_addra_504 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_504 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_504 = InData_Switch[504 : 504];
  assign _zz_addra_505 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_505 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_505 = InData_Switch[505 : 505];
  assign _zz_addra_506 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_506 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_506 = InData_Switch[506 : 506];
  assign _zz_addra_507 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_507 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_507 = InData_Switch[507 : 507];
  assign _zz_addra_508 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_508 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_508 = InData_Switch[508 : 508];
  assign _zz_addra_509 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_509 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_509 = InData_Switch[509 : 509];
  assign _zz_addra_510 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_510 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_510 = InData_Switch[510 : 510];
  assign _zz_addra_511 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_511 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_511 = InData_Switch[511 : 511];
  Weight_Bram xil_SimpleDualBram (
    .clka  (clk                           ), //i
    .addra (xil_SimpleDualBram_addra[10:0]), //i
    .dina  (sData_payload[63:0]           ), //i
    .ena   (xil_SimpleDualBram_ena        ), //i
    .wea   (1'b1                          ), //i
    .addrb (xil_SimpleDualBram_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_doutb[7:0] ), //o
    .clkb  (clk                           )  //i
  );
  Weight_Bram xil_SimpleDualBram_1 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_1_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_1_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_1_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_1_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_2 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_2_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_2_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_2_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_2_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_3 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_3_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_3_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_3_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_3_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_4 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_4_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_4_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_4_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_4_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_5 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_5_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_5_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_5_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_5_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_6 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_6_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_6_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_6_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_6_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_7 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_7_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_7_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_7_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_7_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_8 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_8_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_8_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_8_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_8_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_9 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_9_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_9_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_9_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_9_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_10 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_10_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_10_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_10_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_10_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_11 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_11_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_11_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_11_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_11_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_12 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_12_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_12_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_12_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_12_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_13 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_13_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_13_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_13_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_13_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_14 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_14_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_14_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_14_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_14_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_15 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_15_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_15_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_15_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_15_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_16 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_16_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_16_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_16_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_16_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_17 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_17_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_17_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_17_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_17_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_18 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_18_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_18_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_18_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_18_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_19 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_19_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_19_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_19_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_19_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_20 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_20_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_20_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_20_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_20_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_21 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_21_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_21_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_21_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_21_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_22 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_22_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_22_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_22_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_22_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_23 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_23_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_23_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_23_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_23_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_24 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_24_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_24_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_24_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_24_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_25 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_25_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_25_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_25_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_25_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_26 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_26_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_26_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_26_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_26_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_27 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_27_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_27_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_27_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_27_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_28 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_28_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_28_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_28_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_28_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_29 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_29_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_29_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_29_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_29_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_30 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_30_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_30_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_30_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_30_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_31 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_31_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_31_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_31_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_31_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_32 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_32_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_32_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_32_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_32_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_33 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_33_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_33_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_33_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_33_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_34 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_34_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_34_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_34_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_34_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_35 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_35_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_35_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_35_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_35_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_36 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_36_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_36_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_36_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_36_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_37 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_37_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_37_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_37_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_37_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_38 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_38_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_38_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_38_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_38_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_39 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_39_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_39_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_39_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_39_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_40 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_40_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_40_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_40_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_40_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_41 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_41_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_41_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_41_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_41_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_42 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_42_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_42_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_42_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_42_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_43 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_43_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_43_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_43_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_43_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_44 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_44_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_44_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_44_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_44_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_45 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_45_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_45_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_45_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_45_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_46 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_46_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_46_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_46_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_46_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_47 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_47_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_47_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_47_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_47_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_48 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_48_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_48_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_48_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_48_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_49 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_49_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_49_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_49_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_49_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_50 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_50_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_50_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_50_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_50_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_51 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_51_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_51_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_51_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_51_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_52 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_52_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_52_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_52_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_52_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_53 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_53_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_53_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_53_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_53_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_54 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_54_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_54_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_54_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_54_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_55 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_55_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_55_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_55_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_55_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_56 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_56_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_56_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_56_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_56_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_57 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_57_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_57_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_57_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_57_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_58 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_58_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_58_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_58_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_58_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_59 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_59_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_59_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_59_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_59_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_60 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_60_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_60_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_60_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_60_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_61 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_61_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_61_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_61_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_61_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_62 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_62_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_62_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_62_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_62_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_63 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_63_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_63_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_63_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_63_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_64 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_64_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_64_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_64_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_64_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_65 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_65_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_65_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_65_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_65_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_66 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_66_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_66_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_66_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_66_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_67 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_67_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_67_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_67_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_67_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_68 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_68_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_68_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_68_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_68_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_69 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_69_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_69_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_69_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_69_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_70 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_70_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_70_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_70_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_70_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_71 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_71_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_71_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_71_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_71_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_72 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_72_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_72_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_72_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_72_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_73 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_73_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_73_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_73_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_73_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_74 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_74_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_74_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_74_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_74_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_75 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_75_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_75_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_75_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_75_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_76 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_76_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_76_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_76_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_76_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_77 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_77_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_77_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_77_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_77_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_78 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_78_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_78_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_78_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_78_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_79 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_79_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_79_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_79_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_79_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_80 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_80_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_80_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_80_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_80_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_81 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_81_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_81_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_81_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_81_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_82 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_82_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_82_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_82_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_82_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_83 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_83_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_83_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_83_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_83_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_84 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_84_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_84_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_84_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_84_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_85 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_85_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_85_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_85_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_85_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_86 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_86_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_86_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_86_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_86_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_87 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_87_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_87_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_87_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_87_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_88 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_88_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_88_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_88_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_88_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_89 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_89_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_89_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_89_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_89_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_90 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_90_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_90_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_90_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_90_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_91 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_91_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_91_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_91_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_91_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_92 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_92_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_92_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_92_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_92_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_93 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_93_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_93_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_93_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_93_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_94 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_94_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_94_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_94_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_94_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_95 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_95_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_95_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_95_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_95_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_96 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_96_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_96_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_96_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_96_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_97 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_97_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_97_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_97_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_97_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_98 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_98_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_98_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_98_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_98_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_99 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_99_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_99_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_99_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_99_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_100 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_100_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_100_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_100_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_100_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_101 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_101_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_101_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_101_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_101_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_102 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_102_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_102_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_102_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_102_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_103 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_103_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_103_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_103_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_103_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_104 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_104_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_104_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_104_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_104_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_105 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_105_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_105_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_105_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_105_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_106 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_106_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_106_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_106_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_106_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_107 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_107_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_107_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_107_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_107_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_108 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_108_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_108_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_108_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_108_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_109 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_109_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_109_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_109_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_109_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_110 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_110_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_110_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_110_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_110_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_111 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_111_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_111_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_111_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_111_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_112 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_112_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_112_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_112_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_112_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_113 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_113_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_113_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_113_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_113_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_114 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_114_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_114_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_114_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_114_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_115 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_115_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_115_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_115_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_115_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_116 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_116_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_116_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_116_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_116_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_117 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_117_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_117_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_117_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_117_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_118 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_118_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_118_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_118_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_118_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_119 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_119_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_119_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_119_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_119_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_120 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_120_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_120_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_120_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_120_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_121 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_121_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_121_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_121_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_121_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_122 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_122_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_122_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_122_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_122_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_123 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_123_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_123_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_123_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_123_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_124 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_124_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_124_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_124_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_124_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_125 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_125_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_125_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_125_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_125_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_126 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_126_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_126_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_126_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_126_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_127 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_127_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_127_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_127_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_127_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_128 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_128_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_128_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_128_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_128_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_129 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_129_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_129_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_129_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_129_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_130 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_130_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_130_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_130_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_130_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_131 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_131_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_131_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_131_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_131_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_132 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_132_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_132_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_132_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_132_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_133 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_133_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_133_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_133_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_133_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_134 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_134_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_134_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_134_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_134_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_135 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_135_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_135_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_135_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_135_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_136 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_136_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_136_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_136_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_136_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_137 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_137_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_137_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_137_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_137_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_138 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_138_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_138_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_138_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_138_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_139 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_139_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_139_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_139_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_139_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_140 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_140_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_140_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_140_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_140_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_141 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_141_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_141_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_141_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_141_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_142 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_142_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_142_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_142_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_142_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_143 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_143_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_143_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_143_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_143_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_144 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_144_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_144_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_144_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_144_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_145 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_145_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_145_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_145_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_145_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_146 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_146_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_146_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_146_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_146_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_147 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_147_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_147_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_147_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_147_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_148 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_148_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_148_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_148_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_148_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_149 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_149_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_149_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_149_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_149_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_150 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_150_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_150_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_150_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_150_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_151 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_151_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_151_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_151_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_151_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_152 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_152_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_152_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_152_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_152_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_153 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_153_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_153_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_153_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_153_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_154 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_154_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_154_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_154_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_154_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_155 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_155_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_155_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_155_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_155_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_156 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_156_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_156_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_156_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_156_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_157 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_157_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_157_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_157_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_157_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_158 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_158_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_158_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_158_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_158_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_159 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_159_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_159_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_159_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_159_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_160 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_160_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_160_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_160_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_160_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_161 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_161_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_161_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_161_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_161_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_162 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_162_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_162_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_162_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_162_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_163 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_163_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_163_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_163_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_163_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_164 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_164_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_164_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_164_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_164_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_165 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_165_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_165_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_165_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_165_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_166 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_166_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_166_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_166_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_166_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_167 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_167_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_167_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_167_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_167_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_168 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_168_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_168_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_168_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_168_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_169 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_169_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_169_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_169_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_169_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_170 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_170_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_170_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_170_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_170_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_171 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_171_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_171_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_171_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_171_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_172 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_172_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_172_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_172_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_172_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_173 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_173_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_173_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_173_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_173_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_174 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_174_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_174_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_174_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_174_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_175 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_175_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_175_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_175_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_175_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_176 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_176_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_176_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_176_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_176_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_177 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_177_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_177_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_177_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_177_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_178 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_178_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_178_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_178_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_178_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_179 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_179_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_179_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_179_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_179_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_180 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_180_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_180_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_180_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_180_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_181 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_181_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_181_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_181_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_181_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_182 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_182_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_182_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_182_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_182_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_183 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_183_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_183_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_183_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_183_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_184 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_184_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_184_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_184_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_184_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_185 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_185_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_185_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_185_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_185_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_186 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_186_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_186_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_186_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_186_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_187 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_187_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_187_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_187_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_187_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_188 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_188_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_188_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_188_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_188_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_189 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_189_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_189_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_189_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_189_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_190 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_190_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_190_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_190_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_190_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_191 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_191_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_191_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_191_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_191_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_192 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_192_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_192_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_192_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_192_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_193 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_193_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_193_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_193_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_193_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_194 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_194_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_194_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_194_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_194_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_195 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_195_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_195_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_195_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_195_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_196 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_196_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_196_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_196_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_196_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_197 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_197_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_197_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_197_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_197_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_198 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_198_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_198_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_198_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_198_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_199 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_199_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_199_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_199_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_199_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_200 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_200_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_200_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_200_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_200_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_201 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_201_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_201_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_201_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_201_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_202 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_202_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_202_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_202_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_202_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_203 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_203_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_203_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_203_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_203_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_204 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_204_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_204_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_204_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_204_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_205 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_205_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_205_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_205_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_205_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_206 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_206_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_206_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_206_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_206_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_207 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_207_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_207_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_207_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_207_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_208 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_208_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_208_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_208_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_208_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_209 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_209_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_209_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_209_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_209_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_210 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_210_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_210_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_210_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_210_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_211 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_211_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_211_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_211_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_211_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_212 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_212_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_212_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_212_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_212_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_213 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_213_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_213_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_213_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_213_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_214 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_214_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_214_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_214_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_214_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_215 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_215_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_215_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_215_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_215_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_216 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_216_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_216_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_216_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_216_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_217 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_217_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_217_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_217_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_217_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_218 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_218_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_218_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_218_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_218_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_219 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_219_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_219_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_219_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_219_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_220 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_220_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_220_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_220_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_220_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_221 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_221_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_221_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_221_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_221_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_222 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_222_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_222_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_222_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_222_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_223 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_223_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_223_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_223_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_223_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_224 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_224_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_224_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_224_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_224_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_225 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_225_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_225_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_225_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_225_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_226 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_226_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_226_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_226_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_226_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_227 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_227_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_227_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_227_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_227_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_228 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_228_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_228_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_228_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_228_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_229 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_229_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_229_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_229_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_229_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_230 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_230_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_230_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_230_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_230_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_231 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_231_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_231_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_231_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_231_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_232 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_232_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_232_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_232_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_232_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_233 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_233_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_233_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_233_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_233_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_234 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_234_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_234_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_234_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_234_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_235 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_235_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_235_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_235_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_235_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_236 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_236_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_236_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_236_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_236_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_237 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_237_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_237_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_237_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_237_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_238 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_238_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_238_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_238_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_238_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_239 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_239_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_239_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_239_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_239_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_240 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_240_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_240_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_240_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_240_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_241 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_241_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_241_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_241_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_241_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_242 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_242_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_242_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_242_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_242_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_243 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_243_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_243_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_243_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_243_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_244 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_244_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_244_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_244_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_244_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_245 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_245_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_245_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_245_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_245_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_246 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_246_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_246_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_246_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_246_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_247 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_247_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_247_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_247_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_247_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_248 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_248_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_248_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_248_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_248_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_249 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_249_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_249_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_249_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_249_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_250 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_250_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_250_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_250_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_250_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_251 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_251_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_251_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_251_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_251_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_252 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_252_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_252_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_252_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_252_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_253 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_253_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_253_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_253_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_253_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_254 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_254_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_254_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_254_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_254_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_255 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_255_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_255_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_255_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_255_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_256 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_256_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_256_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_256_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_256_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_257 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_257_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_257_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_257_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_257_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_258 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_258_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_258_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_258_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_258_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_259 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_259_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_259_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_259_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_259_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_260 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_260_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_260_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_260_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_260_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_261 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_261_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_261_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_261_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_261_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_262 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_262_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_262_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_262_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_262_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_263 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_263_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_263_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_263_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_263_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_264 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_264_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_264_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_264_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_264_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_265 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_265_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_265_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_265_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_265_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_266 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_266_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_266_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_266_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_266_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_267 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_267_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_267_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_267_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_267_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_268 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_268_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_268_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_268_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_268_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_269 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_269_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_269_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_269_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_269_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_270 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_270_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_270_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_270_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_270_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_271 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_271_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_271_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_271_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_271_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_272 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_272_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_272_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_272_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_272_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_273 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_273_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_273_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_273_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_273_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_274 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_274_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_274_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_274_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_274_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_275 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_275_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_275_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_275_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_275_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_276 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_276_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_276_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_276_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_276_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_277 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_277_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_277_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_277_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_277_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_278 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_278_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_278_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_278_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_278_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_279 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_279_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_279_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_279_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_279_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_280 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_280_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_280_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_280_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_280_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_281 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_281_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_281_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_281_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_281_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_282 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_282_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_282_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_282_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_282_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_283 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_283_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_283_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_283_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_283_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_284 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_284_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_284_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_284_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_284_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_285 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_285_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_285_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_285_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_285_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_286 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_286_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_286_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_286_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_286_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_287 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_287_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_287_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_287_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_287_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_288 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_288_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_288_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_288_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_288_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_289 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_289_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_289_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_289_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_289_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_290 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_290_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_290_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_290_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_290_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_291 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_291_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_291_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_291_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_291_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_292 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_292_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_292_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_292_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_292_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_293 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_293_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_293_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_293_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_293_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_294 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_294_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_294_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_294_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_294_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_295 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_295_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_295_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_295_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_295_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_296 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_296_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_296_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_296_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_296_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_297 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_297_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_297_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_297_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_297_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_298 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_298_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_298_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_298_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_298_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_299 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_299_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_299_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_299_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_299_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_300 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_300_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_300_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_300_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_300_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_301 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_301_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_301_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_301_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_301_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_302 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_302_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_302_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_302_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_302_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_303 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_303_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_303_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_303_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_303_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_304 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_304_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_304_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_304_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_304_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_305 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_305_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_305_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_305_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_305_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_306 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_306_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_306_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_306_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_306_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_307 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_307_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_307_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_307_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_307_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_308 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_308_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_308_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_308_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_308_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_309 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_309_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_309_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_309_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_309_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_310 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_310_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_310_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_310_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_310_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_311 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_311_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_311_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_311_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_311_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_312 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_312_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_312_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_312_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_312_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_313 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_313_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_313_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_313_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_313_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_314 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_314_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_314_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_314_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_314_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_315 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_315_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_315_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_315_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_315_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_316 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_316_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_316_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_316_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_316_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_317 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_317_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_317_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_317_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_317_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_318 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_318_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_318_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_318_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_318_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_319 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_319_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_319_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_319_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_319_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_320 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_320_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_320_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_320_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_320_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_321 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_321_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_321_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_321_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_321_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_322 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_322_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_322_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_322_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_322_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_323 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_323_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_323_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_323_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_323_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_324 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_324_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_324_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_324_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_324_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_325 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_325_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_325_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_325_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_325_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_326 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_326_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_326_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_326_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_326_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_327 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_327_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_327_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_327_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_327_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_328 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_328_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_328_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_328_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_328_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_329 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_329_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_329_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_329_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_329_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_330 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_330_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_330_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_330_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_330_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_331 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_331_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_331_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_331_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_331_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_332 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_332_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_332_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_332_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_332_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_333 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_333_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_333_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_333_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_333_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_334 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_334_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_334_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_334_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_334_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_335 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_335_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_335_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_335_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_335_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_336 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_336_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_336_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_336_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_336_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_337 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_337_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_337_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_337_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_337_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_338 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_338_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_338_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_338_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_338_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_339 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_339_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_339_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_339_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_339_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_340 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_340_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_340_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_340_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_340_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_341 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_341_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_341_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_341_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_341_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_342 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_342_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_342_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_342_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_342_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_343 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_343_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_343_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_343_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_343_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_344 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_344_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_344_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_344_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_344_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_345 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_345_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_345_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_345_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_345_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_346 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_346_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_346_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_346_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_346_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_347 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_347_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_347_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_347_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_347_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_348 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_348_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_348_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_348_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_348_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_349 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_349_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_349_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_349_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_349_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_350 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_350_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_350_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_350_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_350_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_351 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_351_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_351_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_351_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_351_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_352 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_352_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_352_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_352_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_352_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_353 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_353_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_353_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_353_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_353_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_354 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_354_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_354_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_354_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_354_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_355 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_355_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_355_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_355_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_355_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_356 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_356_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_356_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_356_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_356_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_357 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_357_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_357_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_357_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_357_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_358 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_358_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_358_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_358_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_358_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_359 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_359_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_359_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_359_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_359_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_360 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_360_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_360_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_360_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_360_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_361 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_361_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_361_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_361_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_361_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_362 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_362_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_362_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_362_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_362_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_363 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_363_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_363_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_363_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_363_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_364 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_364_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_364_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_364_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_364_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_365 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_365_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_365_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_365_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_365_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_366 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_366_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_366_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_366_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_366_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_367 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_367_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_367_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_367_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_367_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_368 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_368_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_368_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_368_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_368_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_369 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_369_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_369_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_369_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_369_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_370 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_370_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_370_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_370_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_370_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_371 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_371_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_371_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_371_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_371_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_372 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_372_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_372_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_372_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_372_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_373 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_373_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_373_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_373_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_373_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_374 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_374_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_374_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_374_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_374_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_375 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_375_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_375_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_375_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_375_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_376 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_376_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_376_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_376_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_376_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_377 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_377_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_377_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_377_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_377_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_378 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_378_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_378_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_378_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_378_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_379 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_379_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_379_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_379_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_379_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_380 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_380_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_380_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_380_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_380_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_381 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_381_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_381_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_381_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_381_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_382 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_382_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_382_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_382_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_382_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_383 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_383_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_383_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_383_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_383_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_384 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_384_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_384_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_384_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_384_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_385 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_385_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_385_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_385_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_385_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_386 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_386_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_386_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_386_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_386_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_387 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_387_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_387_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_387_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_387_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_388 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_388_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_388_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_388_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_388_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_389 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_389_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_389_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_389_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_389_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_390 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_390_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_390_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_390_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_390_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_391 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_391_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_391_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_391_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_391_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_392 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_392_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_392_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_392_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_392_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_393 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_393_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_393_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_393_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_393_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_394 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_394_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_394_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_394_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_394_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_395 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_395_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_395_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_395_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_395_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_396 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_396_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_396_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_396_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_396_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_397 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_397_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_397_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_397_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_397_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_398 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_398_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_398_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_398_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_398_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_399 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_399_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_399_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_399_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_399_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_400 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_400_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_400_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_400_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_400_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_401 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_401_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_401_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_401_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_401_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_402 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_402_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_402_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_402_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_402_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_403 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_403_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_403_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_403_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_403_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_404 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_404_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_404_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_404_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_404_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_405 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_405_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_405_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_405_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_405_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_406 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_406_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_406_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_406_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_406_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_407 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_407_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_407_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_407_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_407_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_408 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_408_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_408_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_408_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_408_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_409 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_409_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_409_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_409_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_409_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_410 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_410_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_410_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_410_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_410_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_411 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_411_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_411_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_411_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_411_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_412 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_412_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_412_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_412_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_412_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_413 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_413_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_413_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_413_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_413_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_414 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_414_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_414_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_414_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_414_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_415 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_415_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_415_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_415_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_415_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_416 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_416_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_416_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_416_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_416_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_417 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_417_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_417_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_417_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_417_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_418 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_418_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_418_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_418_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_418_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_419 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_419_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_419_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_419_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_419_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_420 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_420_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_420_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_420_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_420_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_421 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_421_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_421_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_421_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_421_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_422 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_422_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_422_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_422_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_422_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_423 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_423_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_423_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_423_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_423_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_424 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_424_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_424_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_424_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_424_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_425 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_425_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_425_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_425_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_425_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_426 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_426_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_426_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_426_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_426_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_427 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_427_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_427_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_427_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_427_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_428 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_428_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_428_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_428_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_428_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_429 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_429_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_429_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_429_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_429_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_430 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_430_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_430_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_430_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_430_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_431 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_431_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_431_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_431_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_431_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_432 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_432_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_432_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_432_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_432_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_433 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_433_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_433_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_433_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_433_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_434 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_434_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_434_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_434_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_434_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_435 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_435_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_435_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_435_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_435_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_436 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_436_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_436_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_436_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_436_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_437 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_437_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_437_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_437_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_437_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_438 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_438_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_438_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_438_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_438_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_439 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_439_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_439_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_439_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_439_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_440 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_440_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_440_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_440_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_440_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_441 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_441_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_441_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_441_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_441_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_442 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_442_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_442_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_442_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_442_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_443 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_443_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_443_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_443_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_443_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_444 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_444_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_444_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_444_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_444_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_445 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_445_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_445_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_445_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_445_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_446 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_446_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_446_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_446_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_446_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_447 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_447_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_447_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_447_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_447_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_448 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_448_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_448_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_448_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_448_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_449 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_449_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_449_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_449_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_449_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_450 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_450_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_450_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_450_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_450_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_451 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_451_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_451_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_451_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_451_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_452 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_452_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_452_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_452_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_452_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_453 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_453_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_453_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_453_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_453_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_454 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_454_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_454_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_454_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_454_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_455 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_455_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_455_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_455_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_455_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_456 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_456_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_456_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_456_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_456_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_457 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_457_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_457_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_457_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_457_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_458 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_458_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_458_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_458_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_458_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_459 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_459_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_459_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_459_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_459_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_460 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_460_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_460_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_460_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_460_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_461 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_461_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_461_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_461_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_461_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_462 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_462_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_462_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_462_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_462_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_463 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_463_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_463_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_463_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_463_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_464 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_464_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_464_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_464_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_464_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_465 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_465_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_465_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_465_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_465_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_466 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_466_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_466_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_466_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_466_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_467 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_467_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_467_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_467_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_467_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_468 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_468_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_468_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_468_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_468_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_469 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_469_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_469_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_469_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_469_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_470 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_470_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_470_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_470_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_470_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_471 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_471_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_471_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_471_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_471_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_472 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_472_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_472_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_472_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_472_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_473 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_473_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_473_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_473_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_473_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_474 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_474_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_474_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_474_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_474_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_475 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_475_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_475_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_475_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_475_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_476 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_476_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_476_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_476_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_476_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_477 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_477_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_477_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_477_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_477_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_478 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_478_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_478_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_478_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_478_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_479 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_479_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_479_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_479_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_479_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_480 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_480_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_480_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_480_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_480_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_481 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_481_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_481_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_481_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_481_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_482 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_482_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_482_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_482_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_482_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_483 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_483_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_483_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_483_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_483_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_484 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_484_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_484_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_484_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_484_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_485 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_485_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_485_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_485_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_485_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_486 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_486_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_486_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_486_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_486_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_487 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_487_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_487_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_487_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_487_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_488 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_488_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_488_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_488_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_488_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_489 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_489_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_489_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_489_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_489_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_490 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_490_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_490_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_490_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_490_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_491 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_491_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_491_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_491_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_491_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_492 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_492_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_492_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_492_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_492_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_493 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_493_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_493_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_493_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_493_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_494 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_494_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_494_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_494_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_494_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_495 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_495_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_495_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_495_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_495_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_496 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_496_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_496_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_496_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_496_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_497 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_497_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_497_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_497_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_497_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_498 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_498_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_498_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_498_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_498_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_499 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_499_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_499_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_499_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_499_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_500 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_500_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_500_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_500_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_500_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_501 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_501_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_501_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_501_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_501_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_502 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_502_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_502_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_502_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_502_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_503 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_503_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_503_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_503_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_503_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_504 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_504_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_504_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_504_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_504_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_505 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_505_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_505_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_505_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_505_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_506 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_506_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_506_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_506_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_506_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_507 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_507_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_507_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_507_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_507_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_508 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_508_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_508_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_508_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_508_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_509 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_509_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_509_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_509_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_509_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_510 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_510_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_510_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_510_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_510_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  Weight_Bram xil_SimpleDualBram_511 (
    .clka  (clk                               ), //i
    .addra (xil_SimpleDualBram_511_addra[10:0]), //i
    .dina  (sData_payload[63:0]               ), //i
    .ena   (xil_SimpleDualBram_511_ena        ), //i
    .wea   (1'b1                              ), //i
    .addrb (xil_SimpleDualBram_511_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_511_doutb[7:0] ), //o
    .clkb  (clk                               )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      WEIGHT_CACHE_STATUS_IDLE : Fsm_currentState_string = "IDLE        ";
      WEIGHT_CACHE_STATUS_INIT : Fsm_currentState_string = "INIT        ";
      WEIGHT_CACHE_STATUS_CACHE_WEIGHT : Fsm_currentState_string = "CACHE_WEIGHT";
      WEIGHT_CACHE_STATUS_SA_COMPUTE : Fsm_currentState_string = "SA_COMPUTE  ";
      default : Fsm_currentState_string = "????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      WEIGHT_CACHE_STATUS_IDLE : Fsm_nextState_string = "IDLE        ";
      WEIGHT_CACHE_STATUS_INIT : Fsm_nextState_string = "INIT        ";
      WEIGHT_CACHE_STATUS_CACHE_WEIGHT : Fsm_nextState_string = "CACHE_WEIGHT";
      WEIGHT_CACHE_STATUS_SA_COMPUTE : Fsm_nextState_string = "SA_COMPUTE  ";
      default : Fsm_nextState_string = "????????????";
    endcase
  end
  `endif

  assign when_SA3D_WeightCache_l33 = (start && (! start_regNext));
  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & WEIGHT_CACHE_STATUS_IDLE) == WEIGHT_CACHE_STATUS_IDLE) : begin
        if(when_SA3D_WeightCache_l33) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_INIT;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_IDLE;
        end
      end
      (((Fsm_currentState) & WEIGHT_CACHE_STATUS_INIT) == WEIGHT_CACHE_STATUS_INIT) : begin
        if(Fsm_Init_End) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_CACHE_WEIGHT;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_INIT;
        end
      end
      (((Fsm_currentState) & WEIGHT_CACHE_STATUS_CACHE_WEIGHT) == WEIGHT_CACHE_STATUS_CACHE_WEIGHT) : begin
        if(Fsm_Weight_All_Cached) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_SA_COMPUTE;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_CACHE_WEIGHT;
        end
      end
      default : begin
        if(Fsm_SA_Computed) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_IDLE;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_SA_COMPUTE;
        end
      end
    endcase
  end

  assign when_WaCounter_l19 = ((Fsm_currentState & WEIGHT_CACHE_STATUS_INIT) != 4'b0000);
  assign when_WaCounter_l14 = (Init_Count_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l14) begin
      Init_Count_valid = 1'b1;
    end else begin
      Init_Count_valid = 1'b0;
    end
  end

  assign Fsm_Init_End = Init_Count_valid;
  assign Matrix_In_MaxCnt = (Matrix_Row >>> 3);
  assign sData_fire = (sData_valid && sData_ready);
  assign In_Row_Cnt_valid = ((In_Row_Cnt_count == _zz_In_Row_Cnt_valid) && sData_fire);
  assign In_Col_Cnt_valid = ((In_Col_Cnt_count == _zz_In_Col_Cnt_valid) && In_Row_Cnt_valid);
  assign when_WaCounter_l40 = (Raddr_Valid && ((Fsm_currentState & WEIGHT_CACHE_STATUS_SA_COMPUTE) != 4'b0000));
  assign OutRow_Cnt_valid = ((OutRow_Cnt_count == _zz_OutRow_Cnt_valid) && when_WaCounter_l40);
  assign _zz_OutCol_Cnt_count = 4'b1000;
  always @(*) begin
    OutCol_Cnt_valid = ((OutCol_Cnt_count <= _zz_OutCol_Cnt_valid) && OutRow_Cnt_valid);
    if(start) begin
      OutCol_Cnt_valid = 1'b0;
    end
  end

  always @(*) begin
    Col_In_8_Cnt_valid = ((Col_In_8_Cnt_count == 9'h1ff) && In_Row_Cnt_valid);
    if(OutCol_Cnt_valid) begin
      Col_In_8_Cnt_valid = 1'b0;
    end
  end

  assign when_SA3D_WeightCache_l129 = ((Fsm_currentState & WEIGHT_CACHE_STATUS_INIT) != 4'b0000);
  assign when_SA3D_WeightCache_l134 = ((Fsm_currentState & WEIGHT_CACHE_STATUS_INIT) != 4'b0000);
  assign Fsm_Weight_All_Cached = In_Col_Cnt_valid;
  assign Weight_Cached = In_Col_Cnt_valid;
  assign xil_SimpleDualBram_addra = _zz_addra[10:0];
  assign xil_SimpleDualBram_addrb = _zz_addrb[13:0];
  assign sData_fire_1 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_ena = (_zz_ena[0] && sData_fire_1);
  assign mData_0 = xil_SimpleDualBram_doutb;
  assign xil_SimpleDualBram_1_addra = _zz_addra_1[10:0];
  assign xil_SimpleDualBram_1_addrb = _zz_addrb_1[13:0];
  assign sData_fire_2 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_1_ena = (_zz_ena_1[0] && sData_fire_2);
  assign mData_1 = xil_SimpleDualBram_1_doutb;
  assign xil_SimpleDualBram_2_addra = _zz_addra_2[10:0];
  assign xil_SimpleDualBram_2_addrb = _zz_addrb_2[13:0];
  assign sData_fire_3 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_2_ena = (_zz_ena_2[0] && sData_fire_3);
  assign mData_2 = xil_SimpleDualBram_2_doutb;
  assign xil_SimpleDualBram_3_addra = _zz_addra_3[10:0];
  assign xil_SimpleDualBram_3_addrb = _zz_addrb_3[13:0];
  assign sData_fire_4 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_3_ena = (_zz_ena_3[0] && sData_fire_4);
  assign mData_3 = xil_SimpleDualBram_3_doutb;
  assign xil_SimpleDualBram_4_addra = _zz_addra_4[10:0];
  assign xil_SimpleDualBram_4_addrb = _zz_addrb_4[13:0];
  assign sData_fire_5 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_4_ena = (_zz_ena_4[0] && sData_fire_5);
  assign mData_4 = xil_SimpleDualBram_4_doutb;
  assign xil_SimpleDualBram_5_addra = _zz_addra_5[10:0];
  assign xil_SimpleDualBram_5_addrb = _zz_addrb_5[13:0];
  assign sData_fire_6 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_5_ena = (_zz_ena_5[0] && sData_fire_6);
  assign mData_5 = xil_SimpleDualBram_5_doutb;
  assign xil_SimpleDualBram_6_addra = _zz_addra_6[10:0];
  assign xil_SimpleDualBram_6_addrb = _zz_addrb_6[13:0];
  assign sData_fire_7 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_6_ena = (_zz_ena_6[0] && sData_fire_7);
  assign mData_6 = xil_SimpleDualBram_6_doutb;
  assign xil_SimpleDualBram_7_addra = _zz_addra_7[10:0];
  assign xil_SimpleDualBram_7_addrb = _zz_addrb_7[13:0];
  assign sData_fire_8 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_7_ena = (_zz_ena_7[0] && sData_fire_8);
  assign mData_7 = xil_SimpleDualBram_7_doutb;
  assign xil_SimpleDualBram_8_addra = _zz_addra_8[10:0];
  assign xil_SimpleDualBram_8_addrb = _zz_addrb_8[13:0];
  assign sData_fire_9 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_8_ena = (_zz_ena_8[0] && sData_fire_9);
  assign mData_8 = xil_SimpleDualBram_8_doutb;
  assign xil_SimpleDualBram_9_addra = _zz_addra_9[10:0];
  assign xil_SimpleDualBram_9_addrb = _zz_addrb_9[13:0];
  assign sData_fire_10 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_9_ena = (_zz_ena_9[0] && sData_fire_10);
  assign mData_9 = xil_SimpleDualBram_9_doutb;
  assign xil_SimpleDualBram_10_addra = _zz_addra_10[10:0];
  assign xil_SimpleDualBram_10_addrb = _zz_addrb_10[13:0];
  assign sData_fire_11 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_10_ena = (_zz_ena_10[0] && sData_fire_11);
  assign mData_10 = xil_SimpleDualBram_10_doutb;
  assign xil_SimpleDualBram_11_addra = _zz_addra_11[10:0];
  assign xil_SimpleDualBram_11_addrb = _zz_addrb_11[13:0];
  assign sData_fire_12 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_11_ena = (_zz_ena_11[0] && sData_fire_12);
  assign mData_11 = xil_SimpleDualBram_11_doutb;
  assign xil_SimpleDualBram_12_addra = _zz_addra_12[10:0];
  assign xil_SimpleDualBram_12_addrb = _zz_addrb_12[13:0];
  assign sData_fire_13 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_12_ena = (_zz_ena_12[0] && sData_fire_13);
  assign mData_12 = xil_SimpleDualBram_12_doutb;
  assign xil_SimpleDualBram_13_addra = _zz_addra_13[10:0];
  assign xil_SimpleDualBram_13_addrb = _zz_addrb_13[13:0];
  assign sData_fire_14 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_13_ena = (_zz_ena_13[0] && sData_fire_14);
  assign mData_13 = xil_SimpleDualBram_13_doutb;
  assign xil_SimpleDualBram_14_addra = _zz_addra_14[10:0];
  assign xil_SimpleDualBram_14_addrb = _zz_addrb_14[13:0];
  assign sData_fire_15 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_14_ena = (_zz_ena_14[0] && sData_fire_15);
  assign mData_14 = xil_SimpleDualBram_14_doutb;
  assign xil_SimpleDualBram_15_addra = _zz_addra_15[10:0];
  assign xil_SimpleDualBram_15_addrb = _zz_addrb_15[13:0];
  assign sData_fire_16 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_15_ena = (_zz_ena_15[0] && sData_fire_16);
  assign mData_15 = xil_SimpleDualBram_15_doutb;
  assign xil_SimpleDualBram_16_addra = _zz_addra_16[10:0];
  assign xil_SimpleDualBram_16_addrb = _zz_addrb_16[13:0];
  assign sData_fire_17 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_16_ena = (_zz_ena_16[0] && sData_fire_17);
  assign mData_16 = xil_SimpleDualBram_16_doutb;
  assign xil_SimpleDualBram_17_addra = _zz_addra_17[10:0];
  assign xil_SimpleDualBram_17_addrb = _zz_addrb_17[13:0];
  assign sData_fire_18 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_17_ena = (_zz_ena_17[0] && sData_fire_18);
  assign mData_17 = xil_SimpleDualBram_17_doutb;
  assign xil_SimpleDualBram_18_addra = _zz_addra_18[10:0];
  assign xil_SimpleDualBram_18_addrb = _zz_addrb_18[13:0];
  assign sData_fire_19 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_18_ena = (_zz_ena_18[0] && sData_fire_19);
  assign mData_18 = xil_SimpleDualBram_18_doutb;
  assign xil_SimpleDualBram_19_addra = _zz_addra_19[10:0];
  assign xil_SimpleDualBram_19_addrb = _zz_addrb_19[13:0];
  assign sData_fire_20 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_19_ena = (_zz_ena_19[0] && sData_fire_20);
  assign mData_19 = xil_SimpleDualBram_19_doutb;
  assign xil_SimpleDualBram_20_addra = _zz_addra_20[10:0];
  assign xil_SimpleDualBram_20_addrb = _zz_addrb_20[13:0];
  assign sData_fire_21 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_20_ena = (_zz_ena_20[0] && sData_fire_21);
  assign mData_20 = xil_SimpleDualBram_20_doutb;
  assign xil_SimpleDualBram_21_addra = _zz_addra_21[10:0];
  assign xil_SimpleDualBram_21_addrb = _zz_addrb_21[13:0];
  assign sData_fire_22 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_21_ena = (_zz_ena_21[0] && sData_fire_22);
  assign mData_21 = xil_SimpleDualBram_21_doutb;
  assign xil_SimpleDualBram_22_addra = _zz_addra_22[10:0];
  assign xil_SimpleDualBram_22_addrb = _zz_addrb_22[13:0];
  assign sData_fire_23 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_22_ena = (_zz_ena_22[0] && sData_fire_23);
  assign mData_22 = xil_SimpleDualBram_22_doutb;
  assign xil_SimpleDualBram_23_addra = _zz_addra_23[10:0];
  assign xil_SimpleDualBram_23_addrb = _zz_addrb_23[13:0];
  assign sData_fire_24 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_23_ena = (_zz_ena_23[0] && sData_fire_24);
  assign mData_23 = xil_SimpleDualBram_23_doutb;
  assign xil_SimpleDualBram_24_addra = _zz_addra_24[10:0];
  assign xil_SimpleDualBram_24_addrb = _zz_addrb_24[13:0];
  assign sData_fire_25 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_24_ena = (_zz_ena_24[0] && sData_fire_25);
  assign mData_24 = xil_SimpleDualBram_24_doutb;
  assign xil_SimpleDualBram_25_addra = _zz_addra_25[10:0];
  assign xil_SimpleDualBram_25_addrb = _zz_addrb_25[13:0];
  assign sData_fire_26 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_25_ena = (_zz_ena_25[0] && sData_fire_26);
  assign mData_25 = xil_SimpleDualBram_25_doutb;
  assign xil_SimpleDualBram_26_addra = _zz_addra_26[10:0];
  assign xil_SimpleDualBram_26_addrb = _zz_addrb_26[13:0];
  assign sData_fire_27 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_26_ena = (_zz_ena_26[0] && sData_fire_27);
  assign mData_26 = xil_SimpleDualBram_26_doutb;
  assign xil_SimpleDualBram_27_addra = _zz_addra_27[10:0];
  assign xil_SimpleDualBram_27_addrb = _zz_addrb_27[13:0];
  assign sData_fire_28 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_27_ena = (_zz_ena_27[0] && sData_fire_28);
  assign mData_27 = xil_SimpleDualBram_27_doutb;
  assign xil_SimpleDualBram_28_addra = _zz_addra_28[10:0];
  assign xil_SimpleDualBram_28_addrb = _zz_addrb_28[13:0];
  assign sData_fire_29 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_28_ena = (_zz_ena_28[0] && sData_fire_29);
  assign mData_28 = xil_SimpleDualBram_28_doutb;
  assign xil_SimpleDualBram_29_addra = _zz_addra_29[10:0];
  assign xil_SimpleDualBram_29_addrb = _zz_addrb_29[13:0];
  assign sData_fire_30 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_29_ena = (_zz_ena_29[0] && sData_fire_30);
  assign mData_29 = xil_SimpleDualBram_29_doutb;
  assign xil_SimpleDualBram_30_addra = _zz_addra_30[10:0];
  assign xil_SimpleDualBram_30_addrb = _zz_addrb_30[13:0];
  assign sData_fire_31 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_30_ena = (_zz_ena_30[0] && sData_fire_31);
  assign mData_30 = xil_SimpleDualBram_30_doutb;
  assign xil_SimpleDualBram_31_addra = _zz_addra_31[10:0];
  assign xil_SimpleDualBram_31_addrb = _zz_addrb_31[13:0];
  assign sData_fire_32 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_31_ena = (_zz_ena_31[0] && sData_fire_32);
  assign mData_31 = xil_SimpleDualBram_31_doutb;
  assign xil_SimpleDualBram_32_addra = _zz_addra_32[10:0];
  assign xil_SimpleDualBram_32_addrb = _zz_addrb_32[13:0];
  assign sData_fire_33 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_32_ena = (_zz_ena_32[0] && sData_fire_33);
  assign mData_32 = xil_SimpleDualBram_32_doutb;
  assign xil_SimpleDualBram_33_addra = _zz_addra_33[10:0];
  assign xil_SimpleDualBram_33_addrb = _zz_addrb_33[13:0];
  assign sData_fire_34 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_33_ena = (_zz_ena_33[0] && sData_fire_34);
  assign mData_33 = xil_SimpleDualBram_33_doutb;
  assign xil_SimpleDualBram_34_addra = _zz_addra_34[10:0];
  assign xil_SimpleDualBram_34_addrb = _zz_addrb_34[13:0];
  assign sData_fire_35 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_34_ena = (_zz_ena_34[0] && sData_fire_35);
  assign mData_34 = xil_SimpleDualBram_34_doutb;
  assign xil_SimpleDualBram_35_addra = _zz_addra_35[10:0];
  assign xil_SimpleDualBram_35_addrb = _zz_addrb_35[13:0];
  assign sData_fire_36 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_35_ena = (_zz_ena_35[0] && sData_fire_36);
  assign mData_35 = xil_SimpleDualBram_35_doutb;
  assign xil_SimpleDualBram_36_addra = _zz_addra_36[10:0];
  assign xil_SimpleDualBram_36_addrb = _zz_addrb_36[13:0];
  assign sData_fire_37 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_36_ena = (_zz_ena_36[0] && sData_fire_37);
  assign mData_36 = xil_SimpleDualBram_36_doutb;
  assign xil_SimpleDualBram_37_addra = _zz_addra_37[10:0];
  assign xil_SimpleDualBram_37_addrb = _zz_addrb_37[13:0];
  assign sData_fire_38 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_37_ena = (_zz_ena_37[0] && sData_fire_38);
  assign mData_37 = xil_SimpleDualBram_37_doutb;
  assign xil_SimpleDualBram_38_addra = _zz_addra_38[10:0];
  assign xil_SimpleDualBram_38_addrb = _zz_addrb_38[13:0];
  assign sData_fire_39 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_38_ena = (_zz_ena_38[0] && sData_fire_39);
  assign mData_38 = xil_SimpleDualBram_38_doutb;
  assign xil_SimpleDualBram_39_addra = _zz_addra_39[10:0];
  assign xil_SimpleDualBram_39_addrb = _zz_addrb_39[13:0];
  assign sData_fire_40 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_39_ena = (_zz_ena_39[0] && sData_fire_40);
  assign mData_39 = xil_SimpleDualBram_39_doutb;
  assign xil_SimpleDualBram_40_addra = _zz_addra_40[10:0];
  assign xil_SimpleDualBram_40_addrb = _zz_addrb_40[13:0];
  assign sData_fire_41 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_40_ena = (_zz_ena_40[0] && sData_fire_41);
  assign mData_40 = xil_SimpleDualBram_40_doutb;
  assign xil_SimpleDualBram_41_addra = _zz_addra_41[10:0];
  assign xil_SimpleDualBram_41_addrb = _zz_addrb_41[13:0];
  assign sData_fire_42 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_41_ena = (_zz_ena_41[0] && sData_fire_42);
  assign mData_41 = xil_SimpleDualBram_41_doutb;
  assign xil_SimpleDualBram_42_addra = _zz_addra_42[10:0];
  assign xil_SimpleDualBram_42_addrb = _zz_addrb_42[13:0];
  assign sData_fire_43 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_42_ena = (_zz_ena_42[0] && sData_fire_43);
  assign mData_42 = xil_SimpleDualBram_42_doutb;
  assign xil_SimpleDualBram_43_addra = _zz_addra_43[10:0];
  assign xil_SimpleDualBram_43_addrb = _zz_addrb_43[13:0];
  assign sData_fire_44 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_43_ena = (_zz_ena_43[0] && sData_fire_44);
  assign mData_43 = xil_SimpleDualBram_43_doutb;
  assign xil_SimpleDualBram_44_addra = _zz_addra_44[10:0];
  assign xil_SimpleDualBram_44_addrb = _zz_addrb_44[13:0];
  assign sData_fire_45 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_44_ena = (_zz_ena_44[0] && sData_fire_45);
  assign mData_44 = xil_SimpleDualBram_44_doutb;
  assign xil_SimpleDualBram_45_addra = _zz_addra_45[10:0];
  assign xil_SimpleDualBram_45_addrb = _zz_addrb_45[13:0];
  assign sData_fire_46 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_45_ena = (_zz_ena_45[0] && sData_fire_46);
  assign mData_45 = xil_SimpleDualBram_45_doutb;
  assign xil_SimpleDualBram_46_addra = _zz_addra_46[10:0];
  assign xil_SimpleDualBram_46_addrb = _zz_addrb_46[13:0];
  assign sData_fire_47 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_46_ena = (_zz_ena_46[0] && sData_fire_47);
  assign mData_46 = xil_SimpleDualBram_46_doutb;
  assign xil_SimpleDualBram_47_addra = _zz_addra_47[10:0];
  assign xil_SimpleDualBram_47_addrb = _zz_addrb_47[13:0];
  assign sData_fire_48 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_47_ena = (_zz_ena_47[0] && sData_fire_48);
  assign mData_47 = xil_SimpleDualBram_47_doutb;
  assign xil_SimpleDualBram_48_addra = _zz_addra_48[10:0];
  assign xil_SimpleDualBram_48_addrb = _zz_addrb_48[13:0];
  assign sData_fire_49 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_48_ena = (_zz_ena_48[0] && sData_fire_49);
  assign mData_48 = xil_SimpleDualBram_48_doutb;
  assign xil_SimpleDualBram_49_addra = _zz_addra_49[10:0];
  assign xil_SimpleDualBram_49_addrb = _zz_addrb_49[13:0];
  assign sData_fire_50 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_49_ena = (_zz_ena_49[0] && sData_fire_50);
  assign mData_49 = xil_SimpleDualBram_49_doutb;
  assign xil_SimpleDualBram_50_addra = _zz_addra_50[10:0];
  assign xil_SimpleDualBram_50_addrb = _zz_addrb_50[13:0];
  assign sData_fire_51 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_50_ena = (_zz_ena_50[0] && sData_fire_51);
  assign mData_50 = xil_SimpleDualBram_50_doutb;
  assign xil_SimpleDualBram_51_addra = _zz_addra_51[10:0];
  assign xil_SimpleDualBram_51_addrb = _zz_addrb_51[13:0];
  assign sData_fire_52 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_51_ena = (_zz_ena_51[0] && sData_fire_52);
  assign mData_51 = xil_SimpleDualBram_51_doutb;
  assign xil_SimpleDualBram_52_addra = _zz_addra_52[10:0];
  assign xil_SimpleDualBram_52_addrb = _zz_addrb_52[13:0];
  assign sData_fire_53 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_52_ena = (_zz_ena_52[0] && sData_fire_53);
  assign mData_52 = xil_SimpleDualBram_52_doutb;
  assign xil_SimpleDualBram_53_addra = _zz_addra_53[10:0];
  assign xil_SimpleDualBram_53_addrb = _zz_addrb_53[13:0];
  assign sData_fire_54 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_53_ena = (_zz_ena_53[0] && sData_fire_54);
  assign mData_53 = xil_SimpleDualBram_53_doutb;
  assign xil_SimpleDualBram_54_addra = _zz_addra_54[10:0];
  assign xil_SimpleDualBram_54_addrb = _zz_addrb_54[13:0];
  assign sData_fire_55 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_54_ena = (_zz_ena_54[0] && sData_fire_55);
  assign mData_54 = xil_SimpleDualBram_54_doutb;
  assign xil_SimpleDualBram_55_addra = _zz_addra_55[10:0];
  assign xil_SimpleDualBram_55_addrb = _zz_addrb_55[13:0];
  assign sData_fire_56 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_55_ena = (_zz_ena_55[0] && sData_fire_56);
  assign mData_55 = xil_SimpleDualBram_55_doutb;
  assign xil_SimpleDualBram_56_addra = _zz_addra_56[10:0];
  assign xil_SimpleDualBram_56_addrb = _zz_addrb_56[13:0];
  assign sData_fire_57 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_56_ena = (_zz_ena_56[0] && sData_fire_57);
  assign mData_56 = xil_SimpleDualBram_56_doutb;
  assign xil_SimpleDualBram_57_addra = _zz_addra_57[10:0];
  assign xil_SimpleDualBram_57_addrb = _zz_addrb_57[13:0];
  assign sData_fire_58 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_57_ena = (_zz_ena_57[0] && sData_fire_58);
  assign mData_57 = xil_SimpleDualBram_57_doutb;
  assign xil_SimpleDualBram_58_addra = _zz_addra_58[10:0];
  assign xil_SimpleDualBram_58_addrb = _zz_addrb_58[13:0];
  assign sData_fire_59 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_58_ena = (_zz_ena_58[0] && sData_fire_59);
  assign mData_58 = xil_SimpleDualBram_58_doutb;
  assign xil_SimpleDualBram_59_addra = _zz_addra_59[10:0];
  assign xil_SimpleDualBram_59_addrb = _zz_addrb_59[13:0];
  assign sData_fire_60 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_59_ena = (_zz_ena_59[0] && sData_fire_60);
  assign mData_59 = xil_SimpleDualBram_59_doutb;
  assign xil_SimpleDualBram_60_addra = _zz_addra_60[10:0];
  assign xil_SimpleDualBram_60_addrb = _zz_addrb_60[13:0];
  assign sData_fire_61 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_60_ena = (_zz_ena_60[0] && sData_fire_61);
  assign mData_60 = xil_SimpleDualBram_60_doutb;
  assign xil_SimpleDualBram_61_addra = _zz_addra_61[10:0];
  assign xil_SimpleDualBram_61_addrb = _zz_addrb_61[13:0];
  assign sData_fire_62 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_61_ena = (_zz_ena_61[0] && sData_fire_62);
  assign mData_61 = xil_SimpleDualBram_61_doutb;
  assign xil_SimpleDualBram_62_addra = _zz_addra_62[10:0];
  assign xil_SimpleDualBram_62_addrb = _zz_addrb_62[13:0];
  assign sData_fire_63 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_62_ena = (_zz_ena_62[0] && sData_fire_63);
  assign mData_62 = xil_SimpleDualBram_62_doutb;
  assign xil_SimpleDualBram_63_addra = _zz_addra_63[10:0];
  assign xil_SimpleDualBram_63_addrb = _zz_addrb_63[13:0];
  assign sData_fire_64 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_63_ena = (_zz_ena_63[0] && sData_fire_64);
  assign mData_63 = xil_SimpleDualBram_63_doutb;
  assign xil_SimpleDualBram_64_addra = _zz_addra_64[10:0];
  assign xil_SimpleDualBram_64_addrb = _zz_addrb_64[13:0];
  assign sData_fire_65 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_64_ena = (_zz_ena_64[0] && sData_fire_65);
  assign mData_64 = xil_SimpleDualBram_64_doutb;
  assign xil_SimpleDualBram_65_addra = _zz_addra_65[10:0];
  assign xil_SimpleDualBram_65_addrb = _zz_addrb_65[13:0];
  assign sData_fire_66 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_65_ena = (_zz_ena_65[0] && sData_fire_66);
  assign mData_65 = xil_SimpleDualBram_65_doutb;
  assign xil_SimpleDualBram_66_addra = _zz_addra_66[10:0];
  assign xil_SimpleDualBram_66_addrb = _zz_addrb_66[13:0];
  assign sData_fire_67 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_66_ena = (_zz_ena_66[0] && sData_fire_67);
  assign mData_66 = xil_SimpleDualBram_66_doutb;
  assign xil_SimpleDualBram_67_addra = _zz_addra_67[10:0];
  assign xil_SimpleDualBram_67_addrb = _zz_addrb_67[13:0];
  assign sData_fire_68 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_67_ena = (_zz_ena_67[0] && sData_fire_68);
  assign mData_67 = xil_SimpleDualBram_67_doutb;
  assign xil_SimpleDualBram_68_addra = _zz_addra_68[10:0];
  assign xil_SimpleDualBram_68_addrb = _zz_addrb_68[13:0];
  assign sData_fire_69 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_68_ena = (_zz_ena_68[0] && sData_fire_69);
  assign mData_68 = xil_SimpleDualBram_68_doutb;
  assign xil_SimpleDualBram_69_addra = _zz_addra_69[10:0];
  assign xil_SimpleDualBram_69_addrb = _zz_addrb_69[13:0];
  assign sData_fire_70 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_69_ena = (_zz_ena_69[0] && sData_fire_70);
  assign mData_69 = xil_SimpleDualBram_69_doutb;
  assign xil_SimpleDualBram_70_addra = _zz_addra_70[10:0];
  assign xil_SimpleDualBram_70_addrb = _zz_addrb_70[13:0];
  assign sData_fire_71 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_70_ena = (_zz_ena_70[0] && sData_fire_71);
  assign mData_70 = xil_SimpleDualBram_70_doutb;
  assign xil_SimpleDualBram_71_addra = _zz_addra_71[10:0];
  assign xil_SimpleDualBram_71_addrb = _zz_addrb_71[13:0];
  assign sData_fire_72 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_71_ena = (_zz_ena_71[0] && sData_fire_72);
  assign mData_71 = xil_SimpleDualBram_71_doutb;
  assign xil_SimpleDualBram_72_addra = _zz_addra_72[10:0];
  assign xil_SimpleDualBram_72_addrb = _zz_addrb_72[13:0];
  assign sData_fire_73 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_72_ena = (_zz_ena_72[0] && sData_fire_73);
  assign mData_72 = xil_SimpleDualBram_72_doutb;
  assign xil_SimpleDualBram_73_addra = _zz_addra_73[10:0];
  assign xil_SimpleDualBram_73_addrb = _zz_addrb_73[13:0];
  assign sData_fire_74 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_73_ena = (_zz_ena_73[0] && sData_fire_74);
  assign mData_73 = xil_SimpleDualBram_73_doutb;
  assign xil_SimpleDualBram_74_addra = _zz_addra_74[10:0];
  assign xil_SimpleDualBram_74_addrb = _zz_addrb_74[13:0];
  assign sData_fire_75 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_74_ena = (_zz_ena_74[0] && sData_fire_75);
  assign mData_74 = xil_SimpleDualBram_74_doutb;
  assign xil_SimpleDualBram_75_addra = _zz_addra_75[10:0];
  assign xil_SimpleDualBram_75_addrb = _zz_addrb_75[13:0];
  assign sData_fire_76 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_75_ena = (_zz_ena_75[0] && sData_fire_76);
  assign mData_75 = xil_SimpleDualBram_75_doutb;
  assign xil_SimpleDualBram_76_addra = _zz_addra_76[10:0];
  assign xil_SimpleDualBram_76_addrb = _zz_addrb_76[13:0];
  assign sData_fire_77 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_76_ena = (_zz_ena_76[0] && sData_fire_77);
  assign mData_76 = xil_SimpleDualBram_76_doutb;
  assign xil_SimpleDualBram_77_addra = _zz_addra_77[10:0];
  assign xil_SimpleDualBram_77_addrb = _zz_addrb_77[13:0];
  assign sData_fire_78 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_77_ena = (_zz_ena_77[0] && sData_fire_78);
  assign mData_77 = xil_SimpleDualBram_77_doutb;
  assign xil_SimpleDualBram_78_addra = _zz_addra_78[10:0];
  assign xil_SimpleDualBram_78_addrb = _zz_addrb_78[13:0];
  assign sData_fire_79 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_78_ena = (_zz_ena_78[0] && sData_fire_79);
  assign mData_78 = xil_SimpleDualBram_78_doutb;
  assign xil_SimpleDualBram_79_addra = _zz_addra_79[10:0];
  assign xil_SimpleDualBram_79_addrb = _zz_addrb_79[13:0];
  assign sData_fire_80 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_79_ena = (_zz_ena_79[0] && sData_fire_80);
  assign mData_79 = xil_SimpleDualBram_79_doutb;
  assign xil_SimpleDualBram_80_addra = _zz_addra_80[10:0];
  assign xil_SimpleDualBram_80_addrb = _zz_addrb_80[13:0];
  assign sData_fire_81 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_80_ena = (_zz_ena_80[0] && sData_fire_81);
  assign mData_80 = xil_SimpleDualBram_80_doutb;
  assign xil_SimpleDualBram_81_addra = _zz_addra_81[10:0];
  assign xil_SimpleDualBram_81_addrb = _zz_addrb_81[13:0];
  assign sData_fire_82 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_81_ena = (_zz_ena_81[0] && sData_fire_82);
  assign mData_81 = xil_SimpleDualBram_81_doutb;
  assign xil_SimpleDualBram_82_addra = _zz_addra_82[10:0];
  assign xil_SimpleDualBram_82_addrb = _zz_addrb_82[13:0];
  assign sData_fire_83 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_82_ena = (_zz_ena_82[0] && sData_fire_83);
  assign mData_82 = xil_SimpleDualBram_82_doutb;
  assign xil_SimpleDualBram_83_addra = _zz_addra_83[10:0];
  assign xil_SimpleDualBram_83_addrb = _zz_addrb_83[13:0];
  assign sData_fire_84 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_83_ena = (_zz_ena_83[0] && sData_fire_84);
  assign mData_83 = xil_SimpleDualBram_83_doutb;
  assign xil_SimpleDualBram_84_addra = _zz_addra_84[10:0];
  assign xil_SimpleDualBram_84_addrb = _zz_addrb_84[13:0];
  assign sData_fire_85 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_84_ena = (_zz_ena_84[0] && sData_fire_85);
  assign mData_84 = xil_SimpleDualBram_84_doutb;
  assign xil_SimpleDualBram_85_addra = _zz_addra_85[10:0];
  assign xil_SimpleDualBram_85_addrb = _zz_addrb_85[13:0];
  assign sData_fire_86 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_85_ena = (_zz_ena_85[0] && sData_fire_86);
  assign mData_85 = xil_SimpleDualBram_85_doutb;
  assign xil_SimpleDualBram_86_addra = _zz_addra_86[10:0];
  assign xil_SimpleDualBram_86_addrb = _zz_addrb_86[13:0];
  assign sData_fire_87 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_86_ena = (_zz_ena_86[0] && sData_fire_87);
  assign mData_86 = xil_SimpleDualBram_86_doutb;
  assign xil_SimpleDualBram_87_addra = _zz_addra_87[10:0];
  assign xil_SimpleDualBram_87_addrb = _zz_addrb_87[13:0];
  assign sData_fire_88 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_87_ena = (_zz_ena_87[0] && sData_fire_88);
  assign mData_87 = xil_SimpleDualBram_87_doutb;
  assign xil_SimpleDualBram_88_addra = _zz_addra_88[10:0];
  assign xil_SimpleDualBram_88_addrb = _zz_addrb_88[13:0];
  assign sData_fire_89 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_88_ena = (_zz_ena_88[0] && sData_fire_89);
  assign mData_88 = xil_SimpleDualBram_88_doutb;
  assign xil_SimpleDualBram_89_addra = _zz_addra_89[10:0];
  assign xil_SimpleDualBram_89_addrb = _zz_addrb_89[13:0];
  assign sData_fire_90 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_89_ena = (_zz_ena_89[0] && sData_fire_90);
  assign mData_89 = xil_SimpleDualBram_89_doutb;
  assign xil_SimpleDualBram_90_addra = _zz_addra_90[10:0];
  assign xil_SimpleDualBram_90_addrb = _zz_addrb_90[13:0];
  assign sData_fire_91 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_90_ena = (_zz_ena_90[0] && sData_fire_91);
  assign mData_90 = xil_SimpleDualBram_90_doutb;
  assign xil_SimpleDualBram_91_addra = _zz_addra_91[10:0];
  assign xil_SimpleDualBram_91_addrb = _zz_addrb_91[13:0];
  assign sData_fire_92 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_91_ena = (_zz_ena_91[0] && sData_fire_92);
  assign mData_91 = xil_SimpleDualBram_91_doutb;
  assign xil_SimpleDualBram_92_addra = _zz_addra_92[10:0];
  assign xil_SimpleDualBram_92_addrb = _zz_addrb_92[13:0];
  assign sData_fire_93 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_92_ena = (_zz_ena_92[0] && sData_fire_93);
  assign mData_92 = xil_SimpleDualBram_92_doutb;
  assign xil_SimpleDualBram_93_addra = _zz_addra_93[10:0];
  assign xil_SimpleDualBram_93_addrb = _zz_addrb_93[13:0];
  assign sData_fire_94 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_93_ena = (_zz_ena_93[0] && sData_fire_94);
  assign mData_93 = xil_SimpleDualBram_93_doutb;
  assign xil_SimpleDualBram_94_addra = _zz_addra_94[10:0];
  assign xil_SimpleDualBram_94_addrb = _zz_addrb_94[13:0];
  assign sData_fire_95 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_94_ena = (_zz_ena_94[0] && sData_fire_95);
  assign mData_94 = xil_SimpleDualBram_94_doutb;
  assign xil_SimpleDualBram_95_addra = _zz_addra_95[10:0];
  assign xil_SimpleDualBram_95_addrb = _zz_addrb_95[13:0];
  assign sData_fire_96 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_95_ena = (_zz_ena_95[0] && sData_fire_96);
  assign mData_95 = xil_SimpleDualBram_95_doutb;
  assign xil_SimpleDualBram_96_addra = _zz_addra_96[10:0];
  assign xil_SimpleDualBram_96_addrb = _zz_addrb_96[13:0];
  assign sData_fire_97 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_96_ena = (_zz_ena_96[0] && sData_fire_97);
  assign mData_96 = xil_SimpleDualBram_96_doutb;
  assign xil_SimpleDualBram_97_addra = _zz_addra_97[10:0];
  assign xil_SimpleDualBram_97_addrb = _zz_addrb_97[13:0];
  assign sData_fire_98 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_97_ena = (_zz_ena_97[0] && sData_fire_98);
  assign mData_97 = xil_SimpleDualBram_97_doutb;
  assign xil_SimpleDualBram_98_addra = _zz_addra_98[10:0];
  assign xil_SimpleDualBram_98_addrb = _zz_addrb_98[13:0];
  assign sData_fire_99 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_98_ena = (_zz_ena_98[0] && sData_fire_99);
  assign mData_98 = xil_SimpleDualBram_98_doutb;
  assign xil_SimpleDualBram_99_addra = _zz_addra_99[10:0];
  assign xil_SimpleDualBram_99_addrb = _zz_addrb_99[13:0];
  assign sData_fire_100 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_99_ena = (_zz_ena_99[0] && sData_fire_100);
  assign mData_99 = xil_SimpleDualBram_99_doutb;
  assign xil_SimpleDualBram_100_addra = _zz_addra_100[10:0];
  assign xil_SimpleDualBram_100_addrb = _zz_addrb_100[13:0];
  assign sData_fire_101 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_100_ena = (_zz_ena_100[0] && sData_fire_101);
  assign mData_100 = xil_SimpleDualBram_100_doutb;
  assign xil_SimpleDualBram_101_addra = _zz_addra_101[10:0];
  assign xil_SimpleDualBram_101_addrb = _zz_addrb_101[13:0];
  assign sData_fire_102 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_101_ena = (_zz_ena_101[0] && sData_fire_102);
  assign mData_101 = xil_SimpleDualBram_101_doutb;
  assign xil_SimpleDualBram_102_addra = _zz_addra_102[10:0];
  assign xil_SimpleDualBram_102_addrb = _zz_addrb_102[13:0];
  assign sData_fire_103 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_102_ena = (_zz_ena_102[0] && sData_fire_103);
  assign mData_102 = xil_SimpleDualBram_102_doutb;
  assign xil_SimpleDualBram_103_addra = _zz_addra_103[10:0];
  assign xil_SimpleDualBram_103_addrb = _zz_addrb_103[13:0];
  assign sData_fire_104 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_103_ena = (_zz_ena_103[0] && sData_fire_104);
  assign mData_103 = xil_SimpleDualBram_103_doutb;
  assign xil_SimpleDualBram_104_addra = _zz_addra_104[10:0];
  assign xil_SimpleDualBram_104_addrb = _zz_addrb_104[13:0];
  assign sData_fire_105 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_104_ena = (_zz_ena_104[0] && sData_fire_105);
  assign mData_104 = xil_SimpleDualBram_104_doutb;
  assign xil_SimpleDualBram_105_addra = _zz_addra_105[10:0];
  assign xil_SimpleDualBram_105_addrb = _zz_addrb_105[13:0];
  assign sData_fire_106 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_105_ena = (_zz_ena_105[0] && sData_fire_106);
  assign mData_105 = xil_SimpleDualBram_105_doutb;
  assign xil_SimpleDualBram_106_addra = _zz_addra_106[10:0];
  assign xil_SimpleDualBram_106_addrb = _zz_addrb_106[13:0];
  assign sData_fire_107 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_106_ena = (_zz_ena_106[0] && sData_fire_107);
  assign mData_106 = xil_SimpleDualBram_106_doutb;
  assign xil_SimpleDualBram_107_addra = _zz_addra_107[10:0];
  assign xil_SimpleDualBram_107_addrb = _zz_addrb_107[13:0];
  assign sData_fire_108 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_107_ena = (_zz_ena_107[0] && sData_fire_108);
  assign mData_107 = xil_SimpleDualBram_107_doutb;
  assign xil_SimpleDualBram_108_addra = _zz_addra_108[10:0];
  assign xil_SimpleDualBram_108_addrb = _zz_addrb_108[13:0];
  assign sData_fire_109 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_108_ena = (_zz_ena_108[0] && sData_fire_109);
  assign mData_108 = xil_SimpleDualBram_108_doutb;
  assign xil_SimpleDualBram_109_addra = _zz_addra_109[10:0];
  assign xil_SimpleDualBram_109_addrb = _zz_addrb_109[13:0];
  assign sData_fire_110 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_109_ena = (_zz_ena_109[0] && sData_fire_110);
  assign mData_109 = xil_SimpleDualBram_109_doutb;
  assign xil_SimpleDualBram_110_addra = _zz_addra_110[10:0];
  assign xil_SimpleDualBram_110_addrb = _zz_addrb_110[13:0];
  assign sData_fire_111 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_110_ena = (_zz_ena_110[0] && sData_fire_111);
  assign mData_110 = xil_SimpleDualBram_110_doutb;
  assign xil_SimpleDualBram_111_addra = _zz_addra_111[10:0];
  assign xil_SimpleDualBram_111_addrb = _zz_addrb_111[13:0];
  assign sData_fire_112 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_111_ena = (_zz_ena_111[0] && sData_fire_112);
  assign mData_111 = xil_SimpleDualBram_111_doutb;
  assign xil_SimpleDualBram_112_addra = _zz_addra_112[10:0];
  assign xil_SimpleDualBram_112_addrb = _zz_addrb_112[13:0];
  assign sData_fire_113 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_112_ena = (_zz_ena_112[0] && sData_fire_113);
  assign mData_112 = xil_SimpleDualBram_112_doutb;
  assign xil_SimpleDualBram_113_addra = _zz_addra_113[10:0];
  assign xil_SimpleDualBram_113_addrb = _zz_addrb_113[13:0];
  assign sData_fire_114 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_113_ena = (_zz_ena_113[0] && sData_fire_114);
  assign mData_113 = xil_SimpleDualBram_113_doutb;
  assign xil_SimpleDualBram_114_addra = _zz_addra_114[10:0];
  assign xil_SimpleDualBram_114_addrb = _zz_addrb_114[13:0];
  assign sData_fire_115 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_114_ena = (_zz_ena_114[0] && sData_fire_115);
  assign mData_114 = xil_SimpleDualBram_114_doutb;
  assign xil_SimpleDualBram_115_addra = _zz_addra_115[10:0];
  assign xil_SimpleDualBram_115_addrb = _zz_addrb_115[13:0];
  assign sData_fire_116 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_115_ena = (_zz_ena_115[0] && sData_fire_116);
  assign mData_115 = xil_SimpleDualBram_115_doutb;
  assign xil_SimpleDualBram_116_addra = _zz_addra_116[10:0];
  assign xil_SimpleDualBram_116_addrb = _zz_addrb_116[13:0];
  assign sData_fire_117 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_116_ena = (_zz_ena_116[0] && sData_fire_117);
  assign mData_116 = xil_SimpleDualBram_116_doutb;
  assign xil_SimpleDualBram_117_addra = _zz_addra_117[10:0];
  assign xil_SimpleDualBram_117_addrb = _zz_addrb_117[13:0];
  assign sData_fire_118 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_117_ena = (_zz_ena_117[0] && sData_fire_118);
  assign mData_117 = xil_SimpleDualBram_117_doutb;
  assign xil_SimpleDualBram_118_addra = _zz_addra_118[10:0];
  assign xil_SimpleDualBram_118_addrb = _zz_addrb_118[13:0];
  assign sData_fire_119 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_118_ena = (_zz_ena_118[0] && sData_fire_119);
  assign mData_118 = xil_SimpleDualBram_118_doutb;
  assign xil_SimpleDualBram_119_addra = _zz_addra_119[10:0];
  assign xil_SimpleDualBram_119_addrb = _zz_addrb_119[13:0];
  assign sData_fire_120 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_119_ena = (_zz_ena_119[0] && sData_fire_120);
  assign mData_119 = xil_SimpleDualBram_119_doutb;
  assign xil_SimpleDualBram_120_addra = _zz_addra_120[10:0];
  assign xil_SimpleDualBram_120_addrb = _zz_addrb_120[13:0];
  assign sData_fire_121 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_120_ena = (_zz_ena_120[0] && sData_fire_121);
  assign mData_120 = xil_SimpleDualBram_120_doutb;
  assign xil_SimpleDualBram_121_addra = _zz_addra_121[10:0];
  assign xil_SimpleDualBram_121_addrb = _zz_addrb_121[13:0];
  assign sData_fire_122 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_121_ena = (_zz_ena_121[0] && sData_fire_122);
  assign mData_121 = xil_SimpleDualBram_121_doutb;
  assign xil_SimpleDualBram_122_addra = _zz_addra_122[10:0];
  assign xil_SimpleDualBram_122_addrb = _zz_addrb_122[13:0];
  assign sData_fire_123 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_122_ena = (_zz_ena_122[0] && sData_fire_123);
  assign mData_122 = xil_SimpleDualBram_122_doutb;
  assign xil_SimpleDualBram_123_addra = _zz_addra_123[10:0];
  assign xil_SimpleDualBram_123_addrb = _zz_addrb_123[13:0];
  assign sData_fire_124 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_123_ena = (_zz_ena_123[0] && sData_fire_124);
  assign mData_123 = xil_SimpleDualBram_123_doutb;
  assign xil_SimpleDualBram_124_addra = _zz_addra_124[10:0];
  assign xil_SimpleDualBram_124_addrb = _zz_addrb_124[13:0];
  assign sData_fire_125 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_124_ena = (_zz_ena_124[0] && sData_fire_125);
  assign mData_124 = xil_SimpleDualBram_124_doutb;
  assign xil_SimpleDualBram_125_addra = _zz_addra_125[10:0];
  assign xil_SimpleDualBram_125_addrb = _zz_addrb_125[13:0];
  assign sData_fire_126 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_125_ena = (_zz_ena_125[0] && sData_fire_126);
  assign mData_125 = xil_SimpleDualBram_125_doutb;
  assign xil_SimpleDualBram_126_addra = _zz_addra_126[10:0];
  assign xil_SimpleDualBram_126_addrb = _zz_addrb_126[13:0];
  assign sData_fire_127 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_126_ena = (_zz_ena_126[0] && sData_fire_127);
  assign mData_126 = xil_SimpleDualBram_126_doutb;
  assign xil_SimpleDualBram_127_addra = _zz_addra_127[10:0];
  assign xil_SimpleDualBram_127_addrb = _zz_addrb_127[13:0];
  assign sData_fire_128 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_127_ena = (_zz_ena_127[0] && sData_fire_128);
  assign mData_127 = xil_SimpleDualBram_127_doutb;
  assign xil_SimpleDualBram_128_addra = _zz_addra_128[10:0];
  assign xil_SimpleDualBram_128_addrb = _zz_addrb_128[13:0];
  assign sData_fire_129 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_128_ena = (_zz_ena_128[0] && sData_fire_129);
  assign mData_128 = xil_SimpleDualBram_128_doutb;
  assign xil_SimpleDualBram_129_addra = _zz_addra_129[10:0];
  assign xil_SimpleDualBram_129_addrb = _zz_addrb_129[13:0];
  assign sData_fire_130 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_129_ena = (_zz_ena_129[0] && sData_fire_130);
  assign mData_129 = xil_SimpleDualBram_129_doutb;
  assign xil_SimpleDualBram_130_addra = _zz_addra_130[10:0];
  assign xil_SimpleDualBram_130_addrb = _zz_addrb_130[13:0];
  assign sData_fire_131 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_130_ena = (_zz_ena_130[0] && sData_fire_131);
  assign mData_130 = xil_SimpleDualBram_130_doutb;
  assign xil_SimpleDualBram_131_addra = _zz_addra_131[10:0];
  assign xil_SimpleDualBram_131_addrb = _zz_addrb_131[13:0];
  assign sData_fire_132 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_131_ena = (_zz_ena_131[0] && sData_fire_132);
  assign mData_131 = xil_SimpleDualBram_131_doutb;
  assign xil_SimpleDualBram_132_addra = _zz_addra_132[10:0];
  assign xil_SimpleDualBram_132_addrb = _zz_addrb_132[13:0];
  assign sData_fire_133 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_132_ena = (_zz_ena_132[0] && sData_fire_133);
  assign mData_132 = xil_SimpleDualBram_132_doutb;
  assign xil_SimpleDualBram_133_addra = _zz_addra_133[10:0];
  assign xil_SimpleDualBram_133_addrb = _zz_addrb_133[13:0];
  assign sData_fire_134 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_133_ena = (_zz_ena_133[0] && sData_fire_134);
  assign mData_133 = xil_SimpleDualBram_133_doutb;
  assign xil_SimpleDualBram_134_addra = _zz_addra_134[10:0];
  assign xil_SimpleDualBram_134_addrb = _zz_addrb_134[13:0];
  assign sData_fire_135 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_134_ena = (_zz_ena_134[0] && sData_fire_135);
  assign mData_134 = xil_SimpleDualBram_134_doutb;
  assign xil_SimpleDualBram_135_addra = _zz_addra_135[10:0];
  assign xil_SimpleDualBram_135_addrb = _zz_addrb_135[13:0];
  assign sData_fire_136 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_135_ena = (_zz_ena_135[0] && sData_fire_136);
  assign mData_135 = xil_SimpleDualBram_135_doutb;
  assign xil_SimpleDualBram_136_addra = _zz_addra_136[10:0];
  assign xil_SimpleDualBram_136_addrb = _zz_addrb_136[13:0];
  assign sData_fire_137 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_136_ena = (_zz_ena_136[0] && sData_fire_137);
  assign mData_136 = xil_SimpleDualBram_136_doutb;
  assign xil_SimpleDualBram_137_addra = _zz_addra_137[10:0];
  assign xil_SimpleDualBram_137_addrb = _zz_addrb_137[13:0];
  assign sData_fire_138 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_137_ena = (_zz_ena_137[0] && sData_fire_138);
  assign mData_137 = xil_SimpleDualBram_137_doutb;
  assign xil_SimpleDualBram_138_addra = _zz_addra_138[10:0];
  assign xil_SimpleDualBram_138_addrb = _zz_addrb_138[13:0];
  assign sData_fire_139 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_138_ena = (_zz_ena_138[0] && sData_fire_139);
  assign mData_138 = xil_SimpleDualBram_138_doutb;
  assign xil_SimpleDualBram_139_addra = _zz_addra_139[10:0];
  assign xil_SimpleDualBram_139_addrb = _zz_addrb_139[13:0];
  assign sData_fire_140 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_139_ena = (_zz_ena_139[0] && sData_fire_140);
  assign mData_139 = xil_SimpleDualBram_139_doutb;
  assign xil_SimpleDualBram_140_addra = _zz_addra_140[10:0];
  assign xil_SimpleDualBram_140_addrb = _zz_addrb_140[13:0];
  assign sData_fire_141 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_140_ena = (_zz_ena_140[0] && sData_fire_141);
  assign mData_140 = xil_SimpleDualBram_140_doutb;
  assign xil_SimpleDualBram_141_addra = _zz_addra_141[10:0];
  assign xil_SimpleDualBram_141_addrb = _zz_addrb_141[13:0];
  assign sData_fire_142 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_141_ena = (_zz_ena_141[0] && sData_fire_142);
  assign mData_141 = xil_SimpleDualBram_141_doutb;
  assign xil_SimpleDualBram_142_addra = _zz_addra_142[10:0];
  assign xil_SimpleDualBram_142_addrb = _zz_addrb_142[13:0];
  assign sData_fire_143 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_142_ena = (_zz_ena_142[0] && sData_fire_143);
  assign mData_142 = xil_SimpleDualBram_142_doutb;
  assign xil_SimpleDualBram_143_addra = _zz_addra_143[10:0];
  assign xil_SimpleDualBram_143_addrb = _zz_addrb_143[13:0];
  assign sData_fire_144 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_143_ena = (_zz_ena_143[0] && sData_fire_144);
  assign mData_143 = xil_SimpleDualBram_143_doutb;
  assign xil_SimpleDualBram_144_addra = _zz_addra_144[10:0];
  assign xil_SimpleDualBram_144_addrb = _zz_addrb_144[13:0];
  assign sData_fire_145 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_144_ena = (_zz_ena_144[0] && sData_fire_145);
  assign mData_144 = xil_SimpleDualBram_144_doutb;
  assign xil_SimpleDualBram_145_addra = _zz_addra_145[10:0];
  assign xil_SimpleDualBram_145_addrb = _zz_addrb_145[13:0];
  assign sData_fire_146 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_145_ena = (_zz_ena_145[0] && sData_fire_146);
  assign mData_145 = xil_SimpleDualBram_145_doutb;
  assign xil_SimpleDualBram_146_addra = _zz_addra_146[10:0];
  assign xil_SimpleDualBram_146_addrb = _zz_addrb_146[13:0];
  assign sData_fire_147 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_146_ena = (_zz_ena_146[0] && sData_fire_147);
  assign mData_146 = xil_SimpleDualBram_146_doutb;
  assign xil_SimpleDualBram_147_addra = _zz_addra_147[10:0];
  assign xil_SimpleDualBram_147_addrb = _zz_addrb_147[13:0];
  assign sData_fire_148 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_147_ena = (_zz_ena_147[0] && sData_fire_148);
  assign mData_147 = xil_SimpleDualBram_147_doutb;
  assign xil_SimpleDualBram_148_addra = _zz_addra_148[10:0];
  assign xil_SimpleDualBram_148_addrb = _zz_addrb_148[13:0];
  assign sData_fire_149 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_148_ena = (_zz_ena_148[0] && sData_fire_149);
  assign mData_148 = xil_SimpleDualBram_148_doutb;
  assign xil_SimpleDualBram_149_addra = _zz_addra_149[10:0];
  assign xil_SimpleDualBram_149_addrb = _zz_addrb_149[13:0];
  assign sData_fire_150 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_149_ena = (_zz_ena_149[0] && sData_fire_150);
  assign mData_149 = xil_SimpleDualBram_149_doutb;
  assign xil_SimpleDualBram_150_addra = _zz_addra_150[10:0];
  assign xil_SimpleDualBram_150_addrb = _zz_addrb_150[13:0];
  assign sData_fire_151 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_150_ena = (_zz_ena_150[0] && sData_fire_151);
  assign mData_150 = xil_SimpleDualBram_150_doutb;
  assign xil_SimpleDualBram_151_addra = _zz_addra_151[10:0];
  assign xil_SimpleDualBram_151_addrb = _zz_addrb_151[13:0];
  assign sData_fire_152 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_151_ena = (_zz_ena_151[0] && sData_fire_152);
  assign mData_151 = xil_SimpleDualBram_151_doutb;
  assign xil_SimpleDualBram_152_addra = _zz_addra_152[10:0];
  assign xil_SimpleDualBram_152_addrb = _zz_addrb_152[13:0];
  assign sData_fire_153 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_152_ena = (_zz_ena_152[0] && sData_fire_153);
  assign mData_152 = xil_SimpleDualBram_152_doutb;
  assign xil_SimpleDualBram_153_addra = _zz_addra_153[10:0];
  assign xil_SimpleDualBram_153_addrb = _zz_addrb_153[13:0];
  assign sData_fire_154 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_153_ena = (_zz_ena_153[0] && sData_fire_154);
  assign mData_153 = xil_SimpleDualBram_153_doutb;
  assign xil_SimpleDualBram_154_addra = _zz_addra_154[10:0];
  assign xil_SimpleDualBram_154_addrb = _zz_addrb_154[13:0];
  assign sData_fire_155 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_154_ena = (_zz_ena_154[0] && sData_fire_155);
  assign mData_154 = xil_SimpleDualBram_154_doutb;
  assign xil_SimpleDualBram_155_addra = _zz_addra_155[10:0];
  assign xil_SimpleDualBram_155_addrb = _zz_addrb_155[13:0];
  assign sData_fire_156 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_155_ena = (_zz_ena_155[0] && sData_fire_156);
  assign mData_155 = xil_SimpleDualBram_155_doutb;
  assign xil_SimpleDualBram_156_addra = _zz_addra_156[10:0];
  assign xil_SimpleDualBram_156_addrb = _zz_addrb_156[13:0];
  assign sData_fire_157 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_156_ena = (_zz_ena_156[0] && sData_fire_157);
  assign mData_156 = xil_SimpleDualBram_156_doutb;
  assign xil_SimpleDualBram_157_addra = _zz_addra_157[10:0];
  assign xil_SimpleDualBram_157_addrb = _zz_addrb_157[13:0];
  assign sData_fire_158 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_157_ena = (_zz_ena_157[0] && sData_fire_158);
  assign mData_157 = xil_SimpleDualBram_157_doutb;
  assign xil_SimpleDualBram_158_addra = _zz_addra_158[10:0];
  assign xil_SimpleDualBram_158_addrb = _zz_addrb_158[13:0];
  assign sData_fire_159 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_158_ena = (_zz_ena_158[0] && sData_fire_159);
  assign mData_158 = xil_SimpleDualBram_158_doutb;
  assign xil_SimpleDualBram_159_addra = _zz_addra_159[10:0];
  assign xil_SimpleDualBram_159_addrb = _zz_addrb_159[13:0];
  assign sData_fire_160 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_159_ena = (_zz_ena_159[0] && sData_fire_160);
  assign mData_159 = xil_SimpleDualBram_159_doutb;
  assign xil_SimpleDualBram_160_addra = _zz_addra_160[10:0];
  assign xil_SimpleDualBram_160_addrb = _zz_addrb_160[13:0];
  assign sData_fire_161 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_160_ena = (_zz_ena_160[0] && sData_fire_161);
  assign mData_160 = xil_SimpleDualBram_160_doutb;
  assign xil_SimpleDualBram_161_addra = _zz_addra_161[10:0];
  assign xil_SimpleDualBram_161_addrb = _zz_addrb_161[13:0];
  assign sData_fire_162 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_161_ena = (_zz_ena_161[0] && sData_fire_162);
  assign mData_161 = xil_SimpleDualBram_161_doutb;
  assign xil_SimpleDualBram_162_addra = _zz_addra_162[10:0];
  assign xil_SimpleDualBram_162_addrb = _zz_addrb_162[13:0];
  assign sData_fire_163 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_162_ena = (_zz_ena_162[0] && sData_fire_163);
  assign mData_162 = xil_SimpleDualBram_162_doutb;
  assign xil_SimpleDualBram_163_addra = _zz_addra_163[10:0];
  assign xil_SimpleDualBram_163_addrb = _zz_addrb_163[13:0];
  assign sData_fire_164 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_163_ena = (_zz_ena_163[0] && sData_fire_164);
  assign mData_163 = xil_SimpleDualBram_163_doutb;
  assign xil_SimpleDualBram_164_addra = _zz_addra_164[10:0];
  assign xil_SimpleDualBram_164_addrb = _zz_addrb_164[13:0];
  assign sData_fire_165 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_164_ena = (_zz_ena_164[0] && sData_fire_165);
  assign mData_164 = xil_SimpleDualBram_164_doutb;
  assign xil_SimpleDualBram_165_addra = _zz_addra_165[10:0];
  assign xil_SimpleDualBram_165_addrb = _zz_addrb_165[13:0];
  assign sData_fire_166 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_165_ena = (_zz_ena_165[0] && sData_fire_166);
  assign mData_165 = xil_SimpleDualBram_165_doutb;
  assign xil_SimpleDualBram_166_addra = _zz_addra_166[10:0];
  assign xil_SimpleDualBram_166_addrb = _zz_addrb_166[13:0];
  assign sData_fire_167 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_166_ena = (_zz_ena_166[0] && sData_fire_167);
  assign mData_166 = xil_SimpleDualBram_166_doutb;
  assign xil_SimpleDualBram_167_addra = _zz_addra_167[10:0];
  assign xil_SimpleDualBram_167_addrb = _zz_addrb_167[13:0];
  assign sData_fire_168 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_167_ena = (_zz_ena_167[0] && sData_fire_168);
  assign mData_167 = xil_SimpleDualBram_167_doutb;
  assign xil_SimpleDualBram_168_addra = _zz_addra_168[10:0];
  assign xil_SimpleDualBram_168_addrb = _zz_addrb_168[13:0];
  assign sData_fire_169 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_168_ena = (_zz_ena_168[0] && sData_fire_169);
  assign mData_168 = xil_SimpleDualBram_168_doutb;
  assign xil_SimpleDualBram_169_addra = _zz_addra_169[10:0];
  assign xil_SimpleDualBram_169_addrb = _zz_addrb_169[13:0];
  assign sData_fire_170 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_169_ena = (_zz_ena_169[0] && sData_fire_170);
  assign mData_169 = xil_SimpleDualBram_169_doutb;
  assign xil_SimpleDualBram_170_addra = _zz_addra_170[10:0];
  assign xil_SimpleDualBram_170_addrb = _zz_addrb_170[13:0];
  assign sData_fire_171 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_170_ena = (_zz_ena_170[0] && sData_fire_171);
  assign mData_170 = xil_SimpleDualBram_170_doutb;
  assign xil_SimpleDualBram_171_addra = _zz_addra_171[10:0];
  assign xil_SimpleDualBram_171_addrb = _zz_addrb_171[13:0];
  assign sData_fire_172 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_171_ena = (_zz_ena_171[0] && sData_fire_172);
  assign mData_171 = xil_SimpleDualBram_171_doutb;
  assign xil_SimpleDualBram_172_addra = _zz_addra_172[10:0];
  assign xil_SimpleDualBram_172_addrb = _zz_addrb_172[13:0];
  assign sData_fire_173 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_172_ena = (_zz_ena_172[0] && sData_fire_173);
  assign mData_172 = xil_SimpleDualBram_172_doutb;
  assign xil_SimpleDualBram_173_addra = _zz_addra_173[10:0];
  assign xil_SimpleDualBram_173_addrb = _zz_addrb_173[13:0];
  assign sData_fire_174 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_173_ena = (_zz_ena_173[0] && sData_fire_174);
  assign mData_173 = xil_SimpleDualBram_173_doutb;
  assign xil_SimpleDualBram_174_addra = _zz_addra_174[10:0];
  assign xil_SimpleDualBram_174_addrb = _zz_addrb_174[13:0];
  assign sData_fire_175 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_174_ena = (_zz_ena_174[0] && sData_fire_175);
  assign mData_174 = xil_SimpleDualBram_174_doutb;
  assign xil_SimpleDualBram_175_addra = _zz_addra_175[10:0];
  assign xil_SimpleDualBram_175_addrb = _zz_addrb_175[13:0];
  assign sData_fire_176 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_175_ena = (_zz_ena_175[0] && sData_fire_176);
  assign mData_175 = xil_SimpleDualBram_175_doutb;
  assign xil_SimpleDualBram_176_addra = _zz_addra_176[10:0];
  assign xil_SimpleDualBram_176_addrb = _zz_addrb_176[13:0];
  assign sData_fire_177 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_176_ena = (_zz_ena_176[0] && sData_fire_177);
  assign mData_176 = xil_SimpleDualBram_176_doutb;
  assign xil_SimpleDualBram_177_addra = _zz_addra_177[10:0];
  assign xil_SimpleDualBram_177_addrb = _zz_addrb_177[13:0];
  assign sData_fire_178 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_177_ena = (_zz_ena_177[0] && sData_fire_178);
  assign mData_177 = xil_SimpleDualBram_177_doutb;
  assign xil_SimpleDualBram_178_addra = _zz_addra_178[10:0];
  assign xil_SimpleDualBram_178_addrb = _zz_addrb_178[13:0];
  assign sData_fire_179 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_178_ena = (_zz_ena_178[0] && sData_fire_179);
  assign mData_178 = xil_SimpleDualBram_178_doutb;
  assign xil_SimpleDualBram_179_addra = _zz_addra_179[10:0];
  assign xil_SimpleDualBram_179_addrb = _zz_addrb_179[13:0];
  assign sData_fire_180 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_179_ena = (_zz_ena_179[0] && sData_fire_180);
  assign mData_179 = xil_SimpleDualBram_179_doutb;
  assign xil_SimpleDualBram_180_addra = _zz_addra_180[10:0];
  assign xil_SimpleDualBram_180_addrb = _zz_addrb_180[13:0];
  assign sData_fire_181 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_180_ena = (_zz_ena_180[0] && sData_fire_181);
  assign mData_180 = xil_SimpleDualBram_180_doutb;
  assign xil_SimpleDualBram_181_addra = _zz_addra_181[10:0];
  assign xil_SimpleDualBram_181_addrb = _zz_addrb_181[13:0];
  assign sData_fire_182 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_181_ena = (_zz_ena_181[0] && sData_fire_182);
  assign mData_181 = xil_SimpleDualBram_181_doutb;
  assign xil_SimpleDualBram_182_addra = _zz_addra_182[10:0];
  assign xil_SimpleDualBram_182_addrb = _zz_addrb_182[13:0];
  assign sData_fire_183 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_182_ena = (_zz_ena_182[0] && sData_fire_183);
  assign mData_182 = xil_SimpleDualBram_182_doutb;
  assign xil_SimpleDualBram_183_addra = _zz_addra_183[10:0];
  assign xil_SimpleDualBram_183_addrb = _zz_addrb_183[13:0];
  assign sData_fire_184 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_183_ena = (_zz_ena_183[0] && sData_fire_184);
  assign mData_183 = xil_SimpleDualBram_183_doutb;
  assign xil_SimpleDualBram_184_addra = _zz_addra_184[10:0];
  assign xil_SimpleDualBram_184_addrb = _zz_addrb_184[13:0];
  assign sData_fire_185 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_184_ena = (_zz_ena_184[0] && sData_fire_185);
  assign mData_184 = xil_SimpleDualBram_184_doutb;
  assign xil_SimpleDualBram_185_addra = _zz_addra_185[10:0];
  assign xil_SimpleDualBram_185_addrb = _zz_addrb_185[13:0];
  assign sData_fire_186 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_185_ena = (_zz_ena_185[0] && sData_fire_186);
  assign mData_185 = xil_SimpleDualBram_185_doutb;
  assign xil_SimpleDualBram_186_addra = _zz_addra_186[10:0];
  assign xil_SimpleDualBram_186_addrb = _zz_addrb_186[13:0];
  assign sData_fire_187 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_186_ena = (_zz_ena_186[0] && sData_fire_187);
  assign mData_186 = xil_SimpleDualBram_186_doutb;
  assign xil_SimpleDualBram_187_addra = _zz_addra_187[10:0];
  assign xil_SimpleDualBram_187_addrb = _zz_addrb_187[13:0];
  assign sData_fire_188 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_187_ena = (_zz_ena_187[0] && sData_fire_188);
  assign mData_187 = xil_SimpleDualBram_187_doutb;
  assign xil_SimpleDualBram_188_addra = _zz_addra_188[10:0];
  assign xil_SimpleDualBram_188_addrb = _zz_addrb_188[13:0];
  assign sData_fire_189 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_188_ena = (_zz_ena_188[0] && sData_fire_189);
  assign mData_188 = xil_SimpleDualBram_188_doutb;
  assign xil_SimpleDualBram_189_addra = _zz_addra_189[10:0];
  assign xil_SimpleDualBram_189_addrb = _zz_addrb_189[13:0];
  assign sData_fire_190 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_189_ena = (_zz_ena_189[0] && sData_fire_190);
  assign mData_189 = xil_SimpleDualBram_189_doutb;
  assign xil_SimpleDualBram_190_addra = _zz_addra_190[10:0];
  assign xil_SimpleDualBram_190_addrb = _zz_addrb_190[13:0];
  assign sData_fire_191 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_190_ena = (_zz_ena_190[0] && sData_fire_191);
  assign mData_190 = xil_SimpleDualBram_190_doutb;
  assign xil_SimpleDualBram_191_addra = _zz_addra_191[10:0];
  assign xil_SimpleDualBram_191_addrb = _zz_addrb_191[13:0];
  assign sData_fire_192 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_191_ena = (_zz_ena_191[0] && sData_fire_192);
  assign mData_191 = xil_SimpleDualBram_191_doutb;
  assign xil_SimpleDualBram_192_addra = _zz_addra_192[10:0];
  assign xil_SimpleDualBram_192_addrb = _zz_addrb_192[13:0];
  assign sData_fire_193 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_192_ena = (_zz_ena_192[0] && sData_fire_193);
  assign mData_192 = xil_SimpleDualBram_192_doutb;
  assign xil_SimpleDualBram_193_addra = _zz_addra_193[10:0];
  assign xil_SimpleDualBram_193_addrb = _zz_addrb_193[13:0];
  assign sData_fire_194 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_193_ena = (_zz_ena_193[0] && sData_fire_194);
  assign mData_193 = xil_SimpleDualBram_193_doutb;
  assign xil_SimpleDualBram_194_addra = _zz_addra_194[10:0];
  assign xil_SimpleDualBram_194_addrb = _zz_addrb_194[13:0];
  assign sData_fire_195 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_194_ena = (_zz_ena_194[0] && sData_fire_195);
  assign mData_194 = xil_SimpleDualBram_194_doutb;
  assign xil_SimpleDualBram_195_addra = _zz_addra_195[10:0];
  assign xil_SimpleDualBram_195_addrb = _zz_addrb_195[13:0];
  assign sData_fire_196 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_195_ena = (_zz_ena_195[0] && sData_fire_196);
  assign mData_195 = xil_SimpleDualBram_195_doutb;
  assign xil_SimpleDualBram_196_addra = _zz_addra_196[10:0];
  assign xil_SimpleDualBram_196_addrb = _zz_addrb_196[13:0];
  assign sData_fire_197 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_196_ena = (_zz_ena_196[0] && sData_fire_197);
  assign mData_196 = xil_SimpleDualBram_196_doutb;
  assign xil_SimpleDualBram_197_addra = _zz_addra_197[10:0];
  assign xil_SimpleDualBram_197_addrb = _zz_addrb_197[13:0];
  assign sData_fire_198 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_197_ena = (_zz_ena_197[0] && sData_fire_198);
  assign mData_197 = xil_SimpleDualBram_197_doutb;
  assign xil_SimpleDualBram_198_addra = _zz_addra_198[10:0];
  assign xil_SimpleDualBram_198_addrb = _zz_addrb_198[13:0];
  assign sData_fire_199 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_198_ena = (_zz_ena_198[0] && sData_fire_199);
  assign mData_198 = xil_SimpleDualBram_198_doutb;
  assign xil_SimpleDualBram_199_addra = _zz_addra_199[10:0];
  assign xil_SimpleDualBram_199_addrb = _zz_addrb_199[13:0];
  assign sData_fire_200 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_199_ena = (_zz_ena_199[0] && sData_fire_200);
  assign mData_199 = xil_SimpleDualBram_199_doutb;
  assign xil_SimpleDualBram_200_addra = _zz_addra_200[10:0];
  assign xil_SimpleDualBram_200_addrb = _zz_addrb_200[13:0];
  assign sData_fire_201 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_200_ena = (_zz_ena_200[0] && sData_fire_201);
  assign mData_200 = xil_SimpleDualBram_200_doutb;
  assign xil_SimpleDualBram_201_addra = _zz_addra_201[10:0];
  assign xil_SimpleDualBram_201_addrb = _zz_addrb_201[13:0];
  assign sData_fire_202 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_201_ena = (_zz_ena_201[0] && sData_fire_202);
  assign mData_201 = xil_SimpleDualBram_201_doutb;
  assign xil_SimpleDualBram_202_addra = _zz_addra_202[10:0];
  assign xil_SimpleDualBram_202_addrb = _zz_addrb_202[13:0];
  assign sData_fire_203 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_202_ena = (_zz_ena_202[0] && sData_fire_203);
  assign mData_202 = xil_SimpleDualBram_202_doutb;
  assign xil_SimpleDualBram_203_addra = _zz_addra_203[10:0];
  assign xil_SimpleDualBram_203_addrb = _zz_addrb_203[13:0];
  assign sData_fire_204 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_203_ena = (_zz_ena_203[0] && sData_fire_204);
  assign mData_203 = xil_SimpleDualBram_203_doutb;
  assign xil_SimpleDualBram_204_addra = _zz_addra_204[10:0];
  assign xil_SimpleDualBram_204_addrb = _zz_addrb_204[13:0];
  assign sData_fire_205 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_204_ena = (_zz_ena_204[0] && sData_fire_205);
  assign mData_204 = xil_SimpleDualBram_204_doutb;
  assign xil_SimpleDualBram_205_addra = _zz_addra_205[10:0];
  assign xil_SimpleDualBram_205_addrb = _zz_addrb_205[13:0];
  assign sData_fire_206 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_205_ena = (_zz_ena_205[0] && sData_fire_206);
  assign mData_205 = xil_SimpleDualBram_205_doutb;
  assign xil_SimpleDualBram_206_addra = _zz_addra_206[10:0];
  assign xil_SimpleDualBram_206_addrb = _zz_addrb_206[13:0];
  assign sData_fire_207 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_206_ena = (_zz_ena_206[0] && sData_fire_207);
  assign mData_206 = xil_SimpleDualBram_206_doutb;
  assign xil_SimpleDualBram_207_addra = _zz_addra_207[10:0];
  assign xil_SimpleDualBram_207_addrb = _zz_addrb_207[13:0];
  assign sData_fire_208 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_207_ena = (_zz_ena_207[0] && sData_fire_208);
  assign mData_207 = xil_SimpleDualBram_207_doutb;
  assign xil_SimpleDualBram_208_addra = _zz_addra_208[10:0];
  assign xil_SimpleDualBram_208_addrb = _zz_addrb_208[13:0];
  assign sData_fire_209 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_208_ena = (_zz_ena_208[0] && sData_fire_209);
  assign mData_208 = xil_SimpleDualBram_208_doutb;
  assign xil_SimpleDualBram_209_addra = _zz_addra_209[10:0];
  assign xil_SimpleDualBram_209_addrb = _zz_addrb_209[13:0];
  assign sData_fire_210 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_209_ena = (_zz_ena_209[0] && sData_fire_210);
  assign mData_209 = xil_SimpleDualBram_209_doutb;
  assign xil_SimpleDualBram_210_addra = _zz_addra_210[10:0];
  assign xil_SimpleDualBram_210_addrb = _zz_addrb_210[13:0];
  assign sData_fire_211 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_210_ena = (_zz_ena_210[0] && sData_fire_211);
  assign mData_210 = xil_SimpleDualBram_210_doutb;
  assign xil_SimpleDualBram_211_addra = _zz_addra_211[10:0];
  assign xil_SimpleDualBram_211_addrb = _zz_addrb_211[13:0];
  assign sData_fire_212 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_211_ena = (_zz_ena_211[0] && sData_fire_212);
  assign mData_211 = xil_SimpleDualBram_211_doutb;
  assign xil_SimpleDualBram_212_addra = _zz_addra_212[10:0];
  assign xil_SimpleDualBram_212_addrb = _zz_addrb_212[13:0];
  assign sData_fire_213 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_212_ena = (_zz_ena_212[0] && sData_fire_213);
  assign mData_212 = xil_SimpleDualBram_212_doutb;
  assign xil_SimpleDualBram_213_addra = _zz_addra_213[10:0];
  assign xil_SimpleDualBram_213_addrb = _zz_addrb_213[13:0];
  assign sData_fire_214 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_213_ena = (_zz_ena_213[0] && sData_fire_214);
  assign mData_213 = xil_SimpleDualBram_213_doutb;
  assign xil_SimpleDualBram_214_addra = _zz_addra_214[10:0];
  assign xil_SimpleDualBram_214_addrb = _zz_addrb_214[13:0];
  assign sData_fire_215 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_214_ena = (_zz_ena_214[0] && sData_fire_215);
  assign mData_214 = xil_SimpleDualBram_214_doutb;
  assign xil_SimpleDualBram_215_addra = _zz_addra_215[10:0];
  assign xil_SimpleDualBram_215_addrb = _zz_addrb_215[13:0];
  assign sData_fire_216 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_215_ena = (_zz_ena_215[0] && sData_fire_216);
  assign mData_215 = xil_SimpleDualBram_215_doutb;
  assign xil_SimpleDualBram_216_addra = _zz_addra_216[10:0];
  assign xil_SimpleDualBram_216_addrb = _zz_addrb_216[13:0];
  assign sData_fire_217 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_216_ena = (_zz_ena_216[0] && sData_fire_217);
  assign mData_216 = xil_SimpleDualBram_216_doutb;
  assign xil_SimpleDualBram_217_addra = _zz_addra_217[10:0];
  assign xil_SimpleDualBram_217_addrb = _zz_addrb_217[13:0];
  assign sData_fire_218 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_217_ena = (_zz_ena_217[0] && sData_fire_218);
  assign mData_217 = xil_SimpleDualBram_217_doutb;
  assign xil_SimpleDualBram_218_addra = _zz_addra_218[10:0];
  assign xil_SimpleDualBram_218_addrb = _zz_addrb_218[13:0];
  assign sData_fire_219 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_218_ena = (_zz_ena_218[0] && sData_fire_219);
  assign mData_218 = xil_SimpleDualBram_218_doutb;
  assign xil_SimpleDualBram_219_addra = _zz_addra_219[10:0];
  assign xil_SimpleDualBram_219_addrb = _zz_addrb_219[13:0];
  assign sData_fire_220 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_219_ena = (_zz_ena_219[0] && sData_fire_220);
  assign mData_219 = xil_SimpleDualBram_219_doutb;
  assign xil_SimpleDualBram_220_addra = _zz_addra_220[10:0];
  assign xil_SimpleDualBram_220_addrb = _zz_addrb_220[13:0];
  assign sData_fire_221 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_220_ena = (_zz_ena_220[0] && sData_fire_221);
  assign mData_220 = xil_SimpleDualBram_220_doutb;
  assign xil_SimpleDualBram_221_addra = _zz_addra_221[10:0];
  assign xil_SimpleDualBram_221_addrb = _zz_addrb_221[13:0];
  assign sData_fire_222 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_221_ena = (_zz_ena_221[0] && sData_fire_222);
  assign mData_221 = xil_SimpleDualBram_221_doutb;
  assign xil_SimpleDualBram_222_addra = _zz_addra_222[10:0];
  assign xil_SimpleDualBram_222_addrb = _zz_addrb_222[13:0];
  assign sData_fire_223 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_222_ena = (_zz_ena_222[0] && sData_fire_223);
  assign mData_222 = xil_SimpleDualBram_222_doutb;
  assign xil_SimpleDualBram_223_addra = _zz_addra_223[10:0];
  assign xil_SimpleDualBram_223_addrb = _zz_addrb_223[13:0];
  assign sData_fire_224 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_223_ena = (_zz_ena_223[0] && sData_fire_224);
  assign mData_223 = xil_SimpleDualBram_223_doutb;
  assign xil_SimpleDualBram_224_addra = _zz_addra_224[10:0];
  assign xil_SimpleDualBram_224_addrb = _zz_addrb_224[13:0];
  assign sData_fire_225 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_224_ena = (_zz_ena_224[0] && sData_fire_225);
  assign mData_224 = xil_SimpleDualBram_224_doutb;
  assign xil_SimpleDualBram_225_addra = _zz_addra_225[10:0];
  assign xil_SimpleDualBram_225_addrb = _zz_addrb_225[13:0];
  assign sData_fire_226 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_225_ena = (_zz_ena_225[0] && sData_fire_226);
  assign mData_225 = xil_SimpleDualBram_225_doutb;
  assign xil_SimpleDualBram_226_addra = _zz_addra_226[10:0];
  assign xil_SimpleDualBram_226_addrb = _zz_addrb_226[13:0];
  assign sData_fire_227 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_226_ena = (_zz_ena_226[0] && sData_fire_227);
  assign mData_226 = xil_SimpleDualBram_226_doutb;
  assign xil_SimpleDualBram_227_addra = _zz_addra_227[10:0];
  assign xil_SimpleDualBram_227_addrb = _zz_addrb_227[13:0];
  assign sData_fire_228 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_227_ena = (_zz_ena_227[0] && sData_fire_228);
  assign mData_227 = xil_SimpleDualBram_227_doutb;
  assign xil_SimpleDualBram_228_addra = _zz_addra_228[10:0];
  assign xil_SimpleDualBram_228_addrb = _zz_addrb_228[13:0];
  assign sData_fire_229 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_228_ena = (_zz_ena_228[0] && sData_fire_229);
  assign mData_228 = xil_SimpleDualBram_228_doutb;
  assign xil_SimpleDualBram_229_addra = _zz_addra_229[10:0];
  assign xil_SimpleDualBram_229_addrb = _zz_addrb_229[13:0];
  assign sData_fire_230 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_229_ena = (_zz_ena_229[0] && sData_fire_230);
  assign mData_229 = xil_SimpleDualBram_229_doutb;
  assign xil_SimpleDualBram_230_addra = _zz_addra_230[10:0];
  assign xil_SimpleDualBram_230_addrb = _zz_addrb_230[13:0];
  assign sData_fire_231 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_230_ena = (_zz_ena_230[0] && sData_fire_231);
  assign mData_230 = xil_SimpleDualBram_230_doutb;
  assign xil_SimpleDualBram_231_addra = _zz_addra_231[10:0];
  assign xil_SimpleDualBram_231_addrb = _zz_addrb_231[13:0];
  assign sData_fire_232 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_231_ena = (_zz_ena_231[0] && sData_fire_232);
  assign mData_231 = xil_SimpleDualBram_231_doutb;
  assign xil_SimpleDualBram_232_addra = _zz_addra_232[10:0];
  assign xil_SimpleDualBram_232_addrb = _zz_addrb_232[13:0];
  assign sData_fire_233 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_232_ena = (_zz_ena_232[0] && sData_fire_233);
  assign mData_232 = xil_SimpleDualBram_232_doutb;
  assign xil_SimpleDualBram_233_addra = _zz_addra_233[10:0];
  assign xil_SimpleDualBram_233_addrb = _zz_addrb_233[13:0];
  assign sData_fire_234 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_233_ena = (_zz_ena_233[0] && sData_fire_234);
  assign mData_233 = xil_SimpleDualBram_233_doutb;
  assign xil_SimpleDualBram_234_addra = _zz_addra_234[10:0];
  assign xil_SimpleDualBram_234_addrb = _zz_addrb_234[13:0];
  assign sData_fire_235 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_234_ena = (_zz_ena_234[0] && sData_fire_235);
  assign mData_234 = xil_SimpleDualBram_234_doutb;
  assign xil_SimpleDualBram_235_addra = _zz_addra_235[10:0];
  assign xil_SimpleDualBram_235_addrb = _zz_addrb_235[13:0];
  assign sData_fire_236 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_235_ena = (_zz_ena_235[0] && sData_fire_236);
  assign mData_235 = xil_SimpleDualBram_235_doutb;
  assign xil_SimpleDualBram_236_addra = _zz_addra_236[10:0];
  assign xil_SimpleDualBram_236_addrb = _zz_addrb_236[13:0];
  assign sData_fire_237 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_236_ena = (_zz_ena_236[0] && sData_fire_237);
  assign mData_236 = xil_SimpleDualBram_236_doutb;
  assign xil_SimpleDualBram_237_addra = _zz_addra_237[10:0];
  assign xil_SimpleDualBram_237_addrb = _zz_addrb_237[13:0];
  assign sData_fire_238 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_237_ena = (_zz_ena_237[0] && sData_fire_238);
  assign mData_237 = xil_SimpleDualBram_237_doutb;
  assign xil_SimpleDualBram_238_addra = _zz_addra_238[10:0];
  assign xil_SimpleDualBram_238_addrb = _zz_addrb_238[13:0];
  assign sData_fire_239 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_238_ena = (_zz_ena_238[0] && sData_fire_239);
  assign mData_238 = xil_SimpleDualBram_238_doutb;
  assign xil_SimpleDualBram_239_addra = _zz_addra_239[10:0];
  assign xil_SimpleDualBram_239_addrb = _zz_addrb_239[13:0];
  assign sData_fire_240 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_239_ena = (_zz_ena_239[0] && sData_fire_240);
  assign mData_239 = xil_SimpleDualBram_239_doutb;
  assign xil_SimpleDualBram_240_addra = _zz_addra_240[10:0];
  assign xil_SimpleDualBram_240_addrb = _zz_addrb_240[13:0];
  assign sData_fire_241 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_240_ena = (_zz_ena_240[0] && sData_fire_241);
  assign mData_240 = xil_SimpleDualBram_240_doutb;
  assign xil_SimpleDualBram_241_addra = _zz_addra_241[10:0];
  assign xil_SimpleDualBram_241_addrb = _zz_addrb_241[13:0];
  assign sData_fire_242 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_241_ena = (_zz_ena_241[0] && sData_fire_242);
  assign mData_241 = xil_SimpleDualBram_241_doutb;
  assign xil_SimpleDualBram_242_addra = _zz_addra_242[10:0];
  assign xil_SimpleDualBram_242_addrb = _zz_addrb_242[13:0];
  assign sData_fire_243 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_242_ena = (_zz_ena_242[0] && sData_fire_243);
  assign mData_242 = xil_SimpleDualBram_242_doutb;
  assign xil_SimpleDualBram_243_addra = _zz_addra_243[10:0];
  assign xil_SimpleDualBram_243_addrb = _zz_addrb_243[13:0];
  assign sData_fire_244 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_243_ena = (_zz_ena_243[0] && sData_fire_244);
  assign mData_243 = xil_SimpleDualBram_243_doutb;
  assign xil_SimpleDualBram_244_addra = _zz_addra_244[10:0];
  assign xil_SimpleDualBram_244_addrb = _zz_addrb_244[13:0];
  assign sData_fire_245 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_244_ena = (_zz_ena_244[0] && sData_fire_245);
  assign mData_244 = xil_SimpleDualBram_244_doutb;
  assign xil_SimpleDualBram_245_addra = _zz_addra_245[10:0];
  assign xil_SimpleDualBram_245_addrb = _zz_addrb_245[13:0];
  assign sData_fire_246 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_245_ena = (_zz_ena_245[0] && sData_fire_246);
  assign mData_245 = xil_SimpleDualBram_245_doutb;
  assign xil_SimpleDualBram_246_addra = _zz_addra_246[10:0];
  assign xil_SimpleDualBram_246_addrb = _zz_addrb_246[13:0];
  assign sData_fire_247 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_246_ena = (_zz_ena_246[0] && sData_fire_247);
  assign mData_246 = xil_SimpleDualBram_246_doutb;
  assign xil_SimpleDualBram_247_addra = _zz_addra_247[10:0];
  assign xil_SimpleDualBram_247_addrb = _zz_addrb_247[13:0];
  assign sData_fire_248 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_247_ena = (_zz_ena_247[0] && sData_fire_248);
  assign mData_247 = xil_SimpleDualBram_247_doutb;
  assign xil_SimpleDualBram_248_addra = _zz_addra_248[10:0];
  assign xil_SimpleDualBram_248_addrb = _zz_addrb_248[13:0];
  assign sData_fire_249 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_248_ena = (_zz_ena_248[0] && sData_fire_249);
  assign mData_248 = xil_SimpleDualBram_248_doutb;
  assign xil_SimpleDualBram_249_addra = _zz_addra_249[10:0];
  assign xil_SimpleDualBram_249_addrb = _zz_addrb_249[13:0];
  assign sData_fire_250 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_249_ena = (_zz_ena_249[0] && sData_fire_250);
  assign mData_249 = xil_SimpleDualBram_249_doutb;
  assign xil_SimpleDualBram_250_addra = _zz_addra_250[10:0];
  assign xil_SimpleDualBram_250_addrb = _zz_addrb_250[13:0];
  assign sData_fire_251 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_250_ena = (_zz_ena_250[0] && sData_fire_251);
  assign mData_250 = xil_SimpleDualBram_250_doutb;
  assign xil_SimpleDualBram_251_addra = _zz_addra_251[10:0];
  assign xil_SimpleDualBram_251_addrb = _zz_addrb_251[13:0];
  assign sData_fire_252 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_251_ena = (_zz_ena_251[0] && sData_fire_252);
  assign mData_251 = xil_SimpleDualBram_251_doutb;
  assign xil_SimpleDualBram_252_addra = _zz_addra_252[10:0];
  assign xil_SimpleDualBram_252_addrb = _zz_addrb_252[13:0];
  assign sData_fire_253 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_252_ena = (_zz_ena_252[0] && sData_fire_253);
  assign mData_252 = xil_SimpleDualBram_252_doutb;
  assign xil_SimpleDualBram_253_addra = _zz_addra_253[10:0];
  assign xil_SimpleDualBram_253_addrb = _zz_addrb_253[13:0];
  assign sData_fire_254 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_253_ena = (_zz_ena_253[0] && sData_fire_254);
  assign mData_253 = xil_SimpleDualBram_253_doutb;
  assign xil_SimpleDualBram_254_addra = _zz_addra_254[10:0];
  assign xil_SimpleDualBram_254_addrb = _zz_addrb_254[13:0];
  assign sData_fire_255 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_254_ena = (_zz_ena_254[0] && sData_fire_255);
  assign mData_254 = xil_SimpleDualBram_254_doutb;
  assign xil_SimpleDualBram_255_addra = _zz_addra_255[10:0];
  assign xil_SimpleDualBram_255_addrb = _zz_addrb_255[13:0];
  assign sData_fire_256 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_255_ena = (_zz_ena_255[0] && sData_fire_256);
  assign mData_255 = xil_SimpleDualBram_255_doutb;
  assign xil_SimpleDualBram_256_addra = _zz_addra_256[10:0];
  assign xil_SimpleDualBram_256_addrb = _zz_addrb_256[13:0];
  assign sData_fire_257 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_256_ena = (_zz_ena_256[0] && sData_fire_257);
  assign mData_256 = xil_SimpleDualBram_256_doutb;
  assign xil_SimpleDualBram_257_addra = _zz_addra_257[10:0];
  assign xil_SimpleDualBram_257_addrb = _zz_addrb_257[13:0];
  assign sData_fire_258 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_257_ena = (_zz_ena_257[0] && sData_fire_258);
  assign mData_257 = xil_SimpleDualBram_257_doutb;
  assign xil_SimpleDualBram_258_addra = _zz_addra_258[10:0];
  assign xil_SimpleDualBram_258_addrb = _zz_addrb_258[13:0];
  assign sData_fire_259 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_258_ena = (_zz_ena_258[0] && sData_fire_259);
  assign mData_258 = xil_SimpleDualBram_258_doutb;
  assign xil_SimpleDualBram_259_addra = _zz_addra_259[10:0];
  assign xil_SimpleDualBram_259_addrb = _zz_addrb_259[13:0];
  assign sData_fire_260 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_259_ena = (_zz_ena_259[0] && sData_fire_260);
  assign mData_259 = xil_SimpleDualBram_259_doutb;
  assign xil_SimpleDualBram_260_addra = _zz_addra_260[10:0];
  assign xil_SimpleDualBram_260_addrb = _zz_addrb_260[13:0];
  assign sData_fire_261 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_260_ena = (_zz_ena_260[0] && sData_fire_261);
  assign mData_260 = xil_SimpleDualBram_260_doutb;
  assign xil_SimpleDualBram_261_addra = _zz_addra_261[10:0];
  assign xil_SimpleDualBram_261_addrb = _zz_addrb_261[13:0];
  assign sData_fire_262 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_261_ena = (_zz_ena_261[0] && sData_fire_262);
  assign mData_261 = xil_SimpleDualBram_261_doutb;
  assign xil_SimpleDualBram_262_addra = _zz_addra_262[10:0];
  assign xil_SimpleDualBram_262_addrb = _zz_addrb_262[13:0];
  assign sData_fire_263 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_262_ena = (_zz_ena_262[0] && sData_fire_263);
  assign mData_262 = xil_SimpleDualBram_262_doutb;
  assign xil_SimpleDualBram_263_addra = _zz_addra_263[10:0];
  assign xil_SimpleDualBram_263_addrb = _zz_addrb_263[13:0];
  assign sData_fire_264 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_263_ena = (_zz_ena_263[0] && sData_fire_264);
  assign mData_263 = xil_SimpleDualBram_263_doutb;
  assign xil_SimpleDualBram_264_addra = _zz_addra_264[10:0];
  assign xil_SimpleDualBram_264_addrb = _zz_addrb_264[13:0];
  assign sData_fire_265 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_264_ena = (_zz_ena_264[0] && sData_fire_265);
  assign mData_264 = xil_SimpleDualBram_264_doutb;
  assign xil_SimpleDualBram_265_addra = _zz_addra_265[10:0];
  assign xil_SimpleDualBram_265_addrb = _zz_addrb_265[13:0];
  assign sData_fire_266 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_265_ena = (_zz_ena_265[0] && sData_fire_266);
  assign mData_265 = xil_SimpleDualBram_265_doutb;
  assign xil_SimpleDualBram_266_addra = _zz_addra_266[10:0];
  assign xil_SimpleDualBram_266_addrb = _zz_addrb_266[13:0];
  assign sData_fire_267 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_266_ena = (_zz_ena_266[0] && sData_fire_267);
  assign mData_266 = xil_SimpleDualBram_266_doutb;
  assign xil_SimpleDualBram_267_addra = _zz_addra_267[10:0];
  assign xil_SimpleDualBram_267_addrb = _zz_addrb_267[13:0];
  assign sData_fire_268 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_267_ena = (_zz_ena_267[0] && sData_fire_268);
  assign mData_267 = xil_SimpleDualBram_267_doutb;
  assign xil_SimpleDualBram_268_addra = _zz_addra_268[10:0];
  assign xil_SimpleDualBram_268_addrb = _zz_addrb_268[13:0];
  assign sData_fire_269 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_268_ena = (_zz_ena_268[0] && sData_fire_269);
  assign mData_268 = xil_SimpleDualBram_268_doutb;
  assign xil_SimpleDualBram_269_addra = _zz_addra_269[10:0];
  assign xil_SimpleDualBram_269_addrb = _zz_addrb_269[13:0];
  assign sData_fire_270 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_269_ena = (_zz_ena_269[0] && sData_fire_270);
  assign mData_269 = xil_SimpleDualBram_269_doutb;
  assign xil_SimpleDualBram_270_addra = _zz_addra_270[10:0];
  assign xil_SimpleDualBram_270_addrb = _zz_addrb_270[13:0];
  assign sData_fire_271 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_270_ena = (_zz_ena_270[0] && sData_fire_271);
  assign mData_270 = xil_SimpleDualBram_270_doutb;
  assign xil_SimpleDualBram_271_addra = _zz_addra_271[10:0];
  assign xil_SimpleDualBram_271_addrb = _zz_addrb_271[13:0];
  assign sData_fire_272 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_271_ena = (_zz_ena_271[0] && sData_fire_272);
  assign mData_271 = xil_SimpleDualBram_271_doutb;
  assign xil_SimpleDualBram_272_addra = _zz_addra_272[10:0];
  assign xil_SimpleDualBram_272_addrb = _zz_addrb_272[13:0];
  assign sData_fire_273 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_272_ena = (_zz_ena_272[0] && sData_fire_273);
  assign mData_272 = xil_SimpleDualBram_272_doutb;
  assign xil_SimpleDualBram_273_addra = _zz_addra_273[10:0];
  assign xil_SimpleDualBram_273_addrb = _zz_addrb_273[13:0];
  assign sData_fire_274 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_273_ena = (_zz_ena_273[0] && sData_fire_274);
  assign mData_273 = xil_SimpleDualBram_273_doutb;
  assign xil_SimpleDualBram_274_addra = _zz_addra_274[10:0];
  assign xil_SimpleDualBram_274_addrb = _zz_addrb_274[13:0];
  assign sData_fire_275 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_274_ena = (_zz_ena_274[0] && sData_fire_275);
  assign mData_274 = xil_SimpleDualBram_274_doutb;
  assign xil_SimpleDualBram_275_addra = _zz_addra_275[10:0];
  assign xil_SimpleDualBram_275_addrb = _zz_addrb_275[13:0];
  assign sData_fire_276 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_275_ena = (_zz_ena_275[0] && sData_fire_276);
  assign mData_275 = xil_SimpleDualBram_275_doutb;
  assign xil_SimpleDualBram_276_addra = _zz_addra_276[10:0];
  assign xil_SimpleDualBram_276_addrb = _zz_addrb_276[13:0];
  assign sData_fire_277 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_276_ena = (_zz_ena_276[0] && sData_fire_277);
  assign mData_276 = xil_SimpleDualBram_276_doutb;
  assign xil_SimpleDualBram_277_addra = _zz_addra_277[10:0];
  assign xil_SimpleDualBram_277_addrb = _zz_addrb_277[13:0];
  assign sData_fire_278 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_277_ena = (_zz_ena_277[0] && sData_fire_278);
  assign mData_277 = xil_SimpleDualBram_277_doutb;
  assign xil_SimpleDualBram_278_addra = _zz_addra_278[10:0];
  assign xil_SimpleDualBram_278_addrb = _zz_addrb_278[13:0];
  assign sData_fire_279 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_278_ena = (_zz_ena_278[0] && sData_fire_279);
  assign mData_278 = xil_SimpleDualBram_278_doutb;
  assign xil_SimpleDualBram_279_addra = _zz_addra_279[10:0];
  assign xil_SimpleDualBram_279_addrb = _zz_addrb_279[13:0];
  assign sData_fire_280 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_279_ena = (_zz_ena_279[0] && sData_fire_280);
  assign mData_279 = xil_SimpleDualBram_279_doutb;
  assign xil_SimpleDualBram_280_addra = _zz_addra_280[10:0];
  assign xil_SimpleDualBram_280_addrb = _zz_addrb_280[13:0];
  assign sData_fire_281 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_280_ena = (_zz_ena_280[0] && sData_fire_281);
  assign mData_280 = xil_SimpleDualBram_280_doutb;
  assign xil_SimpleDualBram_281_addra = _zz_addra_281[10:0];
  assign xil_SimpleDualBram_281_addrb = _zz_addrb_281[13:0];
  assign sData_fire_282 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_281_ena = (_zz_ena_281[0] && sData_fire_282);
  assign mData_281 = xil_SimpleDualBram_281_doutb;
  assign xil_SimpleDualBram_282_addra = _zz_addra_282[10:0];
  assign xil_SimpleDualBram_282_addrb = _zz_addrb_282[13:0];
  assign sData_fire_283 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_282_ena = (_zz_ena_282[0] && sData_fire_283);
  assign mData_282 = xil_SimpleDualBram_282_doutb;
  assign xil_SimpleDualBram_283_addra = _zz_addra_283[10:0];
  assign xil_SimpleDualBram_283_addrb = _zz_addrb_283[13:0];
  assign sData_fire_284 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_283_ena = (_zz_ena_283[0] && sData_fire_284);
  assign mData_283 = xil_SimpleDualBram_283_doutb;
  assign xil_SimpleDualBram_284_addra = _zz_addra_284[10:0];
  assign xil_SimpleDualBram_284_addrb = _zz_addrb_284[13:0];
  assign sData_fire_285 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_284_ena = (_zz_ena_284[0] && sData_fire_285);
  assign mData_284 = xil_SimpleDualBram_284_doutb;
  assign xil_SimpleDualBram_285_addra = _zz_addra_285[10:0];
  assign xil_SimpleDualBram_285_addrb = _zz_addrb_285[13:0];
  assign sData_fire_286 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_285_ena = (_zz_ena_285[0] && sData_fire_286);
  assign mData_285 = xil_SimpleDualBram_285_doutb;
  assign xil_SimpleDualBram_286_addra = _zz_addra_286[10:0];
  assign xil_SimpleDualBram_286_addrb = _zz_addrb_286[13:0];
  assign sData_fire_287 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_286_ena = (_zz_ena_286[0] && sData_fire_287);
  assign mData_286 = xil_SimpleDualBram_286_doutb;
  assign xil_SimpleDualBram_287_addra = _zz_addra_287[10:0];
  assign xil_SimpleDualBram_287_addrb = _zz_addrb_287[13:0];
  assign sData_fire_288 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_287_ena = (_zz_ena_287[0] && sData_fire_288);
  assign mData_287 = xil_SimpleDualBram_287_doutb;
  assign xil_SimpleDualBram_288_addra = _zz_addra_288[10:0];
  assign xil_SimpleDualBram_288_addrb = _zz_addrb_288[13:0];
  assign sData_fire_289 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_288_ena = (_zz_ena_288[0] && sData_fire_289);
  assign mData_288 = xil_SimpleDualBram_288_doutb;
  assign xil_SimpleDualBram_289_addra = _zz_addra_289[10:0];
  assign xil_SimpleDualBram_289_addrb = _zz_addrb_289[13:0];
  assign sData_fire_290 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_289_ena = (_zz_ena_289[0] && sData_fire_290);
  assign mData_289 = xil_SimpleDualBram_289_doutb;
  assign xil_SimpleDualBram_290_addra = _zz_addra_290[10:0];
  assign xil_SimpleDualBram_290_addrb = _zz_addrb_290[13:0];
  assign sData_fire_291 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_290_ena = (_zz_ena_290[0] && sData_fire_291);
  assign mData_290 = xil_SimpleDualBram_290_doutb;
  assign xil_SimpleDualBram_291_addra = _zz_addra_291[10:0];
  assign xil_SimpleDualBram_291_addrb = _zz_addrb_291[13:0];
  assign sData_fire_292 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_291_ena = (_zz_ena_291[0] && sData_fire_292);
  assign mData_291 = xil_SimpleDualBram_291_doutb;
  assign xil_SimpleDualBram_292_addra = _zz_addra_292[10:0];
  assign xil_SimpleDualBram_292_addrb = _zz_addrb_292[13:0];
  assign sData_fire_293 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_292_ena = (_zz_ena_292[0] && sData_fire_293);
  assign mData_292 = xil_SimpleDualBram_292_doutb;
  assign xil_SimpleDualBram_293_addra = _zz_addra_293[10:0];
  assign xil_SimpleDualBram_293_addrb = _zz_addrb_293[13:0];
  assign sData_fire_294 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_293_ena = (_zz_ena_293[0] && sData_fire_294);
  assign mData_293 = xil_SimpleDualBram_293_doutb;
  assign xil_SimpleDualBram_294_addra = _zz_addra_294[10:0];
  assign xil_SimpleDualBram_294_addrb = _zz_addrb_294[13:0];
  assign sData_fire_295 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_294_ena = (_zz_ena_294[0] && sData_fire_295);
  assign mData_294 = xil_SimpleDualBram_294_doutb;
  assign xil_SimpleDualBram_295_addra = _zz_addra_295[10:0];
  assign xil_SimpleDualBram_295_addrb = _zz_addrb_295[13:0];
  assign sData_fire_296 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_295_ena = (_zz_ena_295[0] && sData_fire_296);
  assign mData_295 = xil_SimpleDualBram_295_doutb;
  assign xil_SimpleDualBram_296_addra = _zz_addra_296[10:0];
  assign xil_SimpleDualBram_296_addrb = _zz_addrb_296[13:0];
  assign sData_fire_297 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_296_ena = (_zz_ena_296[0] && sData_fire_297);
  assign mData_296 = xil_SimpleDualBram_296_doutb;
  assign xil_SimpleDualBram_297_addra = _zz_addra_297[10:0];
  assign xil_SimpleDualBram_297_addrb = _zz_addrb_297[13:0];
  assign sData_fire_298 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_297_ena = (_zz_ena_297[0] && sData_fire_298);
  assign mData_297 = xil_SimpleDualBram_297_doutb;
  assign xil_SimpleDualBram_298_addra = _zz_addra_298[10:0];
  assign xil_SimpleDualBram_298_addrb = _zz_addrb_298[13:0];
  assign sData_fire_299 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_298_ena = (_zz_ena_298[0] && sData_fire_299);
  assign mData_298 = xil_SimpleDualBram_298_doutb;
  assign xil_SimpleDualBram_299_addra = _zz_addra_299[10:0];
  assign xil_SimpleDualBram_299_addrb = _zz_addrb_299[13:0];
  assign sData_fire_300 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_299_ena = (_zz_ena_299[0] && sData_fire_300);
  assign mData_299 = xil_SimpleDualBram_299_doutb;
  assign xil_SimpleDualBram_300_addra = _zz_addra_300[10:0];
  assign xil_SimpleDualBram_300_addrb = _zz_addrb_300[13:0];
  assign sData_fire_301 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_300_ena = (_zz_ena_300[0] && sData_fire_301);
  assign mData_300 = xil_SimpleDualBram_300_doutb;
  assign xil_SimpleDualBram_301_addra = _zz_addra_301[10:0];
  assign xil_SimpleDualBram_301_addrb = _zz_addrb_301[13:0];
  assign sData_fire_302 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_301_ena = (_zz_ena_301[0] && sData_fire_302);
  assign mData_301 = xil_SimpleDualBram_301_doutb;
  assign xil_SimpleDualBram_302_addra = _zz_addra_302[10:0];
  assign xil_SimpleDualBram_302_addrb = _zz_addrb_302[13:0];
  assign sData_fire_303 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_302_ena = (_zz_ena_302[0] && sData_fire_303);
  assign mData_302 = xil_SimpleDualBram_302_doutb;
  assign xil_SimpleDualBram_303_addra = _zz_addra_303[10:0];
  assign xil_SimpleDualBram_303_addrb = _zz_addrb_303[13:0];
  assign sData_fire_304 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_303_ena = (_zz_ena_303[0] && sData_fire_304);
  assign mData_303 = xil_SimpleDualBram_303_doutb;
  assign xil_SimpleDualBram_304_addra = _zz_addra_304[10:0];
  assign xil_SimpleDualBram_304_addrb = _zz_addrb_304[13:0];
  assign sData_fire_305 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_304_ena = (_zz_ena_304[0] && sData_fire_305);
  assign mData_304 = xil_SimpleDualBram_304_doutb;
  assign xil_SimpleDualBram_305_addra = _zz_addra_305[10:0];
  assign xil_SimpleDualBram_305_addrb = _zz_addrb_305[13:0];
  assign sData_fire_306 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_305_ena = (_zz_ena_305[0] && sData_fire_306);
  assign mData_305 = xil_SimpleDualBram_305_doutb;
  assign xil_SimpleDualBram_306_addra = _zz_addra_306[10:0];
  assign xil_SimpleDualBram_306_addrb = _zz_addrb_306[13:0];
  assign sData_fire_307 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_306_ena = (_zz_ena_306[0] && sData_fire_307);
  assign mData_306 = xil_SimpleDualBram_306_doutb;
  assign xil_SimpleDualBram_307_addra = _zz_addra_307[10:0];
  assign xil_SimpleDualBram_307_addrb = _zz_addrb_307[13:0];
  assign sData_fire_308 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_307_ena = (_zz_ena_307[0] && sData_fire_308);
  assign mData_307 = xil_SimpleDualBram_307_doutb;
  assign xil_SimpleDualBram_308_addra = _zz_addra_308[10:0];
  assign xil_SimpleDualBram_308_addrb = _zz_addrb_308[13:0];
  assign sData_fire_309 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_308_ena = (_zz_ena_308[0] && sData_fire_309);
  assign mData_308 = xil_SimpleDualBram_308_doutb;
  assign xil_SimpleDualBram_309_addra = _zz_addra_309[10:0];
  assign xil_SimpleDualBram_309_addrb = _zz_addrb_309[13:0];
  assign sData_fire_310 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_309_ena = (_zz_ena_309[0] && sData_fire_310);
  assign mData_309 = xil_SimpleDualBram_309_doutb;
  assign xil_SimpleDualBram_310_addra = _zz_addra_310[10:0];
  assign xil_SimpleDualBram_310_addrb = _zz_addrb_310[13:0];
  assign sData_fire_311 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_310_ena = (_zz_ena_310[0] && sData_fire_311);
  assign mData_310 = xil_SimpleDualBram_310_doutb;
  assign xil_SimpleDualBram_311_addra = _zz_addra_311[10:0];
  assign xil_SimpleDualBram_311_addrb = _zz_addrb_311[13:0];
  assign sData_fire_312 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_311_ena = (_zz_ena_311[0] && sData_fire_312);
  assign mData_311 = xil_SimpleDualBram_311_doutb;
  assign xil_SimpleDualBram_312_addra = _zz_addra_312[10:0];
  assign xil_SimpleDualBram_312_addrb = _zz_addrb_312[13:0];
  assign sData_fire_313 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_312_ena = (_zz_ena_312[0] && sData_fire_313);
  assign mData_312 = xil_SimpleDualBram_312_doutb;
  assign xil_SimpleDualBram_313_addra = _zz_addra_313[10:0];
  assign xil_SimpleDualBram_313_addrb = _zz_addrb_313[13:0];
  assign sData_fire_314 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_313_ena = (_zz_ena_313[0] && sData_fire_314);
  assign mData_313 = xil_SimpleDualBram_313_doutb;
  assign xil_SimpleDualBram_314_addra = _zz_addra_314[10:0];
  assign xil_SimpleDualBram_314_addrb = _zz_addrb_314[13:0];
  assign sData_fire_315 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_314_ena = (_zz_ena_314[0] && sData_fire_315);
  assign mData_314 = xil_SimpleDualBram_314_doutb;
  assign xil_SimpleDualBram_315_addra = _zz_addra_315[10:0];
  assign xil_SimpleDualBram_315_addrb = _zz_addrb_315[13:0];
  assign sData_fire_316 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_315_ena = (_zz_ena_315[0] && sData_fire_316);
  assign mData_315 = xil_SimpleDualBram_315_doutb;
  assign xil_SimpleDualBram_316_addra = _zz_addra_316[10:0];
  assign xil_SimpleDualBram_316_addrb = _zz_addrb_316[13:0];
  assign sData_fire_317 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_316_ena = (_zz_ena_316[0] && sData_fire_317);
  assign mData_316 = xil_SimpleDualBram_316_doutb;
  assign xil_SimpleDualBram_317_addra = _zz_addra_317[10:0];
  assign xil_SimpleDualBram_317_addrb = _zz_addrb_317[13:0];
  assign sData_fire_318 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_317_ena = (_zz_ena_317[0] && sData_fire_318);
  assign mData_317 = xil_SimpleDualBram_317_doutb;
  assign xil_SimpleDualBram_318_addra = _zz_addra_318[10:0];
  assign xil_SimpleDualBram_318_addrb = _zz_addrb_318[13:0];
  assign sData_fire_319 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_318_ena = (_zz_ena_318[0] && sData_fire_319);
  assign mData_318 = xil_SimpleDualBram_318_doutb;
  assign xil_SimpleDualBram_319_addra = _zz_addra_319[10:0];
  assign xil_SimpleDualBram_319_addrb = _zz_addrb_319[13:0];
  assign sData_fire_320 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_319_ena = (_zz_ena_319[0] && sData_fire_320);
  assign mData_319 = xil_SimpleDualBram_319_doutb;
  assign xil_SimpleDualBram_320_addra = _zz_addra_320[10:0];
  assign xil_SimpleDualBram_320_addrb = _zz_addrb_320[13:0];
  assign sData_fire_321 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_320_ena = (_zz_ena_320[0] && sData_fire_321);
  assign mData_320 = xil_SimpleDualBram_320_doutb;
  assign xil_SimpleDualBram_321_addra = _zz_addra_321[10:0];
  assign xil_SimpleDualBram_321_addrb = _zz_addrb_321[13:0];
  assign sData_fire_322 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_321_ena = (_zz_ena_321[0] && sData_fire_322);
  assign mData_321 = xil_SimpleDualBram_321_doutb;
  assign xil_SimpleDualBram_322_addra = _zz_addra_322[10:0];
  assign xil_SimpleDualBram_322_addrb = _zz_addrb_322[13:0];
  assign sData_fire_323 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_322_ena = (_zz_ena_322[0] && sData_fire_323);
  assign mData_322 = xil_SimpleDualBram_322_doutb;
  assign xil_SimpleDualBram_323_addra = _zz_addra_323[10:0];
  assign xil_SimpleDualBram_323_addrb = _zz_addrb_323[13:0];
  assign sData_fire_324 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_323_ena = (_zz_ena_323[0] && sData_fire_324);
  assign mData_323 = xil_SimpleDualBram_323_doutb;
  assign xil_SimpleDualBram_324_addra = _zz_addra_324[10:0];
  assign xil_SimpleDualBram_324_addrb = _zz_addrb_324[13:0];
  assign sData_fire_325 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_324_ena = (_zz_ena_324[0] && sData_fire_325);
  assign mData_324 = xil_SimpleDualBram_324_doutb;
  assign xil_SimpleDualBram_325_addra = _zz_addra_325[10:0];
  assign xil_SimpleDualBram_325_addrb = _zz_addrb_325[13:0];
  assign sData_fire_326 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_325_ena = (_zz_ena_325[0] && sData_fire_326);
  assign mData_325 = xil_SimpleDualBram_325_doutb;
  assign xil_SimpleDualBram_326_addra = _zz_addra_326[10:0];
  assign xil_SimpleDualBram_326_addrb = _zz_addrb_326[13:0];
  assign sData_fire_327 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_326_ena = (_zz_ena_326[0] && sData_fire_327);
  assign mData_326 = xil_SimpleDualBram_326_doutb;
  assign xil_SimpleDualBram_327_addra = _zz_addra_327[10:0];
  assign xil_SimpleDualBram_327_addrb = _zz_addrb_327[13:0];
  assign sData_fire_328 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_327_ena = (_zz_ena_327[0] && sData_fire_328);
  assign mData_327 = xil_SimpleDualBram_327_doutb;
  assign xil_SimpleDualBram_328_addra = _zz_addra_328[10:0];
  assign xil_SimpleDualBram_328_addrb = _zz_addrb_328[13:0];
  assign sData_fire_329 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_328_ena = (_zz_ena_328[0] && sData_fire_329);
  assign mData_328 = xil_SimpleDualBram_328_doutb;
  assign xil_SimpleDualBram_329_addra = _zz_addra_329[10:0];
  assign xil_SimpleDualBram_329_addrb = _zz_addrb_329[13:0];
  assign sData_fire_330 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_329_ena = (_zz_ena_329[0] && sData_fire_330);
  assign mData_329 = xil_SimpleDualBram_329_doutb;
  assign xil_SimpleDualBram_330_addra = _zz_addra_330[10:0];
  assign xil_SimpleDualBram_330_addrb = _zz_addrb_330[13:0];
  assign sData_fire_331 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_330_ena = (_zz_ena_330[0] && sData_fire_331);
  assign mData_330 = xil_SimpleDualBram_330_doutb;
  assign xil_SimpleDualBram_331_addra = _zz_addra_331[10:0];
  assign xil_SimpleDualBram_331_addrb = _zz_addrb_331[13:0];
  assign sData_fire_332 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_331_ena = (_zz_ena_331[0] && sData_fire_332);
  assign mData_331 = xil_SimpleDualBram_331_doutb;
  assign xil_SimpleDualBram_332_addra = _zz_addra_332[10:0];
  assign xil_SimpleDualBram_332_addrb = _zz_addrb_332[13:0];
  assign sData_fire_333 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_332_ena = (_zz_ena_332[0] && sData_fire_333);
  assign mData_332 = xil_SimpleDualBram_332_doutb;
  assign xil_SimpleDualBram_333_addra = _zz_addra_333[10:0];
  assign xil_SimpleDualBram_333_addrb = _zz_addrb_333[13:0];
  assign sData_fire_334 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_333_ena = (_zz_ena_333[0] && sData_fire_334);
  assign mData_333 = xil_SimpleDualBram_333_doutb;
  assign xil_SimpleDualBram_334_addra = _zz_addra_334[10:0];
  assign xil_SimpleDualBram_334_addrb = _zz_addrb_334[13:0];
  assign sData_fire_335 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_334_ena = (_zz_ena_334[0] && sData_fire_335);
  assign mData_334 = xil_SimpleDualBram_334_doutb;
  assign xil_SimpleDualBram_335_addra = _zz_addra_335[10:0];
  assign xil_SimpleDualBram_335_addrb = _zz_addrb_335[13:0];
  assign sData_fire_336 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_335_ena = (_zz_ena_335[0] && sData_fire_336);
  assign mData_335 = xil_SimpleDualBram_335_doutb;
  assign xil_SimpleDualBram_336_addra = _zz_addra_336[10:0];
  assign xil_SimpleDualBram_336_addrb = _zz_addrb_336[13:0];
  assign sData_fire_337 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_336_ena = (_zz_ena_336[0] && sData_fire_337);
  assign mData_336 = xil_SimpleDualBram_336_doutb;
  assign xil_SimpleDualBram_337_addra = _zz_addra_337[10:0];
  assign xil_SimpleDualBram_337_addrb = _zz_addrb_337[13:0];
  assign sData_fire_338 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_337_ena = (_zz_ena_337[0] && sData_fire_338);
  assign mData_337 = xil_SimpleDualBram_337_doutb;
  assign xil_SimpleDualBram_338_addra = _zz_addra_338[10:0];
  assign xil_SimpleDualBram_338_addrb = _zz_addrb_338[13:0];
  assign sData_fire_339 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_338_ena = (_zz_ena_338[0] && sData_fire_339);
  assign mData_338 = xil_SimpleDualBram_338_doutb;
  assign xil_SimpleDualBram_339_addra = _zz_addra_339[10:0];
  assign xil_SimpleDualBram_339_addrb = _zz_addrb_339[13:0];
  assign sData_fire_340 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_339_ena = (_zz_ena_339[0] && sData_fire_340);
  assign mData_339 = xil_SimpleDualBram_339_doutb;
  assign xil_SimpleDualBram_340_addra = _zz_addra_340[10:0];
  assign xil_SimpleDualBram_340_addrb = _zz_addrb_340[13:0];
  assign sData_fire_341 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_340_ena = (_zz_ena_340[0] && sData_fire_341);
  assign mData_340 = xil_SimpleDualBram_340_doutb;
  assign xil_SimpleDualBram_341_addra = _zz_addra_341[10:0];
  assign xil_SimpleDualBram_341_addrb = _zz_addrb_341[13:0];
  assign sData_fire_342 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_341_ena = (_zz_ena_341[0] && sData_fire_342);
  assign mData_341 = xil_SimpleDualBram_341_doutb;
  assign xil_SimpleDualBram_342_addra = _zz_addra_342[10:0];
  assign xil_SimpleDualBram_342_addrb = _zz_addrb_342[13:0];
  assign sData_fire_343 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_342_ena = (_zz_ena_342[0] && sData_fire_343);
  assign mData_342 = xil_SimpleDualBram_342_doutb;
  assign xil_SimpleDualBram_343_addra = _zz_addra_343[10:0];
  assign xil_SimpleDualBram_343_addrb = _zz_addrb_343[13:0];
  assign sData_fire_344 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_343_ena = (_zz_ena_343[0] && sData_fire_344);
  assign mData_343 = xil_SimpleDualBram_343_doutb;
  assign xil_SimpleDualBram_344_addra = _zz_addra_344[10:0];
  assign xil_SimpleDualBram_344_addrb = _zz_addrb_344[13:0];
  assign sData_fire_345 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_344_ena = (_zz_ena_344[0] && sData_fire_345);
  assign mData_344 = xil_SimpleDualBram_344_doutb;
  assign xil_SimpleDualBram_345_addra = _zz_addra_345[10:0];
  assign xil_SimpleDualBram_345_addrb = _zz_addrb_345[13:0];
  assign sData_fire_346 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_345_ena = (_zz_ena_345[0] && sData_fire_346);
  assign mData_345 = xil_SimpleDualBram_345_doutb;
  assign xil_SimpleDualBram_346_addra = _zz_addra_346[10:0];
  assign xil_SimpleDualBram_346_addrb = _zz_addrb_346[13:0];
  assign sData_fire_347 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_346_ena = (_zz_ena_346[0] && sData_fire_347);
  assign mData_346 = xil_SimpleDualBram_346_doutb;
  assign xil_SimpleDualBram_347_addra = _zz_addra_347[10:0];
  assign xil_SimpleDualBram_347_addrb = _zz_addrb_347[13:0];
  assign sData_fire_348 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_347_ena = (_zz_ena_347[0] && sData_fire_348);
  assign mData_347 = xil_SimpleDualBram_347_doutb;
  assign xil_SimpleDualBram_348_addra = _zz_addra_348[10:0];
  assign xil_SimpleDualBram_348_addrb = _zz_addrb_348[13:0];
  assign sData_fire_349 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_348_ena = (_zz_ena_348[0] && sData_fire_349);
  assign mData_348 = xil_SimpleDualBram_348_doutb;
  assign xil_SimpleDualBram_349_addra = _zz_addra_349[10:0];
  assign xil_SimpleDualBram_349_addrb = _zz_addrb_349[13:0];
  assign sData_fire_350 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_349_ena = (_zz_ena_349[0] && sData_fire_350);
  assign mData_349 = xil_SimpleDualBram_349_doutb;
  assign xil_SimpleDualBram_350_addra = _zz_addra_350[10:0];
  assign xil_SimpleDualBram_350_addrb = _zz_addrb_350[13:0];
  assign sData_fire_351 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_350_ena = (_zz_ena_350[0] && sData_fire_351);
  assign mData_350 = xil_SimpleDualBram_350_doutb;
  assign xil_SimpleDualBram_351_addra = _zz_addra_351[10:0];
  assign xil_SimpleDualBram_351_addrb = _zz_addrb_351[13:0];
  assign sData_fire_352 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_351_ena = (_zz_ena_351[0] && sData_fire_352);
  assign mData_351 = xil_SimpleDualBram_351_doutb;
  assign xil_SimpleDualBram_352_addra = _zz_addra_352[10:0];
  assign xil_SimpleDualBram_352_addrb = _zz_addrb_352[13:0];
  assign sData_fire_353 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_352_ena = (_zz_ena_352[0] && sData_fire_353);
  assign mData_352 = xil_SimpleDualBram_352_doutb;
  assign xil_SimpleDualBram_353_addra = _zz_addra_353[10:0];
  assign xil_SimpleDualBram_353_addrb = _zz_addrb_353[13:0];
  assign sData_fire_354 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_353_ena = (_zz_ena_353[0] && sData_fire_354);
  assign mData_353 = xil_SimpleDualBram_353_doutb;
  assign xil_SimpleDualBram_354_addra = _zz_addra_354[10:0];
  assign xil_SimpleDualBram_354_addrb = _zz_addrb_354[13:0];
  assign sData_fire_355 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_354_ena = (_zz_ena_354[0] && sData_fire_355);
  assign mData_354 = xil_SimpleDualBram_354_doutb;
  assign xil_SimpleDualBram_355_addra = _zz_addra_355[10:0];
  assign xil_SimpleDualBram_355_addrb = _zz_addrb_355[13:0];
  assign sData_fire_356 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_355_ena = (_zz_ena_355[0] && sData_fire_356);
  assign mData_355 = xil_SimpleDualBram_355_doutb;
  assign xil_SimpleDualBram_356_addra = _zz_addra_356[10:0];
  assign xil_SimpleDualBram_356_addrb = _zz_addrb_356[13:0];
  assign sData_fire_357 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_356_ena = (_zz_ena_356[0] && sData_fire_357);
  assign mData_356 = xil_SimpleDualBram_356_doutb;
  assign xil_SimpleDualBram_357_addra = _zz_addra_357[10:0];
  assign xil_SimpleDualBram_357_addrb = _zz_addrb_357[13:0];
  assign sData_fire_358 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_357_ena = (_zz_ena_357[0] && sData_fire_358);
  assign mData_357 = xil_SimpleDualBram_357_doutb;
  assign xil_SimpleDualBram_358_addra = _zz_addra_358[10:0];
  assign xil_SimpleDualBram_358_addrb = _zz_addrb_358[13:0];
  assign sData_fire_359 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_358_ena = (_zz_ena_358[0] && sData_fire_359);
  assign mData_358 = xil_SimpleDualBram_358_doutb;
  assign xil_SimpleDualBram_359_addra = _zz_addra_359[10:0];
  assign xil_SimpleDualBram_359_addrb = _zz_addrb_359[13:0];
  assign sData_fire_360 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_359_ena = (_zz_ena_359[0] && sData_fire_360);
  assign mData_359 = xil_SimpleDualBram_359_doutb;
  assign xil_SimpleDualBram_360_addra = _zz_addra_360[10:0];
  assign xil_SimpleDualBram_360_addrb = _zz_addrb_360[13:0];
  assign sData_fire_361 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_360_ena = (_zz_ena_360[0] && sData_fire_361);
  assign mData_360 = xil_SimpleDualBram_360_doutb;
  assign xil_SimpleDualBram_361_addra = _zz_addra_361[10:0];
  assign xil_SimpleDualBram_361_addrb = _zz_addrb_361[13:0];
  assign sData_fire_362 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_361_ena = (_zz_ena_361[0] && sData_fire_362);
  assign mData_361 = xil_SimpleDualBram_361_doutb;
  assign xil_SimpleDualBram_362_addra = _zz_addra_362[10:0];
  assign xil_SimpleDualBram_362_addrb = _zz_addrb_362[13:0];
  assign sData_fire_363 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_362_ena = (_zz_ena_362[0] && sData_fire_363);
  assign mData_362 = xil_SimpleDualBram_362_doutb;
  assign xil_SimpleDualBram_363_addra = _zz_addra_363[10:0];
  assign xil_SimpleDualBram_363_addrb = _zz_addrb_363[13:0];
  assign sData_fire_364 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_363_ena = (_zz_ena_363[0] && sData_fire_364);
  assign mData_363 = xil_SimpleDualBram_363_doutb;
  assign xil_SimpleDualBram_364_addra = _zz_addra_364[10:0];
  assign xil_SimpleDualBram_364_addrb = _zz_addrb_364[13:0];
  assign sData_fire_365 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_364_ena = (_zz_ena_364[0] && sData_fire_365);
  assign mData_364 = xil_SimpleDualBram_364_doutb;
  assign xil_SimpleDualBram_365_addra = _zz_addra_365[10:0];
  assign xil_SimpleDualBram_365_addrb = _zz_addrb_365[13:0];
  assign sData_fire_366 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_365_ena = (_zz_ena_365[0] && sData_fire_366);
  assign mData_365 = xil_SimpleDualBram_365_doutb;
  assign xil_SimpleDualBram_366_addra = _zz_addra_366[10:0];
  assign xil_SimpleDualBram_366_addrb = _zz_addrb_366[13:0];
  assign sData_fire_367 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_366_ena = (_zz_ena_366[0] && sData_fire_367);
  assign mData_366 = xil_SimpleDualBram_366_doutb;
  assign xil_SimpleDualBram_367_addra = _zz_addra_367[10:0];
  assign xil_SimpleDualBram_367_addrb = _zz_addrb_367[13:0];
  assign sData_fire_368 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_367_ena = (_zz_ena_367[0] && sData_fire_368);
  assign mData_367 = xil_SimpleDualBram_367_doutb;
  assign xil_SimpleDualBram_368_addra = _zz_addra_368[10:0];
  assign xil_SimpleDualBram_368_addrb = _zz_addrb_368[13:0];
  assign sData_fire_369 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_368_ena = (_zz_ena_368[0] && sData_fire_369);
  assign mData_368 = xil_SimpleDualBram_368_doutb;
  assign xil_SimpleDualBram_369_addra = _zz_addra_369[10:0];
  assign xil_SimpleDualBram_369_addrb = _zz_addrb_369[13:0];
  assign sData_fire_370 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_369_ena = (_zz_ena_369[0] && sData_fire_370);
  assign mData_369 = xil_SimpleDualBram_369_doutb;
  assign xil_SimpleDualBram_370_addra = _zz_addra_370[10:0];
  assign xil_SimpleDualBram_370_addrb = _zz_addrb_370[13:0];
  assign sData_fire_371 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_370_ena = (_zz_ena_370[0] && sData_fire_371);
  assign mData_370 = xil_SimpleDualBram_370_doutb;
  assign xil_SimpleDualBram_371_addra = _zz_addra_371[10:0];
  assign xil_SimpleDualBram_371_addrb = _zz_addrb_371[13:0];
  assign sData_fire_372 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_371_ena = (_zz_ena_371[0] && sData_fire_372);
  assign mData_371 = xil_SimpleDualBram_371_doutb;
  assign xil_SimpleDualBram_372_addra = _zz_addra_372[10:0];
  assign xil_SimpleDualBram_372_addrb = _zz_addrb_372[13:0];
  assign sData_fire_373 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_372_ena = (_zz_ena_372[0] && sData_fire_373);
  assign mData_372 = xil_SimpleDualBram_372_doutb;
  assign xil_SimpleDualBram_373_addra = _zz_addra_373[10:0];
  assign xil_SimpleDualBram_373_addrb = _zz_addrb_373[13:0];
  assign sData_fire_374 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_373_ena = (_zz_ena_373[0] && sData_fire_374);
  assign mData_373 = xil_SimpleDualBram_373_doutb;
  assign xil_SimpleDualBram_374_addra = _zz_addra_374[10:0];
  assign xil_SimpleDualBram_374_addrb = _zz_addrb_374[13:0];
  assign sData_fire_375 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_374_ena = (_zz_ena_374[0] && sData_fire_375);
  assign mData_374 = xil_SimpleDualBram_374_doutb;
  assign xil_SimpleDualBram_375_addra = _zz_addra_375[10:0];
  assign xil_SimpleDualBram_375_addrb = _zz_addrb_375[13:0];
  assign sData_fire_376 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_375_ena = (_zz_ena_375[0] && sData_fire_376);
  assign mData_375 = xil_SimpleDualBram_375_doutb;
  assign xil_SimpleDualBram_376_addra = _zz_addra_376[10:0];
  assign xil_SimpleDualBram_376_addrb = _zz_addrb_376[13:0];
  assign sData_fire_377 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_376_ena = (_zz_ena_376[0] && sData_fire_377);
  assign mData_376 = xil_SimpleDualBram_376_doutb;
  assign xil_SimpleDualBram_377_addra = _zz_addra_377[10:0];
  assign xil_SimpleDualBram_377_addrb = _zz_addrb_377[13:0];
  assign sData_fire_378 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_377_ena = (_zz_ena_377[0] && sData_fire_378);
  assign mData_377 = xil_SimpleDualBram_377_doutb;
  assign xil_SimpleDualBram_378_addra = _zz_addra_378[10:0];
  assign xil_SimpleDualBram_378_addrb = _zz_addrb_378[13:0];
  assign sData_fire_379 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_378_ena = (_zz_ena_378[0] && sData_fire_379);
  assign mData_378 = xil_SimpleDualBram_378_doutb;
  assign xil_SimpleDualBram_379_addra = _zz_addra_379[10:0];
  assign xil_SimpleDualBram_379_addrb = _zz_addrb_379[13:0];
  assign sData_fire_380 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_379_ena = (_zz_ena_379[0] && sData_fire_380);
  assign mData_379 = xil_SimpleDualBram_379_doutb;
  assign xil_SimpleDualBram_380_addra = _zz_addra_380[10:0];
  assign xil_SimpleDualBram_380_addrb = _zz_addrb_380[13:0];
  assign sData_fire_381 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_380_ena = (_zz_ena_380[0] && sData_fire_381);
  assign mData_380 = xil_SimpleDualBram_380_doutb;
  assign xil_SimpleDualBram_381_addra = _zz_addra_381[10:0];
  assign xil_SimpleDualBram_381_addrb = _zz_addrb_381[13:0];
  assign sData_fire_382 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_381_ena = (_zz_ena_381[0] && sData_fire_382);
  assign mData_381 = xil_SimpleDualBram_381_doutb;
  assign xil_SimpleDualBram_382_addra = _zz_addra_382[10:0];
  assign xil_SimpleDualBram_382_addrb = _zz_addrb_382[13:0];
  assign sData_fire_383 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_382_ena = (_zz_ena_382[0] && sData_fire_383);
  assign mData_382 = xil_SimpleDualBram_382_doutb;
  assign xil_SimpleDualBram_383_addra = _zz_addra_383[10:0];
  assign xil_SimpleDualBram_383_addrb = _zz_addrb_383[13:0];
  assign sData_fire_384 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_383_ena = (_zz_ena_383[0] && sData_fire_384);
  assign mData_383 = xil_SimpleDualBram_383_doutb;
  assign xil_SimpleDualBram_384_addra = _zz_addra_384[10:0];
  assign xil_SimpleDualBram_384_addrb = _zz_addrb_384[13:0];
  assign sData_fire_385 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_384_ena = (_zz_ena_384[0] && sData_fire_385);
  assign mData_384 = xil_SimpleDualBram_384_doutb;
  assign xil_SimpleDualBram_385_addra = _zz_addra_385[10:0];
  assign xil_SimpleDualBram_385_addrb = _zz_addrb_385[13:0];
  assign sData_fire_386 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_385_ena = (_zz_ena_385[0] && sData_fire_386);
  assign mData_385 = xil_SimpleDualBram_385_doutb;
  assign xil_SimpleDualBram_386_addra = _zz_addra_386[10:0];
  assign xil_SimpleDualBram_386_addrb = _zz_addrb_386[13:0];
  assign sData_fire_387 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_386_ena = (_zz_ena_386[0] && sData_fire_387);
  assign mData_386 = xil_SimpleDualBram_386_doutb;
  assign xil_SimpleDualBram_387_addra = _zz_addra_387[10:0];
  assign xil_SimpleDualBram_387_addrb = _zz_addrb_387[13:0];
  assign sData_fire_388 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_387_ena = (_zz_ena_387[0] && sData_fire_388);
  assign mData_387 = xil_SimpleDualBram_387_doutb;
  assign xil_SimpleDualBram_388_addra = _zz_addra_388[10:0];
  assign xil_SimpleDualBram_388_addrb = _zz_addrb_388[13:0];
  assign sData_fire_389 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_388_ena = (_zz_ena_388[0] && sData_fire_389);
  assign mData_388 = xil_SimpleDualBram_388_doutb;
  assign xil_SimpleDualBram_389_addra = _zz_addra_389[10:0];
  assign xil_SimpleDualBram_389_addrb = _zz_addrb_389[13:0];
  assign sData_fire_390 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_389_ena = (_zz_ena_389[0] && sData_fire_390);
  assign mData_389 = xil_SimpleDualBram_389_doutb;
  assign xil_SimpleDualBram_390_addra = _zz_addra_390[10:0];
  assign xil_SimpleDualBram_390_addrb = _zz_addrb_390[13:0];
  assign sData_fire_391 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_390_ena = (_zz_ena_390[0] && sData_fire_391);
  assign mData_390 = xil_SimpleDualBram_390_doutb;
  assign xil_SimpleDualBram_391_addra = _zz_addra_391[10:0];
  assign xil_SimpleDualBram_391_addrb = _zz_addrb_391[13:0];
  assign sData_fire_392 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_391_ena = (_zz_ena_391[0] && sData_fire_392);
  assign mData_391 = xil_SimpleDualBram_391_doutb;
  assign xil_SimpleDualBram_392_addra = _zz_addra_392[10:0];
  assign xil_SimpleDualBram_392_addrb = _zz_addrb_392[13:0];
  assign sData_fire_393 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_392_ena = (_zz_ena_392[0] && sData_fire_393);
  assign mData_392 = xil_SimpleDualBram_392_doutb;
  assign xil_SimpleDualBram_393_addra = _zz_addra_393[10:0];
  assign xil_SimpleDualBram_393_addrb = _zz_addrb_393[13:0];
  assign sData_fire_394 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_393_ena = (_zz_ena_393[0] && sData_fire_394);
  assign mData_393 = xil_SimpleDualBram_393_doutb;
  assign xil_SimpleDualBram_394_addra = _zz_addra_394[10:0];
  assign xil_SimpleDualBram_394_addrb = _zz_addrb_394[13:0];
  assign sData_fire_395 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_394_ena = (_zz_ena_394[0] && sData_fire_395);
  assign mData_394 = xil_SimpleDualBram_394_doutb;
  assign xil_SimpleDualBram_395_addra = _zz_addra_395[10:0];
  assign xil_SimpleDualBram_395_addrb = _zz_addrb_395[13:0];
  assign sData_fire_396 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_395_ena = (_zz_ena_395[0] && sData_fire_396);
  assign mData_395 = xil_SimpleDualBram_395_doutb;
  assign xil_SimpleDualBram_396_addra = _zz_addra_396[10:0];
  assign xil_SimpleDualBram_396_addrb = _zz_addrb_396[13:0];
  assign sData_fire_397 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_396_ena = (_zz_ena_396[0] && sData_fire_397);
  assign mData_396 = xil_SimpleDualBram_396_doutb;
  assign xil_SimpleDualBram_397_addra = _zz_addra_397[10:0];
  assign xil_SimpleDualBram_397_addrb = _zz_addrb_397[13:0];
  assign sData_fire_398 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_397_ena = (_zz_ena_397[0] && sData_fire_398);
  assign mData_397 = xil_SimpleDualBram_397_doutb;
  assign xil_SimpleDualBram_398_addra = _zz_addra_398[10:0];
  assign xil_SimpleDualBram_398_addrb = _zz_addrb_398[13:0];
  assign sData_fire_399 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_398_ena = (_zz_ena_398[0] && sData_fire_399);
  assign mData_398 = xil_SimpleDualBram_398_doutb;
  assign xil_SimpleDualBram_399_addra = _zz_addra_399[10:0];
  assign xil_SimpleDualBram_399_addrb = _zz_addrb_399[13:0];
  assign sData_fire_400 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_399_ena = (_zz_ena_399[0] && sData_fire_400);
  assign mData_399 = xil_SimpleDualBram_399_doutb;
  assign xil_SimpleDualBram_400_addra = _zz_addra_400[10:0];
  assign xil_SimpleDualBram_400_addrb = _zz_addrb_400[13:0];
  assign sData_fire_401 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_400_ena = (_zz_ena_400[0] && sData_fire_401);
  assign mData_400 = xil_SimpleDualBram_400_doutb;
  assign xil_SimpleDualBram_401_addra = _zz_addra_401[10:0];
  assign xil_SimpleDualBram_401_addrb = _zz_addrb_401[13:0];
  assign sData_fire_402 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_401_ena = (_zz_ena_401[0] && sData_fire_402);
  assign mData_401 = xil_SimpleDualBram_401_doutb;
  assign xil_SimpleDualBram_402_addra = _zz_addra_402[10:0];
  assign xil_SimpleDualBram_402_addrb = _zz_addrb_402[13:0];
  assign sData_fire_403 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_402_ena = (_zz_ena_402[0] && sData_fire_403);
  assign mData_402 = xil_SimpleDualBram_402_doutb;
  assign xil_SimpleDualBram_403_addra = _zz_addra_403[10:0];
  assign xil_SimpleDualBram_403_addrb = _zz_addrb_403[13:0];
  assign sData_fire_404 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_403_ena = (_zz_ena_403[0] && sData_fire_404);
  assign mData_403 = xil_SimpleDualBram_403_doutb;
  assign xil_SimpleDualBram_404_addra = _zz_addra_404[10:0];
  assign xil_SimpleDualBram_404_addrb = _zz_addrb_404[13:0];
  assign sData_fire_405 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_404_ena = (_zz_ena_404[0] && sData_fire_405);
  assign mData_404 = xil_SimpleDualBram_404_doutb;
  assign xil_SimpleDualBram_405_addra = _zz_addra_405[10:0];
  assign xil_SimpleDualBram_405_addrb = _zz_addrb_405[13:0];
  assign sData_fire_406 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_405_ena = (_zz_ena_405[0] && sData_fire_406);
  assign mData_405 = xil_SimpleDualBram_405_doutb;
  assign xil_SimpleDualBram_406_addra = _zz_addra_406[10:0];
  assign xil_SimpleDualBram_406_addrb = _zz_addrb_406[13:0];
  assign sData_fire_407 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_406_ena = (_zz_ena_406[0] && sData_fire_407);
  assign mData_406 = xil_SimpleDualBram_406_doutb;
  assign xil_SimpleDualBram_407_addra = _zz_addra_407[10:0];
  assign xil_SimpleDualBram_407_addrb = _zz_addrb_407[13:0];
  assign sData_fire_408 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_407_ena = (_zz_ena_407[0] && sData_fire_408);
  assign mData_407 = xil_SimpleDualBram_407_doutb;
  assign xil_SimpleDualBram_408_addra = _zz_addra_408[10:0];
  assign xil_SimpleDualBram_408_addrb = _zz_addrb_408[13:0];
  assign sData_fire_409 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_408_ena = (_zz_ena_408[0] && sData_fire_409);
  assign mData_408 = xil_SimpleDualBram_408_doutb;
  assign xil_SimpleDualBram_409_addra = _zz_addra_409[10:0];
  assign xil_SimpleDualBram_409_addrb = _zz_addrb_409[13:0];
  assign sData_fire_410 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_409_ena = (_zz_ena_409[0] && sData_fire_410);
  assign mData_409 = xil_SimpleDualBram_409_doutb;
  assign xil_SimpleDualBram_410_addra = _zz_addra_410[10:0];
  assign xil_SimpleDualBram_410_addrb = _zz_addrb_410[13:0];
  assign sData_fire_411 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_410_ena = (_zz_ena_410[0] && sData_fire_411);
  assign mData_410 = xil_SimpleDualBram_410_doutb;
  assign xil_SimpleDualBram_411_addra = _zz_addra_411[10:0];
  assign xil_SimpleDualBram_411_addrb = _zz_addrb_411[13:0];
  assign sData_fire_412 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_411_ena = (_zz_ena_411[0] && sData_fire_412);
  assign mData_411 = xil_SimpleDualBram_411_doutb;
  assign xil_SimpleDualBram_412_addra = _zz_addra_412[10:0];
  assign xil_SimpleDualBram_412_addrb = _zz_addrb_412[13:0];
  assign sData_fire_413 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_412_ena = (_zz_ena_412[0] && sData_fire_413);
  assign mData_412 = xil_SimpleDualBram_412_doutb;
  assign xil_SimpleDualBram_413_addra = _zz_addra_413[10:0];
  assign xil_SimpleDualBram_413_addrb = _zz_addrb_413[13:0];
  assign sData_fire_414 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_413_ena = (_zz_ena_413[0] && sData_fire_414);
  assign mData_413 = xil_SimpleDualBram_413_doutb;
  assign xil_SimpleDualBram_414_addra = _zz_addra_414[10:0];
  assign xil_SimpleDualBram_414_addrb = _zz_addrb_414[13:0];
  assign sData_fire_415 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_414_ena = (_zz_ena_414[0] && sData_fire_415);
  assign mData_414 = xil_SimpleDualBram_414_doutb;
  assign xil_SimpleDualBram_415_addra = _zz_addra_415[10:0];
  assign xil_SimpleDualBram_415_addrb = _zz_addrb_415[13:0];
  assign sData_fire_416 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_415_ena = (_zz_ena_415[0] && sData_fire_416);
  assign mData_415 = xil_SimpleDualBram_415_doutb;
  assign xil_SimpleDualBram_416_addra = _zz_addra_416[10:0];
  assign xil_SimpleDualBram_416_addrb = _zz_addrb_416[13:0];
  assign sData_fire_417 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_416_ena = (_zz_ena_416[0] && sData_fire_417);
  assign mData_416 = xil_SimpleDualBram_416_doutb;
  assign xil_SimpleDualBram_417_addra = _zz_addra_417[10:0];
  assign xil_SimpleDualBram_417_addrb = _zz_addrb_417[13:0];
  assign sData_fire_418 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_417_ena = (_zz_ena_417[0] && sData_fire_418);
  assign mData_417 = xil_SimpleDualBram_417_doutb;
  assign xil_SimpleDualBram_418_addra = _zz_addra_418[10:0];
  assign xil_SimpleDualBram_418_addrb = _zz_addrb_418[13:0];
  assign sData_fire_419 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_418_ena = (_zz_ena_418[0] && sData_fire_419);
  assign mData_418 = xil_SimpleDualBram_418_doutb;
  assign xil_SimpleDualBram_419_addra = _zz_addra_419[10:0];
  assign xil_SimpleDualBram_419_addrb = _zz_addrb_419[13:0];
  assign sData_fire_420 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_419_ena = (_zz_ena_419[0] && sData_fire_420);
  assign mData_419 = xil_SimpleDualBram_419_doutb;
  assign xil_SimpleDualBram_420_addra = _zz_addra_420[10:0];
  assign xil_SimpleDualBram_420_addrb = _zz_addrb_420[13:0];
  assign sData_fire_421 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_420_ena = (_zz_ena_420[0] && sData_fire_421);
  assign mData_420 = xil_SimpleDualBram_420_doutb;
  assign xil_SimpleDualBram_421_addra = _zz_addra_421[10:0];
  assign xil_SimpleDualBram_421_addrb = _zz_addrb_421[13:0];
  assign sData_fire_422 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_421_ena = (_zz_ena_421[0] && sData_fire_422);
  assign mData_421 = xil_SimpleDualBram_421_doutb;
  assign xil_SimpleDualBram_422_addra = _zz_addra_422[10:0];
  assign xil_SimpleDualBram_422_addrb = _zz_addrb_422[13:0];
  assign sData_fire_423 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_422_ena = (_zz_ena_422[0] && sData_fire_423);
  assign mData_422 = xil_SimpleDualBram_422_doutb;
  assign xil_SimpleDualBram_423_addra = _zz_addra_423[10:0];
  assign xil_SimpleDualBram_423_addrb = _zz_addrb_423[13:0];
  assign sData_fire_424 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_423_ena = (_zz_ena_423[0] && sData_fire_424);
  assign mData_423 = xil_SimpleDualBram_423_doutb;
  assign xil_SimpleDualBram_424_addra = _zz_addra_424[10:0];
  assign xil_SimpleDualBram_424_addrb = _zz_addrb_424[13:0];
  assign sData_fire_425 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_424_ena = (_zz_ena_424[0] && sData_fire_425);
  assign mData_424 = xil_SimpleDualBram_424_doutb;
  assign xil_SimpleDualBram_425_addra = _zz_addra_425[10:0];
  assign xil_SimpleDualBram_425_addrb = _zz_addrb_425[13:0];
  assign sData_fire_426 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_425_ena = (_zz_ena_425[0] && sData_fire_426);
  assign mData_425 = xil_SimpleDualBram_425_doutb;
  assign xil_SimpleDualBram_426_addra = _zz_addra_426[10:0];
  assign xil_SimpleDualBram_426_addrb = _zz_addrb_426[13:0];
  assign sData_fire_427 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_426_ena = (_zz_ena_426[0] && sData_fire_427);
  assign mData_426 = xil_SimpleDualBram_426_doutb;
  assign xil_SimpleDualBram_427_addra = _zz_addra_427[10:0];
  assign xil_SimpleDualBram_427_addrb = _zz_addrb_427[13:0];
  assign sData_fire_428 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_427_ena = (_zz_ena_427[0] && sData_fire_428);
  assign mData_427 = xil_SimpleDualBram_427_doutb;
  assign xil_SimpleDualBram_428_addra = _zz_addra_428[10:0];
  assign xil_SimpleDualBram_428_addrb = _zz_addrb_428[13:0];
  assign sData_fire_429 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_428_ena = (_zz_ena_428[0] && sData_fire_429);
  assign mData_428 = xil_SimpleDualBram_428_doutb;
  assign xil_SimpleDualBram_429_addra = _zz_addra_429[10:0];
  assign xil_SimpleDualBram_429_addrb = _zz_addrb_429[13:0];
  assign sData_fire_430 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_429_ena = (_zz_ena_429[0] && sData_fire_430);
  assign mData_429 = xil_SimpleDualBram_429_doutb;
  assign xil_SimpleDualBram_430_addra = _zz_addra_430[10:0];
  assign xil_SimpleDualBram_430_addrb = _zz_addrb_430[13:0];
  assign sData_fire_431 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_430_ena = (_zz_ena_430[0] && sData_fire_431);
  assign mData_430 = xil_SimpleDualBram_430_doutb;
  assign xil_SimpleDualBram_431_addra = _zz_addra_431[10:0];
  assign xil_SimpleDualBram_431_addrb = _zz_addrb_431[13:0];
  assign sData_fire_432 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_431_ena = (_zz_ena_431[0] && sData_fire_432);
  assign mData_431 = xil_SimpleDualBram_431_doutb;
  assign xil_SimpleDualBram_432_addra = _zz_addra_432[10:0];
  assign xil_SimpleDualBram_432_addrb = _zz_addrb_432[13:0];
  assign sData_fire_433 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_432_ena = (_zz_ena_432[0] && sData_fire_433);
  assign mData_432 = xil_SimpleDualBram_432_doutb;
  assign xil_SimpleDualBram_433_addra = _zz_addra_433[10:0];
  assign xil_SimpleDualBram_433_addrb = _zz_addrb_433[13:0];
  assign sData_fire_434 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_433_ena = (_zz_ena_433[0] && sData_fire_434);
  assign mData_433 = xil_SimpleDualBram_433_doutb;
  assign xil_SimpleDualBram_434_addra = _zz_addra_434[10:0];
  assign xil_SimpleDualBram_434_addrb = _zz_addrb_434[13:0];
  assign sData_fire_435 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_434_ena = (_zz_ena_434[0] && sData_fire_435);
  assign mData_434 = xil_SimpleDualBram_434_doutb;
  assign xil_SimpleDualBram_435_addra = _zz_addra_435[10:0];
  assign xil_SimpleDualBram_435_addrb = _zz_addrb_435[13:0];
  assign sData_fire_436 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_435_ena = (_zz_ena_435[0] && sData_fire_436);
  assign mData_435 = xil_SimpleDualBram_435_doutb;
  assign xil_SimpleDualBram_436_addra = _zz_addra_436[10:0];
  assign xil_SimpleDualBram_436_addrb = _zz_addrb_436[13:0];
  assign sData_fire_437 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_436_ena = (_zz_ena_436[0] && sData_fire_437);
  assign mData_436 = xil_SimpleDualBram_436_doutb;
  assign xil_SimpleDualBram_437_addra = _zz_addra_437[10:0];
  assign xil_SimpleDualBram_437_addrb = _zz_addrb_437[13:0];
  assign sData_fire_438 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_437_ena = (_zz_ena_437[0] && sData_fire_438);
  assign mData_437 = xil_SimpleDualBram_437_doutb;
  assign xil_SimpleDualBram_438_addra = _zz_addra_438[10:0];
  assign xil_SimpleDualBram_438_addrb = _zz_addrb_438[13:0];
  assign sData_fire_439 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_438_ena = (_zz_ena_438[0] && sData_fire_439);
  assign mData_438 = xil_SimpleDualBram_438_doutb;
  assign xil_SimpleDualBram_439_addra = _zz_addra_439[10:0];
  assign xil_SimpleDualBram_439_addrb = _zz_addrb_439[13:0];
  assign sData_fire_440 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_439_ena = (_zz_ena_439[0] && sData_fire_440);
  assign mData_439 = xil_SimpleDualBram_439_doutb;
  assign xil_SimpleDualBram_440_addra = _zz_addra_440[10:0];
  assign xil_SimpleDualBram_440_addrb = _zz_addrb_440[13:0];
  assign sData_fire_441 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_440_ena = (_zz_ena_440[0] && sData_fire_441);
  assign mData_440 = xil_SimpleDualBram_440_doutb;
  assign xil_SimpleDualBram_441_addra = _zz_addra_441[10:0];
  assign xil_SimpleDualBram_441_addrb = _zz_addrb_441[13:0];
  assign sData_fire_442 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_441_ena = (_zz_ena_441[0] && sData_fire_442);
  assign mData_441 = xil_SimpleDualBram_441_doutb;
  assign xil_SimpleDualBram_442_addra = _zz_addra_442[10:0];
  assign xil_SimpleDualBram_442_addrb = _zz_addrb_442[13:0];
  assign sData_fire_443 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_442_ena = (_zz_ena_442[0] && sData_fire_443);
  assign mData_442 = xil_SimpleDualBram_442_doutb;
  assign xil_SimpleDualBram_443_addra = _zz_addra_443[10:0];
  assign xil_SimpleDualBram_443_addrb = _zz_addrb_443[13:0];
  assign sData_fire_444 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_443_ena = (_zz_ena_443[0] && sData_fire_444);
  assign mData_443 = xil_SimpleDualBram_443_doutb;
  assign xil_SimpleDualBram_444_addra = _zz_addra_444[10:0];
  assign xil_SimpleDualBram_444_addrb = _zz_addrb_444[13:0];
  assign sData_fire_445 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_444_ena = (_zz_ena_444[0] && sData_fire_445);
  assign mData_444 = xil_SimpleDualBram_444_doutb;
  assign xil_SimpleDualBram_445_addra = _zz_addra_445[10:0];
  assign xil_SimpleDualBram_445_addrb = _zz_addrb_445[13:0];
  assign sData_fire_446 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_445_ena = (_zz_ena_445[0] && sData_fire_446);
  assign mData_445 = xil_SimpleDualBram_445_doutb;
  assign xil_SimpleDualBram_446_addra = _zz_addra_446[10:0];
  assign xil_SimpleDualBram_446_addrb = _zz_addrb_446[13:0];
  assign sData_fire_447 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_446_ena = (_zz_ena_446[0] && sData_fire_447);
  assign mData_446 = xil_SimpleDualBram_446_doutb;
  assign xil_SimpleDualBram_447_addra = _zz_addra_447[10:0];
  assign xil_SimpleDualBram_447_addrb = _zz_addrb_447[13:0];
  assign sData_fire_448 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_447_ena = (_zz_ena_447[0] && sData_fire_448);
  assign mData_447 = xil_SimpleDualBram_447_doutb;
  assign xil_SimpleDualBram_448_addra = _zz_addra_448[10:0];
  assign xil_SimpleDualBram_448_addrb = _zz_addrb_448[13:0];
  assign sData_fire_449 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_448_ena = (_zz_ena_448[0] && sData_fire_449);
  assign mData_448 = xil_SimpleDualBram_448_doutb;
  assign xil_SimpleDualBram_449_addra = _zz_addra_449[10:0];
  assign xil_SimpleDualBram_449_addrb = _zz_addrb_449[13:0];
  assign sData_fire_450 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_449_ena = (_zz_ena_449[0] && sData_fire_450);
  assign mData_449 = xil_SimpleDualBram_449_doutb;
  assign xil_SimpleDualBram_450_addra = _zz_addra_450[10:0];
  assign xil_SimpleDualBram_450_addrb = _zz_addrb_450[13:0];
  assign sData_fire_451 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_450_ena = (_zz_ena_450[0] && sData_fire_451);
  assign mData_450 = xil_SimpleDualBram_450_doutb;
  assign xil_SimpleDualBram_451_addra = _zz_addra_451[10:0];
  assign xil_SimpleDualBram_451_addrb = _zz_addrb_451[13:0];
  assign sData_fire_452 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_451_ena = (_zz_ena_451[0] && sData_fire_452);
  assign mData_451 = xil_SimpleDualBram_451_doutb;
  assign xil_SimpleDualBram_452_addra = _zz_addra_452[10:0];
  assign xil_SimpleDualBram_452_addrb = _zz_addrb_452[13:0];
  assign sData_fire_453 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_452_ena = (_zz_ena_452[0] && sData_fire_453);
  assign mData_452 = xil_SimpleDualBram_452_doutb;
  assign xil_SimpleDualBram_453_addra = _zz_addra_453[10:0];
  assign xil_SimpleDualBram_453_addrb = _zz_addrb_453[13:0];
  assign sData_fire_454 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_453_ena = (_zz_ena_453[0] && sData_fire_454);
  assign mData_453 = xil_SimpleDualBram_453_doutb;
  assign xil_SimpleDualBram_454_addra = _zz_addra_454[10:0];
  assign xil_SimpleDualBram_454_addrb = _zz_addrb_454[13:0];
  assign sData_fire_455 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_454_ena = (_zz_ena_454[0] && sData_fire_455);
  assign mData_454 = xil_SimpleDualBram_454_doutb;
  assign xil_SimpleDualBram_455_addra = _zz_addra_455[10:0];
  assign xil_SimpleDualBram_455_addrb = _zz_addrb_455[13:0];
  assign sData_fire_456 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_455_ena = (_zz_ena_455[0] && sData_fire_456);
  assign mData_455 = xil_SimpleDualBram_455_doutb;
  assign xil_SimpleDualBram_456_addra = _zz_addra_456[10:0];
  assign xil_SimpleDualBram_456_addrb = _zz_addrb_456[13:0];
  assign sData_fire_457 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_456_ena = (_zz_ena_456[0] && sData_fire_457);
  assign mData_456 = xil_SimpleDualBram_456_doutb;
  assign xil_SimpleDualBram_457_addra = _zz_addra_457[10:0];
  assign xil_SimpleDualBram_457_addrb = _zz_addrb_457[13:0];
  assign sData_fire_458 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_457_ena = (_zz_ena_457[0] && sData_fire_458);
  assign mData_457 = xil_SimpleDualBram_457_doutb;
  assign xil_SimpleDualBram_458_addra = _zz_addra_458[10:0];
  assign xil_SimpleDualBram_458_addrb = _zz_addrb_458[13:0];
  assign sData_fire_459 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_458_ena = (_zz_ena_458[0] && sData_fire_459);
  assign mData_458 = xil_SimpleDualBram_458_doutb;
  assign xil_SimpleDualBram_459_addra = _zz_addra_459[10:0];
  assign xil_SimpleDualBram_459_addrb = _zz_addrb_459[13:0];
  assign sData_fire_460 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_459_ena = (_zz_ena_459[0] && sData_fire_460);
  assign mData_459 = xil_SimpleDualBram_459_doutb;
  assign xil_SimpleDualBram_460_addra = _zz_addra_460[10:0];
  assign xil_SimpleDualBram_460_addrb = _zz_addrb_460[13:0];
  assign sData_fire_461 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_460_ena = (_zz_ena_460[0] && sData_fire_461);
  assign mData_460 = xil_SimpleDualBram_460_doutb;
  assign xil_SimpleDualBram_461_addra = _zz_addra_461[10:0];
  assign xil_SimpleDualBram_461_addrb = _zz_addrb_461[13:0];
  assign sData_fire_462 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_461_ena = (_zz_ena_461[0] && sData_fire_462);
  assign mData_461 = xil_SimpleDualBram_461_doutb;
  assign xil_SimpleDualBram_462_addra = _zz_addra_462[10:0];
  assign xil_SimpleDualBram_462_addrb = _zz_addrb_462[13:0];
  assign sData_fire_463 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_462_ena = (_zz_ena_462[0] && sData_fire_463);
  assign mData_462 = xil_SimpleDualBram_462_doutb;
  assign xil_SimpleDualBram_463_addra = _zz_addra_463[10:0];
  assign xil_SimpleDualBram_463_addrb = _zz_addrb_463[13:0];
  assign sData_fire_464 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_463_ena = (_zz_ena_463[0] && sData_fire_464);
  assign mData_463 = xil_SimpleDualBram_463_doutb;
  assign xil_SimpleDualBram_464_addra = _zz_addra_464[10:0];
  assign xil_SimpleDualBram_464_addrb = _zz_addrb_464[13:0];
  assign sData_fire_465 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_464_ena = (_zz_ena_464[0] && sData_fire_465);
  assign mData_464 = xil_SimpleDualBram_464_doutb;
  assign xil_SimpleDualBram_465_addra = _zz_addra_465[10:0];
  assign xil_SimpleDualBram_465_addrb = _zz_addrb_465[13:0];
  assign sData_fire_466 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_465_ena = (_zz_ena_465[0] && sData_fire_466);
  assign mData_465 = xil_SimpleDualBram_465_doutb;
  assign xil_SimpleDualBram_466_addra = _zz_addra_466[10:0];
  assign xil_SimpleDualBram_466_addrb = _zz_addrb_466[13:0];
  assign sData_fire_467 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_466_ena = (_zz_ena_466[0] && sData_fire_467);
  assign mData_466 = xil_SimpleDualBram_466_doutb;
  assign xil_SimpleDualBram_467_addra = _zz_addra_467[10:0];
  assign xil_SimpleDualBram_467_addrb = _zz_addrb_467[13:0];
  assign sData_fire_468 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_467_ena = (_zz_ena_467[0] && sData_fire_468);
  assign mData_467 = xil_SimpleDualBram_467_doutb;
  assign xil_SimpleDualBram_468_addra = _zz_addra_468[10:0];
  assign xil_SimpleDualBram_468_addrb = _zz_addrb_468[13:0];
  assign sData_fire_469 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_468_ena = (_zz_ena_468[0] && sData_fire_469);
  assign mData_468 = xil_SimpleDualBram_468_doutb;
  assign xil_SimpleDualBram_469_addra = _zz_addra_469[10:0];
  assign xil_SimpleDualBram_469_addrb = _zz_addrb_469[13:0];
  assign sData_fire_470 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_469_ena = (_zz_ena_469[0] && sData_fire_470);
  assign mData_469 = xil_SimpleDualBram_469_doutb;
  assign xil_SimpleDualBram_470_addra = _zz_addra_470[10:0];
  assign xil_SimpleDualBram_470_addrb = _zz_addrb_470[13:0];
  assign sData_fire_471 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_470_ena = (_zz_ena_470[0] && sData_fire_471);
  assign mData_470 = xil_SimpleDualBram_470_doutb;
  assign xil_SimpleDualBram_471_addra = _zz_addra_471[10:0];
  assign xil_SimpleDualBram_471_addrb = _zz_addrb_471[13:0];
  assign sData_fire_472 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_471_ena = (_zz_ena_471[0] && sData_fire_472);
  assign mData_471 = xil_SimpleDualBram_471_doutb;
  assign xil_SimpleDualBram_472_addra = _zz_addra_472[10:0];
  assign xil_SimpleDualBram_472_addrb = _zz_addrb_472[13:0];
  assign sData_fire_473 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_472_ena = (_zz_ena_472[0] && sData_fire_473);
  assign mData_472 = xil_SimpleDualBram_472_doutb;
  assign xil_SimpleDualBram_473_addra = _zz_addra_473[10:0];
  assign xil_SimpleDualBram_473_addrb = _zz_addrb_473[13:0];
  assign sData_fire_474 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_473_ena = (_zz_ena_473[0] && sData_fire_474);
  assign mData_473 = xil_SimpleDualBram_473_doutb;
  assign xil_SimpleDualBram_474_addra = _zz_addra_474[10:0];
  assign xil_SimpleDualBram_474_addrb = _zz_addrb_474[13:0];
  assign sData_fire_475 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_474_ena = (_zz_ena_474[0] && sData_fire_475);
  assign mData_474 = xil_SimpleDualBram_474_doutb;
  assign xil_SimpleDualBram_475_addra = _zz_addra_475[10:0];
  assign xil_SimpleDualBram_475_addrb = _zz_addrb_475[13:0];
  assign sData_fire_476 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_475_ena = (_zz_ena_475[0] && sData_fire_476);
  assign mData_475 = xil_SimpleDualBram_475_doutb;
  assign xil_SimpleDualBram_476_addra = _zz_addra_476[10:0];
  assign xil_SimpleDualBram_476_addrb = _zz_addrb_476[13:0];
  assign sData_fire_477 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_476_ena = (_zz_ena_476[0] && sData_fire_477);
  assign mData_476 = xil_SimpleDualBram_476_doutb;
  assign xil_SimpleDualBram_477_addra = _zz_addra_477[10:0];
  assign xil_SimpleDualBram_477_addrb = _zz_addrb_477[13:0];
  assign sData_fire_478 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_477_ena = (_zz_ena_477[0] && sData_fire_478);
  assign mData_477 = xil_SimpleDualBram_477_doutb;
  assign xil_SimpleDualBram_478_addra = _zz_addra_478[10:0];
  assign xil_SimpleDualBram_478_addrb = _zz_addrb_478[13:0];
  assign sData_fire_479 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_478_ena = (_zz_ena_478[0] && sData_fire_479);
  assign mData_478 = xil_SimpleDualBram_478_doutb;
  assign xil_SimpleDualBram_479_addra = _zz_addra_479[10:0];
  assign xil_SimpleDualBram_479_addrb = _zz_addrb_479[13:0];
  assign sData_fire_480 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_479_ena = (_zz_ena_479[0] && sData_fire_480);
  assign mData_479 = xil_SimpleDualBram_479_doutb;
  assign xil_SimpleDualBram_480_addra = _zz_addra_480[10:0];
  assign xil_SimpleDualBram_480_addrb = _zz_addrb_480[13:0];
  assign sData_fire_481 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_480_ena = (_zz_ena_480[0] && sData_fire_481);
  assign mData_480 = xil_SimpleDualBram_480_doutb;
  assign xil_SimpleDualBram_481_addra = _zz_addra_481[10:0];
  assign xil_SimpleDualBram_481_addrb = _zz_addrb_481[13:0];
  assign sData_fire_482 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_481_ena = (_zz_ena_481[0] && sData_fire_482);
  assign mData_481 = xil_SimpleDualBram_481_doutb;
  assign xil_SimpleDualBram_482_addra = _zz_addra_482[10:0];
  assign xil_SimpleDualBram_482_addrb = _zz_addrb_482[13:0];
  assign sData_fire_483 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_482_ena = (_zz_ena_482[0] && sData_fire_483);
  assign mData_482 = xil_SimpleDualBram_482_doutb;
  assign xil_SimpleDualBram_483_addra = _zz_addra_483[10:0];
  assign xil_SimpleDualBram_483_addrb = _zz_addrb_483[13:0];
  assign sData_fire_484 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_483_ena = (_zz_ena_483[0] && sData_fire_484);
  assign mData_483 = xil_SimpleDualBram_483_doutb;
  assign xil_SimpleDualBram_484_addra = _zz_addra_484[10:0];
  assign xil_SimpleDualBram_484_addrb = _zz_addrb_484[13:0];
  assign sData_fire_485 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_484_ena = (_zz_ena_484[0] && sData_fire_485);
  assign mData_484 = xil_SimpleDualBram_484_doutb;
  assign xil_SimpleDualBram_485_addra = _zz_addra_485[10:0];
  assign xil_SimpleDualBram_485_addrb = _zz_addrb_485[13:0];
  assign sData_fire_486 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_485_ena = (_zz_ena_485[0] && sData_fire_486);
  assign mData_485 = xil_SimpleDualBram_485_doutb;
  assign xil_SimpleDualBram_486_addra = _zz_addra_486[10:0];
  assign xil_SimpleDualBram_486_addrb = _zz_addrb_486[13:0];
  assign sData_fire_487 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_486_ena = (_zz_ena_486[0] && sData_fire_487);
  assign mData_486 = xil_SimpleDualBram_486_doutb;
  assign xil_SimpleDualBram_487_addra = _zz_addra_487[10:0];
  assign xil_SimpleDualBram_487_addrb = _zz_addrb_487[13:0];
  assign sData_fire_488 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_487_ena = (_zz_ena_487[0] && sData_fire_488);
  assign mData_487 = xil_SimpleDualBram_487_doutb;
  assign xil_SimpleDualBram_488_addra = _zz_addra_488[10:0];
  assign xil_SimpleDualBram_488_addrb = _zz_addrb_488[13:0];
  assign sData_fire_489 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_488_ena = (_zz_ena_488[0] && sData_fire_489);
  assign mData_488 = xil_SimpleDualBram_488_doutb;
  assign xil_SimpleDualBram_489_addra = _zz_addra_489[10:0];
  assign xil_SimpleDualBram_489_addrb = _zz_addrb_489[13:0];
  assign sData_fire_490 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_489_ena = (_zz_ena_489[0] && sData_fire_490);
  assign mData_489 = xil_SimpleDualBram_489_doutb;
  assign xil_SimpleDualBram_490_addra = _zz_addra_490[10:0];
  assign xil_SimpleDualBram_490_addrb = _zz_addrb_490[13:0];
  assign sData_fire_491 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_490_ena = (_zz_ena_490[0] && sData_fire_491);
  assign mData_490 = xil_SimpleDualBram_490_doutb;
  assign xil_SimpleDualBram_491_addra = _zz_addra_491[10:0];
  assign xil_SimpleDualBram_491_addrb = _zz_addrb_491[13:0];
  assign sData_fire_492 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_491_ena = (_zz_ena_491[0] && sData_fire_492);
  assign mData_491 = xil_SimpleDualBram_491_doutb;
  assign xil_SimpleDualBram_492_addra = _zz_addra_492[10:0];
  assign xil_SimpleDualBram_492_addrb = _zz_addrb_492[13:0];
  assign sData_fire_493 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_492_ena = (_zz_ena_492[0] && sData_fire_493);
  assign mData_492 = xil_SimpleDualBram_492_doutb;
  assign xil_SimpleDualBram_493_addra = _zz_addra_493[10:0];
  assign xil_SimpleDualBram_493_addrb = _zz_addrb_493[13:0];
  assign sData_fire_494 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_493_ena = (_zz_ena_493[0] && sData_fire_494);
  assign mData_493 = xil_SimpleDualBram_493_doutb;
  assign xil_SimpleDualBram_494_addra = _zz_addra_494[10:0];
  assign xil_SimpleDualBram_494_addrb = _zz_addrb_494[13:0];
  assign sData_fire_495 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_494_ena = (_zz_ena_494[0] && sData_fire_495);
  assign mData_494 = xil_SimpleDualBram_494_doutb;
  assign xil_SimpleDualBram_495_addra = _zz_addra_495[10:0];
  assign xil_SimpleDualBram_495_addrb = _zz_addrb_495[13:0];
  assign sData_fire_496 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_495_ena = (_zz_ena_495[0] && sData_fire_496);
  assign mData_495 = xil_SimpleDualBram_495_doutb;
  assign xil_SimpleDualBram_496_addra = _zz_addra_496[10:0];
  assign xil_SimpleDualBram_496_addrb = _zz_addrb_496[13:0];
  assign sData_fire_497 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_496_ena = (_zz_ena_496[0] && sData_fire_497);
  assign mData_496 = xil_SimpleDualBram_496_doutb;
  assign xil_SimpleDualBram_497_addra = _zz_addra_497[10:0];
  assign xil_SimpleDualBram_497_addrb = _zz_addrb_497[13:0];
  assign sData_fire_498 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_497_ena = (_zz_ena_497[0] && sData_fire_498);
  assign mData_497 = xil_SimpleDualBram_497_doutb;
  assign xil_SimpleDualBram_498_addra = _zz_addra_498[10:0];
  assign xil_SimpleDualBram_498_addrb = _zz_addrb_498[13:0];
  assign sData_fire_499 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_498_ena = (_zz_ena_498[0] && sData_fire_499);
  assign mData_498 = xil_SimpleDualBram_498_doutb;
  assign xil_SimpleDualBram_499_addra = _zz_addra_499[10:0];
  assign xil_SimpleDualBram_499_addrb = _zz_addrb_499[13:0];
  assign sData_fire_500 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_499_ena = (_zz_ena_499[0] && sData_fire_500);
  assign mData_499 = xil_SimpleDualBram_499_doutb;
  assign xil_SimpleDualBram_500_addra = _zz_addra_500[10:0];
  assign xil_SimpleDualBram_500_addrb = _zz_addrb_500[13:0];
  assign sData_fire_501 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_500_ena = (_zz_ena_500[0] && sData_fire_501);
  assign mData_500 = xil_SimpleDualBram_500_doutb;
  assign xil_SimpleDualBram_501_addra = _zz_addra_501[10:0];
  assign xil_SimpleDualBram_501_addrb = _zz_addrb_501[13:0];
  assign sData_fire_502 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_501_ena = (_zz_ena_501[0] && sData_fire_502);
  assign mData_501 = xil_SimpleDualBram_501_doutb;
  assign xil_SimpleDualBram_502_addra = _zz_addra_502[10:0];
  assign xil_SimpleDualBram_502_addrb = _zz_addrb_502[13:0];
  assign sData_fire_503 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_502_ena = (_zz_ena_502[0] && sData_fire_503);
  assign mData_502 = xil_SimpleDualBram_502_doutb;
  assign xil_SimpleDualBram_503_addra = _zz_addra_503[10:0];
  assign xil_SimpleDualBram_503_addrb = _zz_addrb_503[13:0];
  assign sData_fire_504 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_503_ena = (_zz_ena_503[0] && sData_fire_504);
  assign mData_503 = xil_SimpleDualBram_503_doutb;
  assign xil_SimpleDualBram_504_addra = _zz_addra_504[10:0];
  assign xil_SimpleDualBram_504_addrb = _zz_addrb_504[13:0];
  assign sData_fire_505 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_504_ena = (_zz_ena_504[0] && sData_fire_505);
  assign mData_504 = xil_SimpleDualBram_504_doutb;
  assign xil_SimpleDualBram_505_addra = _zz_addra_505[10:0];
  assign xil_SimpleDualBram_505_addrb = _zz_addrb_505[13:0];
  assign sData_fire_506 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_505_ena = (_zz_ena_505[0] && sData_fire_506);
  assign mData_505 = xil_SimpleDualBram_505_doutb;
  assign xil_SimpleDualBram_506_addra = _zz_addra_506[10:0];
  assign xil_SimpleDualBram_506_addrb = _zz_addrb_506[13:0];
  assign sData_fire_507 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_506_ena = (_zz_ena_506[0] && sData_fire_507);
  assign mData_506 = xil_SimpleDualBram_506_doutb;
  assign xil_SimpleDualBram_507_addra = _zz_addra_507[10:0];
  assign xil_SimpleDualBram_507_addrb = _zz_addrb_507[13:0];
  assign sData_fire_508 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_507_ena = (_zz_ena_507[0] && sData_fire_508);
  assign mData_507 = xil_SimpleDualBram_507_doutb;
  assign xil_SimpleDualBram_508_addra = _zz_addra_508[10:0];
  assign xil_SimpleDualBram_508_addrb = _zz_addrb_508[13:0];
  assign sData_fire_509 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_508_ena = (_zz_ena_508[0] && sData_fire_509);
  assign mData_508 = xil_SimpleDualBram_508_doutb;
  assign xil_SimpleDualBram_509_addra = _zz_addra_509[10:0];
  assign xil_SimpleDualBram_509_addrb = _zz_addrb_509[13:0];
  assign sData_fire_510 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_509_ena = (_zz_ena_509[0] && sData_fire_510);
  assign mData_509 = xil_SimpleDualBram_509_doutb;
  assign xil_SimpleDualBram_510_addra = _zz_addra_510[10:0];
  assign xil_SimpleDualBram_510_addrb = _zz_addrb_510[13:0];
  assign sData_fire_511 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_510_ena = (_zz_ena_510[0] && sData_fire_511);
  assign mData_510 = xil_SimpleDualBram_510_doutb;
  assign xil_SimpleDualBram_511_addra = _zz_addra_511[10:0];
  assign xil_SimpleDualBram_511_addrb = _zz_addrb_511[13:0];
  assign sData_fire_512 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_511_ena = (_zz_ena_511[0] && sData_fire_512);
  assign mData_511 = xil_SimpleDualBram_511_doutb;
  assign sData_ready = ((Fsm_currentState & WEIGHT_CACHE_STATUS_CACHE_WEIGHT) != 4'b0000);
  assign Fsm_SA_Computed = LayerEnd;
  always @(*) begin
    case(OutCol_Cnt_count)
      16'h0001 : begin
        MatrixCol_Switch_1[0 : 0] = 1'b1;
        MatrixCol_Switch_1[7 : 1] = 7'h0;
      end
      16'h0002 : begin
        MatrixCol_Switch_1[1 : 0] = 2'b11;
        MatrixCol_Switch_1[7 : 2] = 6'h0;
      end
      16'h0003 : begin
        MatrixCol_Switch_1[2 : 0] = 3'b111;
        MatrixCol_Switch_1[7 : 3] = 5'h0;
      end
      16'h0004 : begin
        MatrixCol_Switch_1[3 : 0] = 4'b1111;
        MatrixCol_Switch_1[7 : 4] = 4'b0000;
      end
      16'h0005 : begin
        MatrixCol_Switch_1[4 : 0] = 5'h1f;
        MatrixCol_Switch_1[7 : 5] = 3'b000;
      end
      16'h0006 : begin
        MatrixCol_Switch_1[5 : 0] = 6'h3f;
        MatrixCol_Switch_1[7 : 6] = 2'b00;
      end
      16'h0007 : begin
        MatrixCol_Switch_1[6 : 0] = 7'h7f;
        MatrixCol_Switch_1[7 : 7] = 1'b0;
      end
      default : begin
        MatrixCol_Switch_1 = 8'hff;
      end
    endcase
  end

  assign MatrixCol_Switch = MatrixCol_Switch_1_regNext;
  always @(posedge clk) begin
    start_regNext <= start;
    MatrixCol_Switch_1_regNext <= MatrixCol_Switch_1;
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= WEIGHT_CACHE_STATUS_IDLE;
      Init_Count_count <= 3'b000;
      InData_Switch <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
      In_Row_Cnt_count <= 16'h0;
      In_Col_Cnt_count <= 16'h0;
      Read_Row_Base_Addr <= 16'h0;
      Write_Row_Base_Addr <= 16'h0;
      OutRow_Cnt_count <= 16'h0;
      OutCol_Cnt_count <= Matrix_Col;
      Col_In_8_Cnt_count <= 9'h0;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l19) begin
        Init_Count_count <= (Init_Count_count + 3'b001);
        if(Init_Count_valid) begin
          Init_Count_count <= 3'b000;
        end
      end
      if(sData_fire) begin
        if(In_Row_Cnt_valid) begin
          In_Row_Cnt_count <= 16'h0;
        end else begin
          In_Row_Cnt_count <= (In_Row_Cnt_count + 16'h0001);
        end
      end
      if(In_Row_Cnt_valid) begin
        if(In_Col_Cnt_valid) begin
          In_Col_Cnt_count <= 16'h0;
        end else begin
          In_Col_Cnt_count <= (In_Col_Cnt_count + 16'h0001);
        end
      end
      if(when_WaCounter_l40) begin
        if(OutRow_Cnt_valid) begin
          OutRow_Cnt_count <= 16'h0;
        end else begin
          OutRow_Cnt_count <= (OutRow_Cnt_count + 16'h0001);
        end
      end
      if(OutRow_Cnt_valid) begin
        if(OutCol_Cnt_valid) begin
          OutCol_Cnt_count <= Matrix_Col;
        end else begin
          OutCol_Cnt_count <= (OutCol_Cnt_count - _zz_OutCol_Cnt_count_1);
        end
      end
      if(start) begin
        OutCol_Cnt_count <= Matrix_Col;
      end
      if(In_Row_Cnt_valid) begin
        if(Col_In_8_Cnt_valid) begin
          Col_In_8_Cnt_count <= 9'h0;
        end else begin
          Col_In_8_Cnt_count <= (Col_In_8_Cnt_count + 9'h001);
        end
      end
      if(OutCol_Cnt_valid) begin
        Col_In_8_Cnt_count <= 9'h0;
        Read_Row_Base_Addr <= 16'h0;
      end else begin
        if(OutRow_Cnt_valid) begin
          Read_Row_Base_Addr <= (Read_Row_Base_Addr + Matrix_Row);
        end
      end
      if(when_SA3D_WeightCache_l129) begin
        InData_Switch <= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
      end else begin
        if(In_Row_Cnt_valid) begin
          InData_Switch <= {InData_Switch[510 : 0],InData_Switch[511 : 511]};
        end
      end
      if(when_SA3D_WeightCache_l134) begin
        Write_Row_Base_Addr <= 16'h0;
      end else begin
        if(Col_In_8_Cnt_valid) begin
          Write_Row_Base_Addr <= (Write_Row_Base_Addr + _zz_Write_Row_Base_Addr);
        end
      end
    end
  end


endmodule
