// Generator : SpinalHDL v1.7.0    git head : eca519e78d4e6022e34911ec300a432ed9db8220
// Component : Tile
// Git hash  : 3f47e2272714eaadc4903fce7d57faff55e9534d

`timescale 1ns/1ps

module Tile (
  input      [63:0]   activate,
  input      [63:0]   weight,
  input               vaild,
  input      [15:0]   signCount,
  output reg [19:0]   PE_OUT_0,
  output reg [19:0]   PE_OUT_1,
  output reg [19:0]   PE_OUT_2,
  output reg [19:0]   PE_OUT_3,
  output reg [19:0]   PE_OUT_4,
  output reg [19:0]   PE_OUT_5,
  output reg [19:0]   PE_OUT_6,
  output reg [19:0]   PE_OUT_7,
  output reg          resultVaild_0,
  output reg          resultVaild_1,
  output reg          resultVaild_2,
  output reg          resultVaild_3,
  output reg          resultVaild_4,
  output reg          resultVaild_5,
  output reg          resultVaild_6,
  output reg          resultVaild_7,
  input               clk,
  input               reset
);

  wire       [7:0]    pE_64_activate;
  wire       [7:0]    pE_64_weight;
  wire       [7:0]    pE_65_activate;
  wire       [7:0]    pE_66_activate;
  wire       [7:0]    pE_67_activate;
  wire       [7:0]    pE_68_activate;
  wire       [7:0]    pE_69_activate;
  wire       [7:0]    pE_70_activate;
  wire       [7:0]    pE_71_activate;
  wire       [7:0]    pE_64_acount;
  wire       [7:0]    pE_64_bcount;
  wire       [19:0]   pE_64_PE_OUT;
  wire                pE_64_finish;
  wire       [7:0]    pE_65_acount;
  wire       [7:0]    pE_65_bcount;
  wire       [19:0]   pE_65_PE_OUT;
  wire                pE_65_finish;
  wire       [7:0]    pE_66_acount;
  wire       [7:0]    pE_66_bcount;
  wire       [19:0]   pE_66_PE_OUT;
  wire                pE_66_finish;
  wire       [7:0]    pE_67_acount;
  wire       [7:0]    pE_67_bcount;
  wire       [19:0]   pE_67_PE_OUT;
  wire                pE_67_finish;
  wire       [7:0]    pE_68_acount;
  wire       [7:0]    pE_68_bcount;
  wire       [19:0]   pE_68_PE_OUT;
  wire                pE_68_finish;
  wire       [7:0]    pE_69_acount;
  wire       [7:0]    pE_69_bcount;
  wire       [19:0]   pE_69_PE_OUT;
  wire                pE_69_finish;
  wire       [7:0]    pE_70_acount;
  wire       [7:0]    pE_70_bcount;
  wire       [19:0]   pE_70_PE_OUT;
  wire                pE_70_finish;
  wire       [7:0]    pE_71_acount;
  wire       [7:0]    pE_71_bcount;
  wire       [19:0]   pE_71_PE_OUT;
  wire                pE_71_finish;
  wire       [7:0]    pE_72_acount;
  wire       [7:0]    pE_72_bcount;
  wire       [19:0]   pE_72_PE_OUT;
  wire                pE_72_finish;
  wire       [7:0]    pE_73_acount;
  wire       [7:0]    pE_73_bcount;
  wire       [19:0]   pE_73_PE_OUT;
  wire                pE_73_finish;
  wire       [7:0]    pE_74_acount;
  wire       [7:0]    pE_74_bcount;
  wire       [19:0]   pE_74_PE_OUT;
  wire                pE_74_finish;
  wire       [7:0]    pE_75_acount;
  wire       [7:0]    pE_75_bcount;
  wire       [19:0]   pE_75_PE_OUT;
  wire                pE_75_finish;
  wire       [7:0]    pE_76_acount;
  wire       [7:0]    pE_76_bcount;
  wire       [19:0]   pE_76_PE_OUT;
  wire                pE_76_finish;
  wire       [7:0]    pE_77_acount;
  wire       [7:0]    pE_77_bcount;
  wire       [19:0]   pE_77_PE_OUT;
  wire                pE_77_finish;
  wire       [7:0]    pE_78_acount;
  wire       [7:0]    pE_78_bcount;
  wire       [19:0]   pE_78_PE_OUT;
  wire                pE_78_finish;
  wire       [7:0]    pE_79_acount;
  wire       [7:0]    pE_79_bcount;
  wire       [19:0]   pE_79_PE_OUT;
  wire                pE_79_finish;
  wire       [7:0]    pE_80_acount;
  wire       [7:0]    pE_80_bcount;
  wire       [19:0]   pE_80_PE_OUT;
  wire                pE_80_finish;
  wire       [7:0]    pE_81_acount;
  wire       [7:0]    pE_81_bcount;
  wire       [19:0]   pE_81_PE_OUT;
  wire                pE_81_finish;
  wire       [7:0]    pE_82_acount;
  wire       [7:0]    pE_82_bcount;
  wire       [19:0]   pE_82_PE_OUT;
  wire                pE_82_finish;
  wire       [7:0]    pE_83_acount;
  wire       [7:0]    pE_83_bcount;
  wire       [19:0]   pE_83_PE_OUT;
  wire                pE_83_finish;
  wire       [7:0]    pE_84_acount;
  wire       [7:0]    pE_84_bcount;
  wire       [19:0]   pE_84_PE_OUT;
  wire                pE_84_finish;
  wire       [7:0]    pE_85_acount;
  wire       [7:0]    pE_85_bcount;
  wire       [19:0]   pE_85_PE_OUT;
  wire                pE_85_finish;
  wire       [7:0]    pE_86_acount;
  wire       [7:0]    pE_86_bcount;
  wire       [19:0]   pE_86_PE_OUT;
  wire                pE_86_finish;
  wire       [7:0]    pE_87_acount;
  wire       [7:0]    pE_87_bcount;
  wire       [19:0]   pE_87_PE_OUT;
  wire                pE_87_finish;
  wire       [7:0]    pE_88_acount;
  wire       [7:0]    pE_88_bcount;
  wire       [19:0]   pE_88_PE_OUT;
  wire                pE_88_finish;
  wire       [7:0]    pE_89_acount;
  wire       [7:0]    pE_89_bcount;
  wire       [19:0]   pE_89_PE_OUT;
  wire                pE_89_finish;
  wire       [7:0]    pE_90_acount;
  wire       [7:0]    pE_90_bcount;
  wire       [19:0]   pE_90_PE_OUT;
  wire                pE_90_finish;
  wire       [7:0]    pE_91_acount;
  wire       [7:0]    pE_91_bcount;
  wire       [19:0]   pE_91_PE_OUT;
  wire                pE_91_finish;
  wire       [7:0]    pE_92_acount;
  wire       [7:0]    pE_92_bcount;
  wire       [19:0]   pE_92_PE_OUT;
  wire                pE_92_finish;
  wire       [7:0]    pE_93_acount;
  wire       [7:0]    pE_93_bcount;
  wire       [19:0]   pE_93_PE_OUT;
  wire                pE_93_finish;
  wire       [7:0]    pE_94_acount;
  wire       [7:0]    pE_94_bcount;
  wire       [19:0]   pE_94_PE_OUT;
  wire                pE_94_finish;
  wire       [7:0]    pE_95_acount;
  wire       [7:0]    pE_95_bcount;
  wire       [19:0]   pE_95_PE_OUT;
  wire                pE_95_finish;
  wire       [7:0]    pE_96_acount;
  wire       [7:0]    pE_96_bcount;
  wire       [19:0]   pE_96_PE_OUT;
  wire                pE_96_finish;
  wire       [7:0]    pE_97_acount;
  wire       [7:0]    pE_97_bcount;
  wire       [19:0]   pE_97_PE_OUT;
  wire                pE_97_finish;
  wire       [7:0]    pE_98_acount;
  wire       [7:0]    pE_98_bcount;
  wire       [19:0]   pE_98_PE_OUT;
  wire                pE_98_finish;
  wire       [7:0]    pE_99_acount;
  wire       [7:0]    pE_99_bcount;
  wire       [19:0]   pE_99_PE_OUT;
  wire                pE_99_finish;
  wire       [7:0]    pE_100_acount;
  wire       [7:0]    pE_100_bcount;
  wire       [19:0]   pE_100_PE_OUT;
  wire                pE_100_finish;
  wire       [7:0]    pE_101_acount;
  wire       [7:0]    pE_101_bcount;
  wire       [19:0]   pE_101_PE_OUT;
  wire                pE_101_finish;
  wire       [7:0]    pE_102_acount;
  wire       [7:0]    pE_102_bcount;
  wire       [19:0]   pE_102_PE_OUT;
  wire                pE_102_finish;
  wire       [7:0]    pE_103_acount;
  wire       [7:0]    pE_103_bcount;
  wire       [19:0]   pE_103_PE_OUT;
  wire                pE_103_finish;
  wire       [7:0]    pE_104_acount;
  wire       [7:0]    pE_104_bcount;
  wire       [19:0]   pE_104_PE_OUT;
  wire                pE_104_finish;
  wire       [7:0]    pE_105_acount;
  wire       [7:0]    pE_105_bcount;
  wire       [19:0]   pE_105_PE_OUT;
  wire                pE_105_finish;
  wire       [7:0]    pE_106_acount;
  wire       [7:0]    pE_106_bcount;
  wire       [19:0]   pE_106_PE_OUT;
  wire                pE_106_finish;
  wire       [7:0]    pE_107_acount;
  wire       [7:0]    pE_107_bcount;
  wire       [19:0]   pE_107_PE_OUT;
  wire                pE_107_finish;
  wire       [7:0]    pE_108_acount;
  wire       [7:0]    pE_108_bcount;
  wire       [19:0]   pE_108_PE_OUT;
  wire                pE_108_finish;
  wire       [7:0]    pE_109_acount;
  wire       [7:0]    pE_109_bcount;
  wire       [19:0]   pE_109_PE_OUT;
  wire                pE_109_finish;
  wire       [7:0]    pE_110_acount;
  wire       [7:0]    pE_110_bcount;
  wire       [19:0]   pE_110_PE_OUT;
  wire                pE_110_finish;
  wire       [7:0]    pE_111_acount;
  wire       [7:0]    pE_111_bcount;
  wire       [19:0]   pE_111_PE_OUT;
  wire                pE_111_finish;
  wire       [7:0]    pE_112_acount;
  wire       [7:0]    pE_112_bcount;
  wire       [19:0]   pE_112_PE_OUT;
  wire                pE_112_finish;
  wire       [7:0]    pE_113_acount;
  wire       [7:0]    pE_113_bcount;
  wire       [19:0]   pE_113_PE_OUT;
  wire                pE_113_finish;
  wire       [7:0]    pE_114_acount;
  wire       [7:0]    pE_114_bcount;
  wire       [19:0]   pE_114_PE_OUT;
  wire                pE_114_finish;
  wire       [7:0]    pE_115_acount;
  wire       [7:0]    pE_115_bcount;
  wire       [19:0]   pE_115_PE_OUT;
  wire                pE_115_finish;
  wire       [7:0]    pE_116_acount;
  wire       [7:0]    pE_116_bcount;
  wire       [19:0]   pE_116_PE_OUT;
  wire                pE_116_finish;
  wire       [7:0]    pE_117_acount;
  wire       [7:0]    pE_117_bcount;
  wire       [19:0]   pE_117_PE_OUT;
  wire                pE_117_finish;
  wire       [7:0]    pE_118_acount;
  wire       [7:0]    pE_118_bcount;
  wire       [19:0]   pE_118_PE_OUT;
  wire                pE_118_finish;
  wire       [7:0]    pE_119_acount;
  wire       [7:0]    pE_119_bcount;
  wire       [19:0]   pE_119_PE_OUT;
  wire                pE_119_finish;
  wire       [7:0]    pE_120_acount;
  wire       [7:0]    pE_120_bcount;
  wire       [19:0]   pE_120_PE_OUT;
  wire                pE_120_finish;
  wire       [7:0]    pE_121_acount;
  wire       [7:0]    pE_121_bcount;
  wire       [19:0]   pE_121_PE_OUT;
  wire                pE_121_finish;
  wire       [7:0]    pE_122_acount;
  wire       [7:0]    pE_122_bcount;
  wire       [19:0]   pE_122_PE_OUT;
  wire                pE_122_finish;
  wire       [7:0]    pE_123_acount;
  wire       [7:0]    pE_123_bcount;
  wire       [19:0]   pE_123_PE_OUT;
  wire                pE_123_finish;
  wire       [7:0]    pE_124_acount;
  wire       [7:0]    pE_124_bcount;
  wire       [19:0]   pE_124_PE_OUT;
  wire                pE_124_finish;
  wire       [7:0]    pE_125_acount;
  wire       [7:0]    pE_125_bcount;
  wire       [19:0]   pE_125_PE_OUT;
  wire                pE_125_finish;
  wire       [7:0]    pE_126_acount;
  wire       [7:0]    pE_126_bcount;
  wire       [19:0]   pE_126_PE_OUT;
  wire                pE_126_finish;
  wire       [7:0]    pE_127_acount;
  wire       [7:0]    pE_127_bcount;
  wire       [19:0]   pE_127_PE_OUT;
  wire                pE_127_finish;
  reg                 vaild_delay_1;
  reg                 vaild_delay_1_1;
  reg                 vaild_delay_2;
  reg                 vaild_delay_1_2;
  reg                 vaild_delay_2_1;
  reg                 vaild_delay_3;
  reg                 vaild_delay_1_3;
  reg                 vaild_delay_2_2;
  reg                 vaild_delay_3_1;
  reg                 vaild_delay_4;
  reg                 vaild_delay_1_4;
  reg                 vaild_delay_2_3;
  reg                 vaild_delay_3_2;
  reg                 vaild_delay_4_1;
  reg                 vaild_delay_5;
  reg                 vaild_delay_1_5;
  reg                 vaild_delay_2_4;
  reg                 vaild_delay_3_3;
  reg                 vaild_delay_4_2;
  reg                 vaild_delay_5_1;
  reg                 vaild_delay_6;
  reg                 vaild_delay_1_6;
  reg                 vaild_delay_2_5;
  reg                 vaild_delay_3_4;
  reg                 vaild_delay_4_3;
  reg                 vaild_delay_5_2;
  reg                 vaild_delay_6_1;
  reg                 vaild_delay_7;
  reg        [7:0]    _zz_weight;
  reg                 vaild_delay_1_7;
  reg        [7:0]    _zz_weight_1;
  reg        [7:0]    _zz_weight_2;
  reg                 vaild_delay_1_8;
  reg                 vaild_delay_2_6;
  reg        [7:0]    _zz_weight_3;
  reg        [7:0]    _zz_weight_4;
  reg        [7:0]    _zz_weight_5;
  reg                 vaild_delay_1_9;
  reg                 vaild_delay_2_7;
  reg                 vaild_delay_3_5;
  reg        [7:0]    _zz_weight_6;
  reg        [7:0]    _zz_weight_7;
  reg        [7:0]    _zz_weight_8;
  reg        [7:0]    _zz_weight_9;
  reg                 vaild_delay_1_10;
  reg                 vaild_delay_2_8;
  reg                 vaild_delay_3_6;
  reg                 vaild_delay_4_4;
  reg        [7:0]    _zz_weight_10;
  reg        [7:0]    _zz_weight_11;
  reg        [7:0]    _zz_weight_12;
  reg        [7:0]    _zz_weight_13;
  reg        [7:0]    _zz_weight_14;
  reg                 vaild_delay_1_11;
  reg                 vaild_delay_2_9;
  reg                 vaild_delay_3_7;
  reg                 vaild_delay_4_5;
  reg                 vaild_delay_5_3;
  reg        [7:0]    _zz_weight_15;
  reg        [7:0]    _zz_weight_16;
  reg        [7:0]    _zz_weight_17;
  reg        [7:0]    _zz_weight_18;
  reg        [7:0]    _zz_weight_19;
  reg        [7:0]    _zz_weight_20;
  reg                 vaild_delay_1_12;
  reg                 vaild_delay_2_10;
  reg                 vaild_delay_3_8;
  reg                 vaild_delay_4_6;
  reg                 vaild_delay_5_4;
  reg                 vaild_delay_6_2;
  reg        [7:0]    _zz_weight_21;
  reg        [7:0]    _zz_weight_22;
  reg        [7:0]    _zz_weight_23;
  reg        [7:0]    _zz_weight_24;
  reg        [7:0]    _zz_weight_25;
  reg        [7:0]    _zz_weight_26;
  reg        [7:0]    _zz_weight_27;
  reg                 vaild_delay_1_13;
  reg                 vaild_delay_2_11;
  reg                 vaild_delay_3_9;
  reg                 vaild_delay_4_7;
  reg                 vaild_delay_5_5;
  reg                 vaild_delay_6_3;
  reg                 vaild_delay_7_1;
  reg                 pE_65_vaild_delay_1;
  reg                 pE_79_vaild_delay_1;
  reg                 pE_80_vaild_delay_1;
  reg                 pE_81_vaild_delay_1;
  reg                 pE_82_vaild_delay_1;
  reg                 pE_83_vaild_delay_1;
  reg                 pE_84_vaild_delay_1;
  reg                 pE_66_vaild_delay_1;
  reg                 pE_86_vaild_delay_1;
  reg                 pE_87_vaild_delay_1;
  reg                 pE_88_vaild_delay_1;
  reg                 pE_89_vaild_delay_1;
  reg                 pE_90_vaild_delay_1;
  reg                 pE_91_vaild_delay_1;
  reg                 pE_67_vaild_delay_1;
  reg                 pE_93_vaild_delay_1;
  reg                 pE_94_vaild_delay_1;
  reg                 pE_95_vaild_delay_1;
  reg                 pE_96_vaild_delay_1;
  reg                 pE_97_vaild_delay_1;
  reg                 pE_98_vaild_delay_1;
  reg                 pE_68_vaild_delay_1;
  reg                 pE_100_vaild_delay_1;
  reg                 pE_101_vaild_delay_1;
  reg                 pE_102_vaild_delay_1;
  reg                 pE_103_vaild_delay_1;
  reg                 pE_104_vaild_delay_1;
  reg                 pE_105_vaild_delay_1;
  reg                 pE_69_vaild_delay_1;
  reg                 pE_107_vaild_delay_1;
  reg                 pE_108_vaild_delay_1;
  reg                 pE_109_vaild_delay_1;
  reg                 pE_110_vaild_delay_1;
  reg                 pE_111_vaild_delay_1;
  reg                 pE_112_vaild_delay_1;
  reg                 pE_70_vaild_delay_1;
  reg                 pE_114_vaild_delay_1;
  reg                 pE_115_vaild_delay_1;
  reg                 pE_116_vaild_delay_1;
  reg                 pE_117_vaild_delay_1;
  reg                 pE_118_vaild_delay_1;
  reg                 pE_119_vaild_delay_1;
  reg                 pE_71_vaild_delay_1;
  reg                 pE_121_vaild_delay_1;
  reg                 pE_122_vaild_delay_1;
  reg                 pE_123_vaild_delay_1;
  reg                 pE_124_vaild_delay_1;
  reg                 pE_125_vaild_delay_1;
  reg                 pE_126_vaild_delay_1;
  wire                when_Tile_l68;
  wire                when_Tile_l68_1;
  wire                when_Tile_l68_2;
  wire                when_Tile_l68_3;
  wire                when_Tile_l68_4;
  wire                when_Tile_l68_5;
  wire                when_Tile_l68_6;
  wire                when_Tile_l68_7;
  wire                when_Tile_l68_8;
  wire                when_Tile_l68_9;
  wire                when_Tile_l68_10;
  wire                when_Tile_l68_11;
  wire                when_Tile_l68_12;
  wire                when_Tile_l68_13;
  wire                when_Tile_l68_14;
  wire                when_Tile_l68_15;
  wire                when_Tile_l68_16;
  wire                when_Tile_l68_17;
  wire                when_Tile_l68_18;
  wire                when_Tile_l68_19;
  wire                when_Tile_l68_20;
  wire                when_Tile_l68_21;
  wire                when_Tile_l68_22;
  wire                when_Tile_l68_23;
  wire                when_Tile_l68_24;
  wire                when_Tile_l68_25;
  wire                when_Tile_l68_26;
  wire                when_Tile_l68_27;
  wire                when_Tile_l68_28;
  wire                when_Tile_l68_29;
  wire                when_Tile_l68_30;
  wire                when_Tile_l68_31;
  wire                when_Tile_l68_32;
  wire                when_Tile_l68_33;
  wire                when_Tile_l68_34;
  wire                when_Tile_l68_35;
  wire                when_Tile_l68_36;
  wire                when_Tile_l68_37;
  wire                when_Tile_l68_38;
  wire                when_Tile_l68_39;
  wire                when_Tile_l68_40;
  wire                when_Tile_l68_41;
  wire                when_Tile_l68_42;
  wire                when_Tile_l68_43;
  wire                when_Tile_l68_44;
  wire                when_Tile_l68_45;
  wire                when_Tile_l68_46;
  wire                when_Tile_l68_47;
  wire                when_Tile_l68_48;
  wire                when_Tile_l68_49;
  wire                when_Tile_l68_50;
  wire                when_Tile_l68_51;
  wire                when_Tile_l68_52;
  wire                when_Tile_l68_53;
  wire                when_Tile_l68_54;
  wire                when_Tile_l68_55;
  wire                when_Tile_l68_56;
  wire                when_Tile_l68_57;
  wire                when_Tile_l68_58;
  wire                when_Tile_l68_59;
  wire                when_Tile_l68_60;
  wire                when_Tile_l68_61;
  wire                when_Tile_l68_62;
  wire                when_Tile_l68_63;

  PE pE_64 (
    .activate  (pE_64_activate[7:0]), //i
    .weight    (pE_64_weight[7:0]  ), //i
    .vaild     (vaild              ), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_64_acount[7:0]  ), //o
    .bcount    (pE_64_bcount[7:0]  ), //o
    .PE_OUT    (pE_64_PE_OUT[19:0] ), //o
    .finish    (pE_64_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_65 (
    .activate  (pE_65_activate[7:0]), //i
    .weight    (pE_64_bcount[7:0]  ), //i
    .vaild     (vaild_delay_1      ), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_65_acount[7:0]  ), //o
    .bcount    (pE_65_bcount[7:0]  ), //o
    .PE_OUT    (pE_65_PE_OUT[19:0] ), //o
    .finish    (pE_65_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_66 (
    .activate  (pE_66_activate[7:0]), //i
    .weight    (pE_65_bcount[7:0]  ), //i
    .vaild     (vaild_delay_2      ), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_66_acount[7:0]  ), //o
    .bcount    (pE_66_bcount[7:0]  ), //o
    .PE_OUT    (pE_66_PE_OUT[19:0] ), //o
    .finish    (pE_66_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_67 (
    .activate  (pE_67_activate[7:0]), //i
    .weight    (pE_66_bcount[7:0]  ), //i
    .vaild     (vaild_delay_3      ), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_67_acount[7:0]  ), //o
    .bcount    (pE_67_bcount[7:0]  ), //o
    .PE_OUT    (pE_67_PE_OUT[19:0] ), //o
    .finish    (pE_67_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_68 (
    .activate  (pE_68_activate[7:0]), //i
    .weight    (pE_67_bcount[7:0]  ), //i
    .vaild     (vaild_delay_4      ), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_68_acount[7:0]  ), //o
    .bcount    (pE_68_bcount[7:0]  ), //o
    .PE_OUT    (pE_68_PE_OUT[19:0] ), //o
    .finish    (pE_68_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_69 (
    .activate  (pE_69_activate[7:0]), //i
    .weight    (pE_68_bcount[7:0]  ), //i
    .vaild     (vaild_delay_5      ), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_69_acount[7:0]  ), //o
    .bcount    (pE_69_bcount[7:0]  ), //o
    .PE_OUT    (pE_69_PE_OUT[19:0] ), //o
    .finish    (pE_69_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_70 (
    .activate  (pE_70_activate[7:0]), //i
    .weight    (pE_69_bcount[7:0]  ), //i
    .vaild     (vaild_delay_6      ), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_70_acount[7:0]  ), //o
    .bcount    (pE_70_bcount[7:0]  ), //o
    .PE_OUT    (pE_70_PE_OUT[19:0] ), //o
    .finish    (pE_70_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_71 (
    .activate  (pE_71_activate[7:0]), //i
    .weight    (pE_70_bcount[7:0]  ), //i
    .vaild     (vaild_delay_7      ), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_71_acount[7:0]  ), //o
    .bcount    (pE_71_bcount[7:0]  ), //o
    .PE_OUT    (pE_71_PE_OUT[19:0] ), //o
    .finish    (pE_71_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_72 (
    .activate  (pE_64_acount[7:0] ), //i
    .weight    (_zz_weight[7:0]   ), //i
    .vaild     (vaild_delay_1_7   ), //i
    .signCount (signCount[15:0]   ), //i
    .acount    (pE_72_acount[7:0] ), //o
    .bcount    (pE_72_bcount[7:0] ), //o
    .PE_OUT    (pE_72_PE_OUT[19:0]), //o
    .finish    (pE_72_finish      ), //o
    .clk       (clk               ), //i
    .reset     (reset             )  //i
  );
  PE pE_73 (
    .activate  (pE_72_acount[7:0] ), //i
    .weight    (_zz_weight_2[7:0] ), //i
    .vaild     (vaild_delay_2_6   ), //i
    .signCount (signCount[15:0]   ), //i
    .acount    (pE_73_acount[7:0] ), //o
    .bcount    (pE_73_bcount[7:0] ), //o
    .PE_OUT    (pE_73_PE_OUT[19:0]), //o
    .finish    (pE_73_finish      ), //o
    .clk       (clk               ), //i
    .reset     (reset             )  //i
  );
  PE pE_74 (
    .activate  (pE_73_acount[7:0] ), //i
    .weight    (_zz_weight_5[7:0] ), //i
    .vaild     (vaild_delay_3_5   ), //i
    .signCount (signCount[15:0]   ), //i
    .acount    (pE_74_acount[7:0] ), //o
    .bcount    (pE_74_bcount[7:0] ), //o
    .PE_OUT    (pE_74_PE_OUT[19:0]), //o
    .finish    (pE_74_finish      ), //o
    .clk       (clk               ), //i
    .reset     (reset             )  //i
  );
  PE pE_75 (
    .activate  (pE_74_acount[7:0] ), //i
    .weight    (_zz_weight_9[7:0] ), //i
    .vaild     (vaild_delay_4_4   ), //i
    .signCount (signCount[15:0]   ), //i
    .acount    (pE_75_acount[7:0] ), //o
    .bcount    (pE_75_bcount[7:0] ), //o
    .PE_OUT    (pE_75_PE_OUT[19:0]), //o
    .finish    (pE_75_finish      ), //o
    .clk       (clk               ), //i
    .reset     (reset             )  //i
  );
  PE pE_76 (
    .activate  (pE_75_acount[7:0] ), //i
    .weight    (_zz_weight_14[7:0]), //i
    .vaild     (vaild_delay_5_3   ), //i
    .signCount (signCount[15:0]   ), //i
    .acount    (pE_76_acount[7:0] ), //o
    .bcount    (pE_76_bcount[7:0] ), //o
    .PE_OUT    (pE_76_PE_OUT[19:0]), //o
    .finish    (pE_76_finish      ), //o
    .clk       (clk               ), //i
    .reset     (reset             )  //i
  );
  PE pE_77 (
    .activate  (pE_76_acount[7:0] ), //i
    .weight    (_zz_weight_20[7:0]), //i
    .vaild     (vaild_delay_6_2   ), //i
    .signCount (signCount[15:0]   ), //i
    .acount    (pE_77_acount[7:0] ), //o
    .bcount    (pE_77_bcount[7:0] ), //o
    .PE_OUT    (pE_77_PE_OUT[19:0]), //o
    .finish    (pE_77_finish      ), //o
    .clk       (clk               ), //i
    .reset     (reset             )  //i
  );
  PE pE_78 (
    .activate  (pE_77_acount[7:0] ), //i
    .weight    (_zz_weight_27[7:0]), //i
    .vaild     (vaild_delay_7_1   ), //i
    .signCount (signCount[15:0]   ), //i
    .acount    (pE_78_acount[7:0] ), //o
    .bcount    (pE_78_bcount[7:0] ), //o
    .PE_OUT    (pE_78_PE_OUT[19:0]), //o
    .finish    (pE_78_finish      ), //o
    .clk       (clk               ), //i
    .reset     (reset             )  //i
  );
  PE pE_79 (
    .activate  (pE_65_acount[7:0]  ), //i
    .weight    (pE_72_bcount[7:0]  ), //i
    .vaild     (pE_65_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_79_acount[7:0]  ), //o
    .bcount    (pE_79_bcount[7:0]  ), //o
    .PE_OUT    (pE_79_PE_OUT[19:0] ), //o
    .finish    (pE_79_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_80 (
    .activate  (pE_79_acount[7:0]  ), //i
    .weight    (pE_73_bcount[7:0]  ), //i
    .vaild     (pE_79_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_80_acount[7:0]  ), //o
    .bcount    (pE_80_bcount[7:0]  ), //o
    .PE_OUT    (pE_80_PE_OUT[19:0] ), //o
    .finish    (pE_80_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_81 (
    .activate  (pE_80_acount[7:0]  ), //i
    .weight    (pE_74_bcount[7:0]  ), //i
    .vaild     (pE_80_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_81_acount[7:0]  ), //o
    .bcount    (pE_81_bcount[7:0]  ), //o
    .PE_OUT    (pE_81_PE_OUT[19:0] ), //o
    .finish    (pE_81_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_82 (
    .activate  (pE_81_acount[7:0]  ), //i
    .weight    (pE_75_bcount[7:0]  ), //i
    .vaild     (pE_81_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_82_acount[7:0]  ), //o
    .bcount    (pE_82_bcount[7:0]  ), //o
    .PE_OUT    (pE_82_PE_OUT[19:0] ), //o
    .finish    (pE_82_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_83 (
    .activate  (pE_82_acount[7:0]  ), //i
    .weight    (pE_76_bcount[7:0]  ), //i
    .vaild     (pE_82_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_83_acount[7:0]  ), //o
    .bcount    (pE_83_bcount[7:0]  ), //o
    .PE_OUT    (pE_83_PE_OUT[19:0] ), //o
    .finish    (pE_83_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_84 (
    .activate  (pE_83_acount[7:0]  ), //i
    .weight    (pE_77_bcount[7:0]  ), //i
    .vaild     (pE_83_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_84_acount[7:0]  ), //o
    .bcount    (pE_84_bcount[7:0]  ), //o
    .PE_OUT    (pE_84_PE_OUT[19:0] ), //o
    .finish    (pE_84_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_85 (
    .activate  (pE_84_acount[7:0]  ), //i
    .weight    (pE_78_bcount[7:0]  ), //i
    .vaild     (pE_84_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_85_acount[7:0]  ), //o
    .bcount    (pE_85_bcount[7:0]  ), //o
    .PE_OUT    (pE_85_PE_OUT[19:0] ), //o
    .finish    (pE_85_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_86 (
    .activate  (pE_66_acount[7:0]  ), //i
    .weight    (pE_79_bcount[7:0]  ), //i
    .vaild     (pE_66_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_86_acount[7:0]  ), //o
    .bcount    (pE_86_bcount[7:0]  ), //o
    .PE_OUT    (pE_86_PE_OUT[19:0] ), //o
    .finish    (pE_86_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_87 (
    .activate  (pE_86_acount[7:0]  ), //i
    .weight    (pE_80_bcount[7:0]  ), //i
    .vaild     (pE_86_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_87_acount[7:0]  ), //o
    .bcount    (pE_87_bcount[7:0]  ), //o
    .PE_OUT    (pE_87_PE_OUT[19:0] ), //o
    .finish    (pE_87_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_88 (
    .activate  (pE_87_acount[7:0]  ), //i
    .weight    (pE_81_bcount[7:0]  ), //i
    .vaild     (pE_87_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_88_acount[7:0]  ), //o
    .bcount    (pE_88_bcount[7:0]  ), //o
    .PE_OUT    (pE_88_PE_OUT[19:0] ), //o
    .finish    (pE_88_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_89 (
    .activate  (pE_88_acount[7:0]  ), //i
    .weight    (pE_82_bcount[7:0]  ), //i
    .vaild     (pE_88_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_89_acount[7:0]  ), //o
    .bcount    (pE_89_bcount[7:0]  ), //o
    .PE_OUT    (pE_89_PE_OUT[19:0] ), //o
    .finish    (pE_89_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_90 (
    .activate  (pE_89_acount[7:0]  ), //i
    .weight    (pE_83_bcount[7:0]  ), //i
    .vaild     (pE_89_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_90_acount[7:0]  ), //o
    .bcount    (pE_90_bcount[7:0]  ), //o
    .PE_OUT    (pE_90_PE_OUT[19:0] ), //o
    .finish    (pE_90_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_91 (
    .activate  (pE_90_acount[7:0]  ), //i
    .weight    (pE_84_bcount[7:0]  ), //i
    .vaild     (pE_90_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_91_acount[7:0]  ), //o
    .bcount    (pE_91_bcount[7:0]  ), //o
    .PE_OUT    (pE_91_PE_OUT[19:0] ), //o
    .finish    (pE_91_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_92 (
    .activate  (pE_91_acount[7:0]  ), //i
    .weight    (pE_85_bcount[7:0]  ), //i
    .vaild     (pE_91_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_92_acount[7:0]  ), //o
    .bcount    (pE_92_bcount[7:0]  ), //o
    .PE_OUT    (pE_92_PE_OUT[19:0] ), //o
    .finish    (pE_92_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_93 (
    .activate  (pE_67_acount[7:0]  ), //i
    .weight    (pE_86_bcount[7:0]  ), //i
    .vaild     (pE_67_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_93_acount[7:0]  ), //o
    .bcount    (pE_93_bcount[7:0]  ), //o
    .PE_OUT    (pE_93_PE_OUT[19:0] ), //o
    .finish    (pE_93_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_94 (
    .activate  (pE_93_acount[7:0]  ), //i
    .weight    (pE_87_bcount[7:0]  ), //i
    .vaild     (pE_93_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_94_acount[7:0]  ), //o
    .bcount    (pE_94_bcount[7:0]  ), //o
    .PE_OUT    (pE_94_PE_OUT[19:0] ), //o
    .finish    (pE_94_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_95 (
    .activate  (pE_94_acount[7:0]  ), //i
    .weight    (pE_88_bcount[7:0]  ), //i
    .vaild     (pE_94_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_95_acount[7:0]  ), //o
    .bcount    (pE_95_bcount[7:0]  ), //o
    .PE_OUT    (pE_95_PE_OUT[19:0] ), //o
    .finish    (pE_95_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_96 (
    .activate  (pE_95_acount[7:0]  ), //i
    .weight    (pE_89_bcount[7:0]  ), //i
    .vaild     (pE_95_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_96_acount[7:0]  ), //o
    .bcount    (pE_96_bcount[7:0]  ), //o
    .PE_OUT    (pE_96_PE_OUT[19:0] ), //o
    .finish    (pE_96_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_97 (
    .activate  (pE_96_acount[7:0]  ), //i
    .weight    (pE_90_bcount[7:0]  ), //i
    .vaild     (pE_96_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_97_acount[7:0]  ), //o
    .bcount    (pE_97_bcount[7:0]  ), //o
    .PE_OUT    (pE_97_PE_OUT[19:0] ), //o
    .finish    (pE_97_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_98 (
    .activate  (pE_97_acount[7:0]  ), //i
    .weight    (pE_91_bcount[7:0]  ), //i
    .vaild     (pE_97_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_98_acount[7:0]  ), //o
    .bcount    (pE_98_bcount[7:0]  ), //o
    .PE_OUT    (pE_98_PE_OUT[19:0] ), //o
    .finish    (pE_98_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_99 (
    .activate  (pE_98_acount[7:0]  ), //i
    .weight    (pE_92_bcount[7:0]  ), //i
    .vaild     (pE_98_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_99_acount[7:0]  ), //o
    .bcount    (pE_99_bcount[7:0]  ), //o
    .PE_OUT    (pE_99_PE_OUT[19:0] ), //o
    .finish    (pE_99_finish       ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_100 (
    .activate  (pE_68_acount[7:0]  ), //i
    .weight    (pE_93_bcount[7:0]  ), //i
    .vaild     (pE_68_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_100_acount[7:0] ), //o
    .bcount    (pE_100_bcount[7:0] ), //o
    .PE_OUT    (pE_100_PE_OUT[19:0]), //o
    .finish    (pE_100_finish      ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_101 (
    .activate  (pE_100_acount[7:0]  ), //i
    .weight    (pE_94_bcount[7:0]   ), //i
    .vaild     (pE_100_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_101_acount[7:0]  ), //o
    .bcount    (pE_101_bcount[7:0]  ), //o
    .PE_OUT    (pE_101_PE_OUT[19:0] ), //o
    .finish    (pE_101_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_102 (
    .activate  (pE_101_acount[7:0]  ), //i
    .weight    (pE_95_bcount[7:0]   ), //i
    .vaild     (pE_101_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_102_acount[7:0]  ), //o
    .bcount    (pE_102_bcount[7:0]  ), //o
    .PE_OUT    (pE_102_PE_OUT[19:0] ), //o
    .finish    (pE_102_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_103 (
    .activate  (pE_102_acount[7:0]  ), //i
    .weight    (pE_96_bcount[7:0]   ), //i
    .vaild     (pE_102_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_103_acount[7:0]  ), //o
    .bcount    (pE_103_bcount[7:0]  ), //o
    .PE_OUT    (pE_103_PE_OUT[19:0] ), //o
    .finish    (pE_103_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_104 (
    .activate  (pE_103_acount[7:0]  ), //i
    .weight    (pE_97_bcount[7:0]   ), //i
    .vaild     (pE_103_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_104_acount[7:0]  ), //o
    .bcount    (pE_104_bcount[7:0]  ), //o
    .PE_OUT    (pE_104_PE_OUT[19:0] ), //o
    .finish    (pE_104_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_105 (
    .activate  (pE_104_acount[7:0]  ), //i
    .weight    (pE_98_bcount[7:0]   ), //i
    .vaild     (pE_104_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_105_acount[7:0]  ), //o
    .bcount    (pE_105_bcount[7:0]  ), //o
    .PE_OUT    (pE_105_PE_OUT[19:0] ), //o
    .finish    (pE_105_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_106 (
    .activate  (pE_105_acount[7:0]  ), //i
    .weight    (pE_99_bcount[7:0]   ), //i
    .vaild     (pE_105_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_106_acount[7:0]  ), //o
    .bcount    (pE_106_bcount[7:0]  ), //o
    .PE_OUT    (pE_106_PE_OUT[19:0] ), //o
    .finish    (pE_106_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_107 (
    .activate  (pE_69_acount[7:0]  ), //i
    .weight    (pE_100_bcount[7:0] ), //i
    .vaild     (pE_69_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_107_acount[7:0] ), //o
    .bcount    (pE_107_bcount[7:0] ), //o
    .PE_OUT    (pE_107_PE_OUT[19:0]), //o
    .finish    (pE_107_finish      ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_108 (
    .activate  (pE_107_acount[7:0]  ), //i
    .weight    (pE_101_bcount[7:0]  ), //i
    .vaild     (pE_107_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_108_acount[7:0]  ), //o
    .bcount    (pE_108_bcount[7:0]  ), //o
    .PE_OUT    (pE_108_PE_OUT[19:0] ), //o
    .finish    (pE_108_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_109 (
    .activate  (pE_108_acount[7:0]  ), //i
    .weight    (pE_102_bcount[7:0]  ), //i
    .vaild     (pE_108_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_109_acount[7:0]  ), //o
    .bcount    (pE_109_bcount[7:0]  ), //o
    .PE_OUT    (pE_109_PE_OUT[19:0] ), //o
    .finish    (pE_109_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_110 (
    .activate  (pE_109_acount[7:0]  ), //i
    .weight    (pE_103_bcount[7:0]  ), //i
    .vaild     (pE_109_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_110_acount[7:0]  ), //o
    .bcount    (pE_110_bcount[7:0]  ), //o
    .PE_OUT    (pE_110_PE_OUT[19:0] ), //o
    .finish    (pE_110_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_111 (
    .activate  (pE_110_acount[7:0]  ), //i
    .weight    (pE_104_bcount[7:0]  ), //i
    .vaild     (pE_110_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_111_acount[7:0]  ), //o
    .bcount    (pE_111_bcount[7:0]  ), //o
    .PE_OUT    (pE_111_PE_OUT[19:0] ), //o
    .finish    (pE_111_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_112 (
    .activate  (pE_111_acount[7:0]  ), //i
    .weight    (pE_105_bcount[7:0]  ), //i
    .vaild     (pE_111_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_112_acount[7:0]  ), //o
    .bcount    (pE_112_bcount[7:0]  ), //o
    .PE_OUT    (pE_112_PE_OUT[19:0] ), //o
    .finish    (pE_112_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_113 (
    .activate  (pE_112_acount[7:0]  ), //i
    .weight    (pE_106_bcount[7:0]  ), //i
    .vaild     (pE_112_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_113_acount[7:0]  ), //o
    .bcount    (pE_113_bcount[7:0]  ), //o
    .PE_OUT    (pE_113_PE_OUT[19:0] ), //o
    .finish    (pE_113_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_114 (
    .activate  (pE_70_acount[7:0]  ), //i
    .weight    (pE_107_bcount[7:0] ), //i
    .vaild     (pE_70_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_114_acount[7:0] ), //o
    .bcount    (pE_114_bcount[7:0] ), //o
    .PE_OUT    (pE_114_PE_OUT[19:0]), //o
    .finish    (pE_114_finish      ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_115 (
    .activate  (pE_114_acount[7:0]  ), //i
    .weight    (pE_108_bcount[7:0]  ), //i
    .vaild     (pE_114_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_115_acount[7:0]  ), //o
    .bcount    (pE_115_bcount[7:0]  ), //o
    .PE_OUT    (pE_115_PE_OUT[19:0] ), //o
    .finish    (pE_115_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_116 (
    .activate  (pE_115_acount[7:0]  ), //i
    .weight    (pE_109_bcount[7:0]  ), //i
    .vaild     (pE_115_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_116_acount[7:0]  ), //o
    .bcount    (pE_116_bcount[7:0]  ), //o
    .PE_OUT    (pE_116_PE_OUT[19:0] ), //o
    .finish    (pE_116_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_117 (
    .activate  (pE_116_acount[7:0]  ), //i
    .weight    (pE_110_bcount[7:0]  ), //i
    .vaild     (pE_116_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_117_acount[7:0]  ), //o
    .bcount    (pE_117_bcount[7:0]  ), //o
    .PE_OUT    (pE_117_PE_OUT[19:0] ), //o
    .finish    (pE_117_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_118 (
    .activate  (pE_117_acount[7:0]  ), //i
    .weight    (pE_111_bcount[7:0]  ), //i
    .vaild     (pE_117_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_118_acount[7:0]  ), //o
    .bcount    (pE_118_bcount[7:0]  ), //o
    .PE_OUT    (pE_118_PE_OUT[19:0] ), //o
    .finish    (pE_118_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_119 (
    .activate  (pE_118_acount[7:0]  ), //i
    .weight    (pE_112_bcount[7:0]  ), //i
    .vaild     (pE_118_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_119_acount[7:0]  ), //o
    .bcount    (pE_119_bcount[7:0]  ), //o
    .PE_OUT    (pE_119_PE_OUT[19:0] ), //o
    .finish    (pE_119_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_120 (
    .activate  (pE_119_acount[7:0]  ), //i
    .weight    (pE_113_bcount[7:0]  ), //i
    .vaild     (pE_119_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_120_acount[7:0]  ), //o
    .bcount    (pE_120_bcount[7:0]  ), //o
    .PE_OUT    (pE_120_PE_OUT[19:0] ), //o
    .finish    (pE_120_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_121 (
    .activate  (pE_71_acount[7:0]  ), //i
    .weight    (pE_114_bcount[7:0] ), //i
    .vaild     (pE_71_vaild_delay_1), //i
    .signCount (signCount[15:0]    ), //i
    .acount    (pE_121_acount[7:0] ), //o
    .bcount    (pE_121_bcount[7:0] ), //o
    .PE_OUT    (pE_121_PE_OUT[19:0]), //o
    .finish    (pE_121_finish      ), //o
    .clk       (clk                ), //i
    .reset     (reset              )  //i
  );
  PE pE_122 (
    .activate  (pE_121_acount[7:0]  ), //i
    .weight    (pE_115_bcount[7:0]  ), //i
    .vaild     (pE_121_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_122_acount[7:0]  ), //o
    .bcount    (pE_122_bcount[7:0]  ), //o
    .PE_OUT    (pE_122_PE_OUT[19:0] ), //o
    .finish    (pE_122_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_123 (
    .activate  (pE_122_acount[7:0]  ), //i
    .weight    (pE_116_bcount[7:0]  ), //i
    .vaild     (pE_122_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_123_acount[7:0]  ), //o
    .bcount    (pE_123_bcount[7:0]  ), //o
    .PE_OUT    (pE_123_PE_OUT[19:0] ), //o
    .finish    (pE_123_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_124 (
    .activate  (pE_123_acount[7:0]  ), //i
    .weight    (pE_117_bcount[7:0]  ), //i
    .vaild     (pE_123_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_124_acount[7:0]  ), //o
    .bcount    (pE_124_bcount[7:0]  ), //o
    .PE_OUT    (pE_124_PE_OUT[19:0] ), //o
    .finish    (pE_124_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_125 (
    .activate  (pE_124_acount[7:0]  ), //i
    .weight    (pE_118_bcount[7:0]  ), //i
    .vaild     (pE_124_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_125_acount[7:0]  ), //o
    .bcount    (pE_125_bcount[7:0]  ), //o
    .PE_OUT    (pE_125_PE_OUT[19:0] ), //o
    .finish    (pE_125_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_126 (
    .activate  (pE_125_acount[7:0]  ), //i
    .weight    (pE_119_bcount[7:0]  ), //i
    .vaild     (pE_125_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_126_acount[7:0]  ), //o
    .bcount    (pE_126_bcount[7:0]  ), //o
    .PE_OUT    (pE_126_PE_OUT[19:0] ), //o
    .finish    (pE_126_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  PE pE_127 (
    .activate  (pE_126_acount[7:0]  ), //i
    .weight    (pE_120_bcount[7:0]  ), //i
    .vaild     (pE_126_vaild_delay_1), //i
    .signCount (signCount[15:0]     ), //i
    .acount    (pE_127_acount[7:0]  ), //o
    .bcount    (pE_127_bcount[7:0]  ), //o
    .PE_OUT    (pE_127_PE_OUT[19:0] ), //o
    .finish    (pE_127_finish       ), //o
    .clk       (clk                 ), //i
    .reset     (reset               )  //i
  );
  always @(*) begin
    PE_OUT_0 = 20'h0;
    if(when_Tile_l68) begin
      PE_OUT_0 = pE_64_PE_OUT;
    end
    if(when_Tile_l68_1) begin
      PE_OUT_0 = pE_72_PE_OUT;
    end
    if(when_Tile_l68_2) begin
      PE_OUT_0 = pE_73_PE_OUT;
    end
    if(when_Tile_l68_3) begin
      PE_OUT_0 = pE_74_PE_OUT;
    end
    if(when_Tile_l68_4) begin
      PE_OUT_0 = pE_75_PE_OUT;
    end
    if(when_Tile_l68_5) begin
      PE_OUT_0 = pE_76_PE_OUT;
    end
    if(when_Tile_l68_6) begin
      PE_OUT_0 = pE_77_PE_OUT;
    end
    if(when_Tile_l68_7) begin
      PE_OUT_0 = pE_78_PE_OUT;
    end
  end

  always @(*) begin
    resultVaild_0 = 1'b0;
    if(when_Tile_l68) begin
      resultVaild_0 = pE_64_finish;
    end
    if(when_Tile_l68_1) begin
      resultVaild_0 = pE_72_finish;
    end
    if(when_Tile_l68_2) begin
      resultVaild_0 = pE_73_finish;
    end
    if(when_Tile_l68_3) begin
      resultVaild_0 = pE_74_finish;
    end
    if(when_Tile_l68_4) begin
      resultVaild_0 = pE_75_finish;
    end
    if(when_Tile_l68_5) begin
      resultVaild_0 = pE_76_finish;
    end
    if(when_Tile_l68_6) begin
      resultVaild_0 = pE_77_finish;
    end
    if(when_Tile_l68_7) begin
      resultVaild_0 = pE_78_finish;
    end
  end

  always @(*) begin
    PE_OUT_1 = 20'h0;
    if(when_Tile_l68_8) begin
      PE_OUT_1 = pE_65_PE_OUT;
    end
    if(when_Tile_l68_9) begin
      PE_OUT_1 = pE_79_PE_OUT;
    end
    if(when_Tile_l68_10) begin
      PE_OUT_1 = pE_80_PE_OUT;
    end
    if(when_Tile_l68_11) begin
      PE_OUT_1 = pE_81_PE_OUT;
    end
    if(when_Tile_l68_12) begin
      PE_OUT_1 = pE_82_PE_OUT;
    end
    if(when_Tile_l68_13) begin
      PE_OUT_1 = pE_83_PE_OUT;
    end
    if(when_Tile_l68_14) begin
      PE_OUT_1 = pE_84_PE_OUT;
    end
    if(when_Tile_l68_15) begin
      PE_OUT_1 = pE_85_PE_OUT;
    end
  end

  always @(*) begin
    resultVaild_1 = 1'b0;
    if(when_Tile_l68_8) begin
      resultVaild_1 = pE_65_finish;
    end
    if(when_Tile_l68_9) begin
      resultVaild_1 = pE_79_finish;
    end
    if(when_Tile_l68_10) begin
      resultVaild_1 = pE_80_finish;
    end
    if(when_Tile_l68_11) begin
      resultVaild_1 = pE_81_finish;
    end
    if(when_Tile_l68_12) begin
      resultVaild_1 = pE_82_finish;
    end
    if(when_Tile_l68_13) begin
      resultVaild_1 = pE_83_finish;
    end
    if(when_Tile_l68_14) begin
      resultVaild_1 = pE_84_finish;
    end
    if(when_Tile_l68_15) begin
      resultVaild_1 = pE_85_finish;
    end
  end

  always @(*) begin
    PE_OUT_2 = 20'h0;
    if(when_Tile_l68_16) begin
      PE_OUT_2 = pE_66_PE_OUT;
    end
    if(when_Tile_l68_17) begin
      PE_OUT_2 = pE_86_PE_OUT;
    end
    if(when_Tile_l68_18) begin
      PE_OUT_2 = pE_87_PE_OUT;
    end
    if(when_Tile_l68_19) begin
      PE_OUT_2 = pE_88_PE_OUT;
    end
    if(when_Tile_l68_20) begin
      PE_OUT_2 = pE_89_PE_OUT;
    end
    if(when_Tile_l68_21) begin
      PE_OUT_2 = pE_90_PE_OUT;
    end
    if(when_Tile_l68_22) begin
      PE_OUT_2 = pE_91_PE_OUT;
    end
    if(when_Tile_l68_23) begin
      PE_OUT_2 = pE_92_PE_OUT;
    end
  end

  always @(*) begin
    resultVaild_2 = 1'b0;
    if(when_Tile_l68_16) begin
      resultVaild_2 = pE_66_finish;
    end
    if(when_Tile_l68_17) begin
      resultVaild_2 = pE_86_finish;
    end
    if(when_Tile_l68_18) begin
      resultVaild_2 = pE_87_finish;
    end
    if(when_Tile_l68_19) begin
      resultVaild_2 = pE_88_finish;
    end
    if(when_Tile_l68_20) begin
      resultVaild_2 = pE_89_finish;
    end
    if(when_Tile_l68_21) begin
      resultVaild_2 = pE_90_finish;
    end
    if(when_Tile_l68_22) begin
      resultVaild_2 = pE_91_finish;
    end
    if(when_Tile_l68_23) begin
      resultVaild_2 = pE_92_finish;
    end
  end

  always @(*) begin
    PE_OUT_3 = 20'h0;
    if(when_Tile_l68_24) begin
      PE_OUT_3 = pE_67_PE_OUT;
    end
    if(when_Tile_l68_25) begin
      PE_OUT_3 = pE_93_PE_OUT;
    end
    if(when_Tile_l68_26) begin
      PE_OUT_3 = pE_94_PE_OUT;
    end
    if(when_Tile_l68_27) begin
      PE_OUT_3 = pE_95_PE_OUT;
    end
    if(when_Tile_l68_28) begin
      PE_OUT_3 = pE_96_PE_OUT;
    end
    if(when_Tile_l68_29) begin
      PE_OUT_3 = pE_97_PE_OUT;
    end
    if(when_Tile_l68_30) begin
      PE_OUT_3 = pE_98_PE_OUT;
    end
    if(when_Tile_l68_31) begin
      PE_OUT_3 = pE_99_PE_OUT;
    end
  end

  always @(*) begin
    resultVaild_3 = 1'b0;
    if(when_Tile_l68_24) begin
      resultVaild_3 = pE_67_finish;
    end
    if(when_Tile_l68_25) begin
      resultVaild_3 = pE_93_finish;
    end
    if(when_Tile_l68_26) begin
      resultVaild_3 = pE_94_finish;
    end
    if(when_Tile_l68_27) begin
      resultVaild_3 = pE_95_finish;
    end
    if(when_Tile_l68_28) begin
      resultVaild_3 = pE_96_finish;
    end
    if(when_Tile_l68_29) begin
      resultVaild_3 = pE_97_finish;
    end
    if(when_Tile_l68_30) begin
      resultVaild_3 = pE_98_finish;
    end
    if(when_Tile_l68_31) begin
      resultVaild_3 = pE_99_finish;
    end
  end

  always @(*) begin
    PE_OUT_4 = 20'h0;
    if(when_Tile_l68_32) begin
      PE_OUT_4 = pE_68_PE_OUT;
    end
    if(when_Tile_l68_33) begin
      PE_OUT_4 = pE_100_PE_OUT;
    end
    if(when_Tile_l68_34) begin
      PE_OUT_4 = pE_101_PE_OUT;
    end
    if(when_Tile_l68_35) begin
      PE_OUT_4 = pE_102_PE_OUT;
    end
    if(when_Tile_l68_36) begin
      PE_OUT_4 = pE_103_PE_OUT;
    end
    if(when_Tile_l68_37) begin
      PE_OUT_4 = pE_104_PE_OUT;
    end
    if(when_Tile_l68_38) begin
      PE_OUT_4 = pE_105_PE_OUT;
    end
    if(when_Tile_l68_39) begin
      PE_OUT_4 = pE_106_PE_OUT;
    end
  end

  always @(*) begin
    resultVaild_4 = 1'b0;
    if(when_Tile_l68_32) begin
      resultVaild_4 = pE_68_finish;
    end
    if(when_Tile_l68_33) begin
      resultVaild_4 = pE_100_finish;
    end
    if(when_Tile_l68_34) begin
      resultVaild_4 = pE_101_finish;
    end
    if(when_Tile_l68_35) begin
      resultVaild_4 = pE_102_finish;
    end
    if(when_Tile_l68_36) begin
      resultVaild_4 = pE_103_finish;
    end
    if(when_Tile_l68_37) begin
      resultVaild_4 = pE_104_finish;
    end
    if(when_Tile_l68_38) begin
      resultVaild_4 = pE_105_finish;
    end
    if(when_Tile_l68_39) begin
      resultVaild_4 = pE_106_finish;
    end
  end

  always @(*) begin
    PE_OUT_5 = 20'h0;
    if(when_Tile_l68_40) begin
      PE_OUT_5 = pE_69_PE_OUT;
    end
    if(when_Tile_l68_41) begin
      PE_OUT_5 = pE_107_PE_OUT;
    end
    if(when_Tile_l68_42) begin
      PE_OUT_5 = pE_108_PE_OUT;
    end
    if(when_Tile_l68_43) begin
      PE_OUT_5 = pE_109_PE_OUT;
    end
    if(when_Tile_l68_44) begin
      PE_OUT_5 = pE_110_PE_OUT;
    end
    if(when_Tile_l68_45) begin
      PE_OUT_5 = pE_111_PE_OUT;
    end
    if(when_Tile_l68_46) begin
      PE_OUT_5 = pE_112_PE_OUT;
    end
    if(when_Tile_l68_47) begin
      PE_OUT_5 = pE_113_PE_OUT;
    end
  end

  always @(*) begin
    resultVaild_5 = 1'b0;
    if(when_Tile_l68_40) begin
      resultVaild_5 = pE_69_finish;
    end
    if(when_Tile_l68_41) begin
      resultVaild_5 = pE_107_finish;
    end
    if(when_Tile_l68_42) begin
      resultVaild_5 = pE_108_finish;
    end
    if(when_Tile_l68_43) begin
      resultVaild_5 = pE_109_finish;
    end
    if(when_Tile_l68_44) begin
      resultVaild_5 = pE_110_finish;
    end
    if(when_Tile_l68_45) begin
      resultVaild_5 = pE_111_finish;
    end
    if(when_Tile_l68_46) begin
      resultVaild_5 = pE_112_finish;
    end
    if(when_Tile_l68_47) begin
      resultVaild_5 = pE_113_finish;
    end
  end

  always @(*) begin
    PE_OUT_6 = 20'h0;
    if(when_Tile_l68_48) begin
      PE_OUT_6 = pE_70_PE_OUT;
    end
    if(when_Tile_l68_49) begin
      PE_OUT_6 = pE_114_PE_OUT;
    end
    if(when_Tile_l68_50) begin
      PE_OUT_6 = pE_115_PE_OUT;
    end
    if(when_Tile_l68_51) begin
      PE_OUT_6 = pE_116_PE_OUT;
    end
    if(when_Tile_l68_52) begin
      PE_OUT_6 = pE_117_PE_OUT;
    end
    if(when_Tile_l68_53) begin
      PE_OUT_6 = pE_118_PE_OUT;
    end
    if(when_Tile_l68_54) begin
      PE_OUT_6 = pE_119_PE_OUT;
    end
    if(when_Tile_l68_55) begin
      PE_OUT_6 = pE_120_PE_OUT;
    end
  end

  always @(*) begin
    resultVaild_6 = 1'b0;
    if(when_Tile_l68_48) begin
      resultVaild_6 = pE_70_finish;
    end
    if(when_Tile_l68_49) begin
      resultVaild_6 = pE_114_finish;
    end
    if(when_Tile_l68_50) begin
      resultVaild_6 = pE_115_finish;
    end
    if(when_Tile_l68_51) begin
      resultVaild_6 = pE_116_finish;
    end
    if(when_Tile_l68_52) begin
      resultVaild_6 = pE_117_finish;
    end
    if(when_Tile_l68_53) begin
      resultVaild_6 = pE_118_finish;
    end
    if(when_Tile_l68_54) begin
      resultVaild_6 = pE_119_finish;
    end
    if(when_Tile_l68_55) begin
      resultVaild_6 = pE_120_finish;
    end
  end

  always @(*) begin
    PE_OUT_7 = 20'h0;
    if(when_Tile_l68_56) begin
      PE_OUT_7 = pE_71_PE_OUT;
    end
    if(when_Tile_l68_57) begin
      PE_OUT_7 = pE_121_PE_OUT;
    end
    if(when_Tile_l68_58) begin
      PE_OUT_7 = pE_122_PE_OUT;
    end
    if(when_Tile_l68_59) begin
      PE_OUT_7 = pE_123_PE_OUT;
    end
    if(when_Tile_l68_60) begin
      PE_OUT_7 = pE_124_PE_OUT;
    end
    if(when_Tile_l68_61) begin
      PE_OUT_7 = pE_125_PE_OUT;
    end
    if(when_Tile_l68_62) begin
      PE_OUT_7 = pE_126_PE_OUT;
    end
    if(when_Tile_l68_63) begin
      PE_OUT_7 = pE_127_PE_OUT;
    end
  end

  always @(*) begin
    resultVaild_7 = 1'b0;
    if(when_Tile_l68_56) begin
      resultVaild_7 = pE_71_finish;
    end
    if(when_Tile_l68_57) begin
      resultVaild_7 = pE_121_finish;
    end
    if(when_Tile_l68_58) begin
      resultVaild_7 = pE_122_finish;
    end
    if(when_Tile_l68_59) begin
      resultVaild_7 = pE_123_finish;
    end
    if(when_Tile_l68_60) begin
      resultVaild_7 = pE_124_finish;
    end
    if(when_Tile_l68_61) begin
      resultVaild_7 = pE_125_finish;
    end
    if(when_Tile_l68_62) begin
      resultVaild_7 = pE_126_finish;
    end
    if(when_Tile_l68_63) begin
      resultVaild_7 = pE_127_finish;
    end
  end

  assign pE_64_weight = weight[7 : 0];
  assign pE_64_activate = activate[7 : 0];
  assign pE_65_activate = activate[15 : 8];
  assign pE_66_activate = activate[23 : 16];
  assign pE_67_activate = activate[31 : 24];
  assign pE_68_activate = activate[39 : 32];
  assign pE_69_activate = activate[47 : 40];
  assign pE_70_activate = activate[55 : 48];
  assign pE_71_activate = activate[63 : 56];
  assign when_Tile_l68 = (pE_64_finish == 1'b1);
  assign when_Tile_l68_1 = (pE_72_finish == 1'b1);
  assign when_Tile_l68_2 = (pE_73_finish == 1'b1);
  assign when_Tile_l68_3 = (pE_74_finish == 1'b1);
  assign when_Tile_l68_4 = (pE_75_finish == 1'b1);
  assign when_Tile_l68_5 = (pE_76_finish == 1'b1);
  assign when_Tile_l68_6 = (pE_77_finish == 1'b1);
  assign when_Tile_l68_7 = (pE_78_finish == 1'b1);
  assign when_Tile_l68_8 = (pE_65_finish == 1'b1);
  assign when_Tile_l68_9 = (pE_79_finish == 1'b1);
  assign when_Tile_l68_10 = (pE_80_finish == 1'b1);
  assign when_Tile_l68_11 = (pE_81_finish == 1'b1);
  assign when_Tile_l68_12 = (pE_82_finish == 1'b1);
  assign when_Tile_l68_13 = (pE_83_finish == 1'b1);
  assign when_Tile_l68_14 = (pE_84_finish == 1'b1);
  assign when_Tile_l68_15 = (pE_85_finish == 1'b1);
  assign when_Tile_l68_16 = (pE_66_finish == 1'b1);
  assign when_Tile_l68_17 = (pE_86_finish == 1'b1);
  assign when_Tile_l68_18 = (pE_87_finish == 1'b1);
  assign when_Tile_l68_19 = (pE_88_finish == 1'b1);
  assign when_Tile_l68_20 = (pE_89_finish == 1'b1);
  assign when_Tile_l68_21 = (pE_90_finish == 1'b1);
  assign when_Tile_l68_22 = (pE_91_finish == 1'b1);
  assign when_Tile_l68_23 = (pE_92_finish == 1'b1);
  assign when_Tile_l68_24 = (pE_67_finish == 1'b1);
  assign when_Tile_l68_25 = (pE_93_finish == 1'b1);
  assign when_Tile_l68_26 = (pE_94_finish == 1'b1);
  assign when_Tile_l68_27 = (pE_95_finish == 1'b1);
  assign when_Tile_l68_28 = (pE_96_finish == 1'b1);
  assign when_Tile_l68_29 = (pE_97_finish == 1'b1);
  assign when_Tile_l68_30 = (pE_98_finish == 1'b1);
  assign when_Tile_l68_31 = (pE_99_finish == 1'b1);
  assign when_Tile_l68_32 = (pE_68_finish == 1'b1);
  assign when_Tile_l68_33 = (pE_100_finish == 1'b1);
  assign when_Tile_l68_34 = (pE_101_finish == 1'b1);
  assign when_Tile_l68_35 = (pE_102_finish == 1'b1);
  assign when_Tile_l68_36 = (pE_103_finish == 1'b1);
  assign when_Tile_l68_37 = (pE_104_finish == 1'b1);
  assign when_Tile_l68_38 = (pE_105_finish == 1'b1);
  assign when_Tile_l68_39 = (pE_106_finish == 1'b1);
  assign when_Tile_l68_40 = (pE_69_finish == 1'b1);
  assign when_Tile_l68_41 = (pE_107_finish == 1'b1);
  assign when_Tile_l68_42 = (pE_108_finish == 1'b1);
  assign when_Tile_l68_43 = (pE_109_finish == 1'b1);
  assign when_Tile_l68_44 = (pE_110_finish == 1'b1);
  assign when_Tile_l68_45 = (pE_111_finish == 1'b1);
  assign when_Tile_l68_46 = (pE_112_finish == 1'b1);
  assign when_Tile_l68_47 = (pE_113_finish == 1'b1);
  assign when_Tile_l68_48 = (pE_70_finish == 1'b1);
  assign when_Tile_l68_49 = (pE_114_finish == 1'b1);
  assign when_Tile_l68_50 = (pE_115_finish == 1'b1);
  assign when_Tile_l68_51 = (pE_116_finish == 1'b1);
  assign when_Tile_l68_52 = (pE_117_finish == 1'b1);
  assign when_Tile_l68_53 = (pE_118_finish == 1'b1);
  assign when_Tile_l68_54 = (pE_119_finish == 1'b1);
  assign when_Tile_l68_55 = (pE_120_finish == 1'b1);
  assign when_Tile_l68_56 = (pE_71_finish == 1'b1);
  assign when_Tile_l68_57 = (pE_121_finish == 1'b1);
  assign when_Tile_l68_58 = (pE_122_finish == 1'b1);
  assign when_Tile_l68_59 = (pE_123_finish == 1'b1);
  assign when_Tile_l68_60 = (pE_124_finish == 1'b1);
  assign when_Tile_l68_61 = (pE_125_finish == 1'b1);
  assign when_Tile_l68_62 = (pE_126_finish == 1'b1);
  assign when_Tile_l68_63 = (pE_127_finish == 1'b1);
  always @(posedge clk) begin
    vaild_delay_1 <= vaild;
    vaild_delay_1_1 <= vaild;
    vaild_delay_2 <= vaild_delay_1_1;
    vaild_delay_1_2 <= vaild;
    vaild_delay_2_1 <= vaild_delay_1_2;
    vaild_delay_3 <= vaild_delay_2_1;
    vaild_delay_1_3 <= vaild;
    vaild_delay_2_2 <= vaild_delay_1_3;
    vaild_delay_3_1 <= vaild_delay_2_2;
    vaild_delay_4 <= vaild_delay_3_1;
    vaild_delay_1_4 <= vaild;
    vaild_delay_2_3 <= vaild_delay_1_4;
    vaild_delay_3_2 <= vaild_delay_2_3;
    vaild_delay_4_1 <= vaild_delay_3_2;
    vaild_delay_5 <= vaild_delay_4_1;
    vaild_delay_1_5 <= vaild;
    vaild_delay_2_4 <= vaild_delay_1_5;
    vaild_delay_3_3 <= vaild_delay_2_4;
    vaild_delay_4_2 <= vaild_delay_3_3;
    vaild_delay_5_1 <= vaild_delay_4_2;
    vaild_delay_6 <= vaild_delay_5_1;
    vaild_delay_1_6 <= vaild;
    vaild_delay_2_5 <= vaild_delay_1_6;
    vaild_delay_3_4 <= vaild_delay_2_5;
    vaild_delay_4_3 <= vaild_delay_3_4;
    vaild_delay_5_2 <= vaild_delay_4_3;
    vaild_delay_6_1 <= vaild_delay_5_2;
    vaild_delay_7 <= vaild_delay_6_1;
    _zz_weight <= weight[15 : 8];
    vaild_delay_1_7 <= vaild;
    _zz_weight_1 <= weight[23 : 16];
    _zz_weight_2 <= _zz_weight_1;
    vaild_delay_1_8 <= vaild;
    vaild_delay_2_6 <= vaild_delay_1_8;
    _zz_weight_3 <= weight[31 : 24];
    _zz_weight_4 <= _zz_weight_3;
    _zz_weight_5 <= _zz_weight_4;
    vaild_delay_1_9 <= vaild;
    vaild_delay_2_7 <= vaild_delay_1_9;
    vaild_delay_3_5 <= vaild_delay_2_7;
    _zz_weight_6 <= weight[39 : 32];
    _zz_weight_7 <= _zz_weight_6;
    _zz_weight_8 <= _zz_weight_7;
    _zz_weight_9 <= _zz_weight_8;
    vaild_delay_1_10 <= vaild;
    vaild_delay_2_8 <= vaild_delay_1_10;
    vaild_delay_3_6 <= vaild_delay_2_8;
    vaild_delay_4_4 <= vaild_delay_3_6;
    _zz_weight_10 <= weight[47 : 40];
    _zz_weight_11 <= _zz_weight_10;
    _zz_weight_12 <= _zz_weight_11;
    _zz_weight_13 <= _zz_weight_12;
    _zz_weight_14 <= _zz_weight_13;
    vaild_delay_1_11 <= vaild;
    vaild_delay_2_9 <= vaild_delay_1_11;
    vaild_delay_3_7 <= vaild_delay_2_9;
    vaild_delay_4_5 <= vaild_delay_3_7;
    vaild_delay_5_3 <= vaild_delay_4_5;
    _zz_weight_15 <= weight[55 : 48];
    _zz_weight_16 <= _zz_weight_15;
    _zz_weight_17 <= _zz_weight_16;
    _zz_weight_18 <= _zz_weight_17;
    _zz_weight_19 <= _zz_weight_18;
    _zz_weight_20 <= _zz_weight_19;
    vaild_delay_1_12 <= vaild;
    vaild_delay_2_10 <= vaild_delay_1_12;
    vaild_delay_3_8 <= vaild_delay_2_10;
    vaild_delay_4_6 <= vaild_delay_3_8;
    vaild_delay_5_4 <= vaild_delay_4_6;
    vaild_delay_6_2 <= vaild_delay_5_4;
    _zz_weight_21 <= weight[63 : 56];
    _zz_weight_22 <= _zz_weight_21;
    _zz_weight_23 <= _zz_weight_22;
    _zz_weight_24 <= _zz_weight_23;
    _zz_weight_25 <= _zz_weight_24;
    _zz_weight_26 <= _zz_weight_25;
    _zz_weight_27 <= _zz_weight_26;
    vaild_delay_1_13 <= vaild;
    vaild_delay_2_11 <= vaild_delay_1_13;
    vaild_delay_3_9 <= vaild_delay_2_11;
    vaild_delay_4_7 <= vaild_delay_3_9;
    vaild_delay_5_5 <= vaild_delay_4_7;
    vaild_delay_6_3 <= vaild_delay_5_5;
    vaild_delay_7_1 <= vaild_delay_6_3;
    pE_65_vaild_delay_1 <= vaild_delay_1;
    pE_79_vaild_delay_1 <= pE_65_vaild_delay_1;
    pE_80_vaild_delay_1 <= pE_79_vaild_delay_1;
    pE_81_vaild_delay_1 <= pE_80_vaild_delay_1;
    pE_82_vaild_delay_1 <= pE_81_vaild_delay_1;
    pE_83_vaild_delay_1 <= pE_82_vaild_delay_1;
    pE_84_vaild_delay_1 <= pE_83_vaild_delay_1;
    pE_66_vaild_delay_1 <= vaild_delay_2;
    pE_86_vaild_delay_1 <= pE_66_vaild_delay_1;
    pE_87_vaild_delay_1 <= pE_86_vaild_delay_1;
    pE_88_vaild_delay_1 <= pE_87_vaild_delay_1;
    pE_89_vaild_delay_1 <= pE_88_vaild_delay_1;
    pE_90_vaild_delay_1 <= pE_89_vaild_delay_1;
    pE_91_vaild_delay_1 <= pE_90_vaild_delay_1;
    pE_67_vaild_delay_1 <= vaild_delay_3;
    pE_93_vaild_delay_1 <= pE_67_vaild_delay_1;
    pE_94_vaild_delay_1 <= pE_93_vaild_delay_1;
    pE_95_vaild_delay_1 <= pE_94_vaild_delay_1;
    pE_96_vaild_delay_1 <= pE_95_vaild_delay_1;
    pE_97_vaild_delay_1 <= pE_96_vaild_delay_1;
    pE_98_vaild_delay_1 <= pE_97_vaild_delay_1;
    pE_68_vaild_delay_1 <= vaild_delay_4;
    pE_100_vaild_delay_1 <= pE_68_vaild_delay_1;
    pE_101_vaild_delay_1 <= pE_100_vaild_delay_1;
    pE_102_vaild_delay_1 <= pE_101_vaild_delay_1;
    pE_103_vaild_delay_1 <= pE_102_vaild_delay_1;
    pE_104_vaild_delay_1 <= pE_103_vaild_delay_1;
    pE_105_vaild_delay_1 <= pE_104_vaild_delay_1;
    pE_69_vaild_delay_1 <= vaild_delay_5;
    pE_107_vaild_delay_1 <= pE_69_vaild_delay_1;
    pE_108_vaild_delay_1 <= pE_107_vaild_delay_1;
    pE_109_vaild_delay_1 <= pE_108_vaild_delay_1;
    pE_110_vaild_delay_1 <= pE_109_vaild_delay_1;
    pE_111_vaild_delay_1 <= pE_110_vaild_delay_1;
    pE_112_vaild_delay_1 <= pE_111_vaild_delay_1;
    pE_70_vaild_delay_1 <= vaild_delay_6;
    pE_114_vaild_delay_1 <= pE_70_vaild_delay_1;
    pE_115_vaild_delay_1 <= pE_114_vaild_delay_1;
    pE_116_vaild_delay_1 <= pE_115_vaild_delay_1;
    pE_117_vaild_delay_1 <= pE_116_vaild_delay_1;
    pE_118_vaild_delay_1 <= pE_117_vaild_delay_1;
    pE_119_vaild_delay_1 <= pE_118_vaild_delay_1;
    pE_71_vaild_delay_1 <= vaild_delay_7;
    pE_121_vaild_delay_1 <= pE_71_vaild_delay_1;
    pE_122_vaild_delay_1 <= pE_121_vaild_delay_1;
    pE_123_vaild_delay_1 <= pE_122_vaild_delay_1;
    pE_124_vaild_delay_1 <= pE_123_vaild_delay_1;
    pE_125_vaild_delay_1 <= pE_124_vaild_delay_1;
    pE_126_vaild_delay_1 <= pE_125_vaild_delay_1;
  end


endmodule

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

//PE replaced by PE

module PE (
  input      [7:0]    activate,
  input      [7:0]    weight,
  input               vaild,
  input      [15:0]   signCount,
  output     [7:0]    acount,
  output     [7:0]    bcount,
  output reg [19:0]   PE_OUT,
  output              finish,
  input               clk,
  input               reset
);

  wire       [15:0]   dsp_P;
  wire       [19:0]   _zz_reg1;
  reg        [19:0]   reg1;
  reg                 vaild_regNext;
  reg                 vaild_regNext_1;
  reg                 vaild_regNext_1_regNext;
  reg        [15:0]   finishCnt_count;
  reg                 finishCnt_valid;
  wire                when_WaCounter_l13;
  reg        [7:0]    activate_regNext;
  reg        [7:0]    weight_regNext;

  assign _zz_reg1 = {4'd0, dsp_P};
  dsp_marco dsp (
    .CLK (clk          ), //i
    .A   (activate[7:0]), //i
    .B   (weight[7:0]  ), //i
    .P   (dsp_P[15:0]  )  //o
  );
  assign when_WaCounter_l13 = (finishCnt_count == signCount);
  always @(*) begin
    if(when_WaCounter_l13) begin
      finishCnt_valid = 1'b1;
    end else begin
      finishCnt_valid = 1'b0;
    end
  end

  assign finish = finishCnt_valid;
  always @(*) begin
    if(finishCnt_valid) begin
      PE_OUT = reg1;
    end else begin
      PE_OUT = 20'h0;
    end
  end

  assign acount = activate_regNext;
  assign bcount = weight_regNext;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      reg1 <= 20'h0;
      finishCnt_count <= 16'h0;
    end else begin
      if(vaild_regNext) begin
        reg1 <= (_zz_reg1 + reg1);
      end
      if(vaild_regNext_1_regNext) begin
        finishCnt_count <= (finishCnt_count + 16'h0001);
        if(finishCnt_valid) begin
          finishCnt_count <= 16'h0;
        end
      end
      if(finishCnt_valid) begin
        reg1 <= {4'b0000,dsp_P};
      end
    end
  end

  always @(posedge clk) begin
    vaild_regNext <= vaild;
    vaild_regNext_1 <= vaild;
    vaild_regNext_1_regNext <= vaild_regNext_1;
    activate_regNext <= activate;
    weight_regNext <= weight;
  end


endmodule
