// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : Weight_Cache
// Git hash  : 3ff479e98fb57df10a7ff9265112a692f55de7c4

`timescale 1ns/1ps

module Weight_Cache (
  input               start,
  input               sData_valid,
  output              sData_ready,
  input      [63:0]   sData_payload,
  input      [15:0]   Matrix_Row,
  input      [15:0]   Matrix_Col,
  output     [7:0]    mData_0,
  output     [7:0]    mData_1,
  output     [7:0]    mData_2,
  output     [7:0]    mData_3,
  output     [7:0]    mData_4,
  output     [7:0]    mData_5,
  output     [7:0]    mData_6,
  output     [7:0]    mData_7,
  output     [7:0]    mData_8,
  output     [7:0]    mData_9,
  output     [7:0]    mData_10,
  output     [7:0]    mData_11,
  output     [7:0]    mData_12,
  output     [7:0]    mData_13,
  output     [7:0]    mData_14,
  output     [7:0]    mData_15,
  output     [7:0]    mData_16,
  output     [7:0]    mData_17,
  output     [7:0]    mData_18,
  output     [7:0]    mData_19,
  output     [7:0]    mData_20,
  output     [7:0]    mData_21,
  output     [7:0]    mData_22,
  output     [7:0]    mData_23,
  output     [7:0]    mData_24,
  output     [7:0]    mData_25,
  output     [7:0]    mData_26,
  output     [7:0]    mData_27,
  output     [7:0]    mData_28,
  output     [7:0]    mData_29,
  output     [7:0]    mData_30,
  output     [7:0]    mData_31,
  output     [7:0]    mData_32,
  output     [7:0]    mData_33,
  output     [7:0]    mData_34,
  output     [7:0]    mData_35,
  output     [7:0]    mData_36,
  output     [7:0]    mData_37,
  output     [7:0]    mData_38,
  output     [7:0]    mData_39,
  output     [7:0]    mData_40,
  output     [7:0]    mData_41,
  output     [7:0]    mData_42,
  output     [7:0]    mData_43,
  output     [7:0]    mData_44,
  output     [7:0]    mData_45,
  output     [7:0]    mData_46,
  output     [7:0]    mData_47,
  output     [7:0]    mData_48,
  output     [7:0]    mData_49,
  output     [7:0]    mData_50,
  output     [7:0]    mData_51,
  output     [7:0]    mData_52,
  output     [7:0]    mData_53,
  output     [7:0]    mData_54,
  output     [7:0]    mData_55,
  output     [7:0]    mData_56,
  output     [7:0]    mData_57,
  output     [7:0]    mData_58,
  output     [7:0]    mData_59,
  output     [7:0]    mData_60,
  output     [7:0]    mData_61,
  output     [7:0]    mData_62,
  output     [7:0]    mData_63,
  input               Raddr_Valid,
  output              Weight_Cached,
  input               LayerEnd,
  output     [7:0]    MatrixCol_Switch,
  input               clk,
  input               reset
);
  localparam WEIGHT_CACHE_STATUS_IDLE = 4'd1;
  localparam WEIGHT_CACHE_STATUS_INIT = 4'd2;
  localparam WEIGHT_CACHE_STATUS_CACHE_WEIGHT = 4'd4;
  localparam WEIGHT_CACHE_STATUS_SA_COMPUTE = 4'd8;

  wire       [10:0]   xil_SimpleDualBram_addra;
  wire                xil_SimpleDualBram_ena;
  wire       [13:0]   xil_SimpleDualBram_addrb;
  wire       [10:0]   xil_SimpleDualBram_1_addra;
  wire                xil_SimpleDualBram_1_ena;
  wire       [13:0]   xil_SimpleDualBram_1_addrb;
  wire       [10:0]   xil_SimpleDualBram_2_addra;
  wire                xil_SimpleDualBram_2_ena;
  wire       [13:0]   xil_SimpleDualBram_2_addrb;
  wire       [10:0]   xil_SimpleDualBram_3_addra;
  wire                xil_SimpleDualBram_3_ena;
  wire       [13:0]   xil_SimpleDualBram_3_addrb;
  wire       [10:0]   xil_SimpleDualBram_4_addra;
  wire                xil_SimpleDualBram_4_ena;
  wire       [13:0]   xil_SimpleDualBram_4_addrb;
  wire       [10:0]   xil_SimpleDualBram_5_addra;
  wire                xil_SimpleDualBram_5_ena;
  wire       [13:0]   xil_SimpleDualBram_5_addrb;
  wire       [10:0]   xil_SimpleDualBram_6_addra;
  wire                xil_SimpleDualBram_6_ena;
  wire       [13:0]   xil_SimpleDualBram_6_addrb;
  wire       [10:0]   xil_SimpleDualBram_7_addra;
  wire                xil_SimpleDualBram_7_ena;
  wire       [13:0]   xil_SimpleDualBram_7_addrb;
  wire       [10:0]   xil_SimpleDualBram_8_addra;
  wire                xil_SimpleDualBram_8_ena;
  wire       [13:0]   xil_SimpleDualBram_8_addrb;
  wire       [10:0]   xil_SimpleDualBram_9_addra;
  wire                xil_SimpleDualBram_9_ena;
  wire       [13:0]   xil_SimpleDualBram_9_addrb;
  wire       [10:0]   xil_SimpleDualBram_10_addra;
  wire                xil_SimpleDualBram_10_ena;
  wire       [13:0]   xil_SimpleDualBram_10_addrb;
  wire       [10:0]   xil_SimpleDualBram_11_addra;
  wire                xil_SimpleDualBram_11_ena;
  wire       [13:0]   xil_SimpleDualBram_11_addrb;
  wire       [10:0]   xil_SimpleDualBram_12_addra;
  wire                xil_SimpleDualBram_12_ena;
  wire       [13:0]   xil_SimpleDualBram_12_addrb;
  wire       [10:0]   xil_SimpleDualBram_13_addra;
  wire                xil_SimpleDualBram_13_ena;
  wire       [13:0]   xil_SimpleDualBram_13_addrb;
  wire       [10:0]   xil_SimpleDualBram_14_addra;
  wire                xil_SimpleDualBram_14_ena;
  wire       [13:0]   xil_SimpleDualBram_14_addrb;
  wire       [10:0]   xil_SimpleDualBram_15_addra;
  wire                xil_SimpleDualBram_15_ena;
  wire       [13:0]   xil_SimpleDualBram_15_addrb;
  wire       [10:0]   xil_SimpleDualBram_16_addra;
  wire                xil_SimpleDualBram_16_ena;
  wire       [13:0]   xil_SimpleDualBram_16_addrb;
  wire       [10:0]   xil_SimpleDualBram_17_addra;
  wire                xil_SimpleDualBram_17_ena;
  wire       [13:0]   xil_SimpleDualBram_17_addrb;
  wire       [10:0]   xil_SimpleDualBram_18_addra;
  wire                xil_SimpleDualBram_18_ena;
  wire       [13:0]   xil_SimpleDualBram_18_addrb;
  wire       [10:0]   xil_SimpleDualBram_19_addra;
  wire                xil_SimpleDualBram_19_ena;
  wire       [13:0]   xil_SimpleDualBram_19_addrb;
  wire       [10:0]   xil_SimpleDualBram_20_addra;
  wire                xil_SimpleDualBram_20_ena;
  wire       [13:0]   xil_SimpleDualBram_20_addrb;
  wire       [10:0]   xil_SimpleDualBram_21_addra;
  wire                xil_SimpleDualBram_21_ena;
  wire       [13:0]   xil_SimpleDualBram_21_addrb;
  wire       [10:0]   xil_SimpleDualBram_22_addra;
  wire                xil_SimpleDualBram_22_ena;
  wire       [13:0]   xil_SimpleDualBram_22_addrb;
  wire       [10:0]   xil_SimpleDualBram_23_addra;
  wire                xil_SimpleDualBram_23_ena;
  wire       [13:0]   xil_SimpleDualBram_23_addrb;
  wire       [10:0]   xil_SimpleDualBram_24_addra;
  wire                xil_SimpleDualBram_24_ena;
  wire       [13:0]   xil_SimpleDualBram_24_addrb;
  wire       [10:0]   xil_SimpleDualBram_25_addra;
  wire                xil_SimpleDualBram_25_ena;
  wire       [13:0]   xil_SimpleDualBram_25_addrb;
  wire       [10:0]   xil_SimpleDualBram_26_addra;
  wire                xil_SimpleDualBram_26_ena;
  wire       [13:0]   xil_SimpleDualBram_26_addrb;
  wire       [10:0]   xil_SimpleDualBram_27_addra;
  wire                xil_SimpleDualBram_27_ena;
  wire       [13:0]   xil_SimpleDualBram_27_addrb;
  wire       [10:0]   xil_SimpleDualBram_28_addra;
  wire                xil_SimpleDualBram_28_ena;
  wire       [13:0]   xil_SimpleDualBram_28_addrb;
  wire       [10:0]   xil_SimpleDualBram_29_addra;
  wire                xil_SimpleDualBram_29_ena;
  wire       [13:0]   xil_SimpleDualBram_29_addrb;
  wire       [10:0]   xil_SimpleDualBram_30_addra;
  wire                xil_SimpleDualBram_30_ena;
  wire       [13:0]   xil_SimpleDualBram_30_addrb;
  wire       [10:0]   xil_SimpleDualBram_31_addra;
  wire                xil_SimpleDualBram_31_ena;
  wire       [13:0]   xil_SimpleDualBram_31_addrb;
  wire       [10:0]   xil_SimpleDualBram_32_addra;
  wire                xil_SimpleDualBram_32_ena;
  wire       [13:0]   xil_SimpleDualBram_32_addrb;
  wire       [10:0]   xil_SimpleDualBram_33_addra;
  wire                xil_SimpleDualBram_33_ena;
  wire       [13:0]   xil_SimpleDualBram_33_addrb;
  wire       [10:0]   xil_SimpleDualBram_34_addra;
  wire                xil_SimpleDualBram_34_ena;
  wire       [13:0]   xil_SimpleDualBram_34_addrb;
  wire       [10:0]   xil_SimpleDualBram_35_addra;
  wire                xil_SimpleDualBram_35_ena;
  wire       [13:0]   xil_SimpleDualBram_35_addrb;
  wire       [10:0]   xil_SimpleDualBram_36_addra;
  wire                xil_SimpleDualBram_36_ena;
  wire       [13:0]   xil_SimpleDualBram_36_addrb;
  wire       [10:0]   xil_SimpleDualBram_37_addra;
  wire                xil_SimpleDualBram_37_ena;
  wire       [13:0]   xil_SimpleDualBram_37_addrb;
  wire       [10:0]   xil_SimpleDualBram_38_addra;
  wire                xil_SimpleDualBram_38_ena;
  wire       [13:0]   xil_SimpleDualBram_38_addrb;
  wire       [10:0]   xil_SimpleDualBram_39_addra;
  wire                xil_SimpleDualBram_39_ena;
  wire       [13:0]   xil_SimpleDualBram_39_addrb;
  wire       [10:0]   xil_SimpleDualBram_40_addra;
  wire                xil_SimpleDualBram_40_ena;
  wire       [13:0]   xil_SimpleDualBram_40_addrb;
  wire       [10:0]   xil_SimpleDualBram_41_addra;
  wire                xil_SimpleDualBram_41_ena;
  wire       [13:0]   xil_SimpleDualBram_41_addrb;
  wire       [10:0]   xil_SimpleDualBram_42_addra;
  wire                xil_SimpleDualBram_42_ena;
  wire       [13:0]   xil_SimpleDualBram_42_addrb;
  wire       [10:0]   xil_SimpleDualBram_43_addra;
  wire                xil_SimpleDualBram_43_ena;
  wire       [13:0]   xil_SimpleDualBram_43_addrb;
  wire       [10:0]   xil_SimpleDualBram_44_addra;
  wire                xil_SimpleDualBram_44_ena;
  wire       [13:0]   xil_SimpleDualBram_44_addrb;
  wire       [10:0]   xil_SimpleDualBram_45_addra;
  wire                xil_SimpleDualBram_45_ena;
  wire       [13:0]   xil_SimpleDualBram_45_addrb;
  wire       [10:0]   xil_SimpleDualBram_46_addra;
  wire                xil_SimpleDualBram_46_ena;
  wire       [13:0]   xil_SimpleDualBram_46_addrb;
  wire       [10:0]   xil_SimpleDualBram_47_addra;
  wire                xil_SimpleDualBram_47_ena;
  wire       [13:0]   xil_SimpleDualBram_47_addrb;
  wire       [10:0]   xil_SimpleDualBram_48_addra;
  wire                xil_SimpleDualBram_48_ena;
  wire       [13:0]   xil_SimpleDualBram_48_addrb;
  wire       [10:0]   xil_SimpleDualBram_49_addra;
  wire                xil_SimpleDualBram_49_ena;
  wire       [13:0]   xil_SimpleDualBram_49_addrb;
  wire       [10:0]   xil_SimpleDualBram_50_addra;
  wire                xil_SimpleDualBram_50_ena;
  wire       [13:0]   xil_SimpleDualBram_50_addrb;
  wire       [10:0]   xil_SimpleDualBram_51_addra;
  wire                xil_SimpleDualBram_51_ena;
  wire       [13:0]   xil_SimpleDualBram_51_addrb;
  wire       [10:0]   xil_SimpleDualBram_52_addra;
  wire                xil_SimpleDualBram_52_ena;
  wire       [13:0]   xil_SimpleDualBram_52_addrb;
  wire       [10:0]   xil_SimpleDualBram_53_addra;
  wire                xil_SimpleDualBram_53_ena;
  wire       [13:0]   xil_SimpleDualBram_53_addrb;
  wire       [10:0]   xil_SimpleDualBram_54_addra;
  wire                xil_SimpleDualBram_54_ena;
  wire       [13:0]   xil_SimpleDualBram_54_addrb;
  wire       [10:0]   xil_SimpleDualBram_55_addra;
  wire                xil_SimpleDualBram_55_ena;
  wire       [13:0]   xil_SimpleDualBram_55_addrb;
  wire       [10:0]   xil_SimpleDualBram_56_addra;
  wire                xil_SimpleDualBram_56_ena;
  wire       [13:0]   xil_SimpleDualBram_56_addrb;
  wire       [10:0]   xil_SimpleDualBram_57_addra;
  wire                xil_SimpleDualBram_57_ena;
  wire       [13:0]   xil_SimpleDualBram_57_addrb;
  wire       [10:0]   xil_SimpleDualBram_58_addra;
  wire                xil_SimpleDualBram_58_ena;
  wire       [13:0]   xil_SimpleDualBram_58_addrb;
  wire       [10:0]   xil_SimpleDualBram_59_addra;
  wire                xil_SimpleDualBram_59_ena;
  wire       [13:0]   xil_SimpleDualBram_59_addrb;
  wire       [10:0]   xil_SimpleDualBram_60_addra;
  wire                xil_SimpleDualBram_60_ena;
  wire       [13:0]   xil_SimpleDualBram_60_addrb;
  wire       [10:0]   xil_SimpleDualBram_61_addra;
  wire                xil_SimpleDualBram_61_ena;
  wire       [13:0]   xil_SimpleDualBram_61_addrb;
  wire       [10:0]   xil_SimpleDualBram_62_addra;
  wire                xil_SimpleDualBram_62_ena;
  wire       [13:0]   xil_SimpleDualBram_62_addrb;
  wire       [10:0]   xil_SimpleDualBram_63_addra;
  wire                xil_SimpleDualBram_63_ena;
  wire       [13:0]   xil_SimpleDualBram_63_addrb;
  wire       [7:0]    xil_SimpleDualBram_doutb;
  wire       [7:0]    xil_SimpleDualBram_1_doutb;
  wire       [7:0]    xil_SimpleDualBram_2_doutb;
  wire       [7:0]    xil_SimpleDualBram_3_doutb;
  wire       [7:0]    xil_SimpleDualBram_4_doutb;
  wire       [7:0]    xil_SimpleDualBram_5_doutb;
  wire       [7:0]    xil_SimpleDualBram_6_doutb;
  wire       [7:0]    xil_SimpleDualBram_7_doutb;
  wire       [7:0]    xil_SimpleDualBram_8_doutb;
  wire       [7:0]    xil_SimpleDualBram_9_doutb;
  wire       [7:0]    xil_SimpleDualBram_10_doutb;
  wire       [7:0]    xil_SimpleDualBram_11_doutb;
  wire       [7:0]    xil_SimpleDualBram_12_doutb;
  wire       [7:0]    xil_SimpleDualBram_13_doutb;
  wire       [7:0]    xil_SimpleDualBram_14_doutb;
  wire       [7:0]    xil_SimpleDualBram_15_doutb;
  wire       [7:0]    xil_SimpleDualBram_16_doutb;
  wire       [7:0]    xil_SimpleDualBram_17_doutb;
  wire       [7:0]    xil_SimpleDualBram_18_doutb;
  wire       [7:0]    xil_SimpleDualBram_19_doutb;
  wire       [7:0]    xil_SimpleDualBram_20_doutb;
  wire       [7:0]    xil_SimpleDualBram_21_doutb;
  wire       [7:0]    xil_SimpleDualBram_22_doutb;
  wire       [7:0]    xil_SimpleDualBram_23_doutb;
  wire       [7:0]    xil_SimpleDualBram_24_doutb;
  wire       [7:0]    xil_SimpleDualBram_25_doutb;
  wire       [7:0]    xil_SimpleDualBram_26_doutb;
  wire       [7:0]    xil_SimpleDualBram_27_doutb;
  wire       [7:0]    xil_SimpleDualBram_28_doutb;
  wire       [7:0]    xil_SimpleDualBram_29_doutb;
  wire       [7:0]    xil_SimpleDualBram_30_doutb;
  wire       [7:0]    xil_SimpleDualBram_31_doutb;
  wire       [7:0]    xil_SimpleDualBram_32_doutb;
  wire       [7:0]    xil_SimpleDualBram_33_doutb;
  wire       [7:0]    xil_SimpleDualBram_34_doutb;
  wire       [7:0]    xil_SimpleDualBram_35_doutb;
  wire       [7:0]    xil_SimpleDualBram_36_doutb;
  wire       [7:0]    xil_SimpleDualBram_37_doutb;
  wire       [7:0]    xil_SimpleDualBram_38_doutb;
  wire       [7:0]    xil_SimpleDualBram_39_doutb;
  wire       [7:0]    xil_SimpleDualBram_40_doutb;
  wire       [7:0]    xil_SimpleDualBram_41_doutb;
  wire       [7:0]    xil_SimpleDualBram_42_doutb;
  wire       [7:0]    xil_SimpleDualBram_43_doutb;
  wire       [7:0]    xil_SimpleDualBram_44_doutb;
  wire       [7:0]    xil_SimpleDualBram_45_doutb;
  wire       [7:0]    xil_SimpleDualBram_46_doutb;
  wire       [7:0]    xil_SimpleDualBram_47_doutb;
  wire       [7:0]    xil_SimpleDualBram_48_doutb;
  wire       [7:0]    xil_SimpleDualBram_49_doutb;
  wire       [7:0]    xil_SimpleDualBram_50_doutb;
  wire       [7:0]    xil_SimpleDualBram_51_doutb;
  wire       [7:0]    xil_SimpleDualBram_52_doutb;
  wire       [7:0]    xil_SimpleDualBram_53_doutb;
  wire       [7:0]    xil_SimpleDualBram_54_doutb;
  wire       [7:0]    xil_SimpleDualBram_55_doutb;
  wire       [7:0]    xil_SimpleDualBram_56_doutb;
  wire       [7:0]    xil_SimpleDualBram_57_doutb;
  wire       [7:0]    xil_SimpleDualBram_58_doutb;
  wire       [7:0]    xil_SimpleDualBram_59_doutb;
  wire       [7:0]    xil_SimpleDualBram_60_doutb;
  wire       [7:0]    xil_SimpleDualBram_61_doutb;
  wire       [7:0]    xil_SimpleDualBram_62_doutb;
  wire       [7:0]    xil_SimpleDualBram_63_doutb;
  wire       [15:0]   _zz_In_Row_Cnt_valid;
  wire       [12:0]   _zz_In_Row_Cnt_valid_1;
  wire       [15:0]   _zz_In_Col_Cnt_valid;
  wire       [15:0]   _zz_OutRow_Cnt_valid;
  wire       [15:0]   _zz_OutCol_Cnt_valid;
  wire       [15:0]   _zz_OutCol_Cnt_count_1;
  wire       [15:0]   _zz_Write_Row_Base_Addr;
  wire       [15:0]   _zz_addra;
  wire       [15:0]   _zz_addrb;
  wire       [0:0]    _zz_ena;
  wire       [15:0]   _zz_addra_1;
  wire       [15:0]   _zz_addrb_1;
  wire       [0:0]    _zz_ena_1;
  wire       [15:0]   _zz_addra_2;
  wire       [15:0]   _zz_addrb_2;
  wire       [0:0]    _zz_ena_2;
  wire       [15:0]   _zz_addra_3;
  wire       [15:0]   _zz_addrb_3;
  wire       [0:0]    _zz_ena_3;
  wire       [15:0]   _zz_addra_4;
  wire       [15:0]   _zz_addrb_4;
  wire       [0:0]    _zz_ena_4;
  wire       [15:0]   _zz_addra_5;
  wire       [15:0]   _zz_addrb_5;
  wire       [0:0]    _zz_ena_5;
  wire       [15:0]   _zz_addra_6;
  wire       [15:0]   _zz_addrb_6;
  wire       [0:0]    _zz_ena_6;
  wire       [15:0]   _zz_addra_7;
  wire       [15:0]   _zz_addrb_7;
  wire       [0:0]    _zz_ena_7;
  wire       [15:0]   _zz_addra_8;
  wire       [15:0]   _zz_addrb_8;
  wire       [0:0]    _zz_ena_8;
  wire       [15:0]   _zz_addra_9;
  wire       [15:0]   _zz_addrb_9;
  wire       [0:0]    _zz_ena_9;
  wire       [15:0]   _zz_addra_10;
  wire       [15:0]   _zz_addrb_10;
  wire       [0:0]    _zz_ena_10;
  wire       [15:0]   _zz_addra_11;
  wire       [15:0]   _zz_addrb_11;
  wire       [0:0]    _zz_ena_11;
  wire       [15:0]   _zz_addra_12;
  wire       [15:0]   _zz_addrb_12;
  wire       [0:0]    _zz_ena_12;
  wire       [15:0]   _zz_addra_13;
  wire       [15:0]   _zz_addrb_13;
  wire       [0:0]    _zz_ena_13;
  wire       [15:0]   _zz_addra_14;
  wire       [15:0]   _zz_addrb_14;
  wire       [0:0]    _zz_ena_14;
  wire       [15:0]   _zz_addra_15;
  wire       [15:0]   _zz_addrb_15;
  wire       [0:0]    _zz_ena_15;
  wire       [15:0]   _zz_addra_16;
  wire       [15:0]   _zz_addrb_16;
  wire       [0:0]    _zz_ena_16;
  wire       [15:0]   _zz_addra_17;
  wire       [15:0]   _zz_addrb_17;
  wire       [0:0]    _zz_ena_17;
  wire       [15:0]   _zz_addra_18;
  wire       [15:0]   _zz_addrb_18;
  wire       [0:0]    _zz_ena_18;
  wire       [15:0]   _zz_addra_19;
  wire       [15:0]   _zz_addrb_19;
  wire       [0:0]    _zz_ena_19;
  wire       [15:0]   _zz_addra_20;
  wire       [15:0]   _zz_addrb_20;
  wire       [0:0]    _zz_ena_20;
  wire       [15:0]   _zz_addra_21;
  wire       [15:0]   _zz_addrb_21;
  wire       [0:0]    _zz_ena_21;
  wire       [15:0]   _zz_addra_22;
  wire       [15:0]   _zz_addrb_22;
  wire       [0:0]    _zz_ena_22;
  wire       [15:0]   _zz_addra_23;
  wire       [15:0]   _zz_addrb_23;
  wire       [0:0]    _zz_ena_23;
  wire       [15:0]   _zz_addra_24;
  wire       [15:0]   _zz_addrb_24;
  wire       [0:0]    _zz_ena_24;
  wire       [15:0]   _zz_addra_25;
  wire       [15:0]   _zz_addrb_25;
  wire       [0:0]    _zz_ena_25;
  wire       [15:0]   _zz_addra_26;
  wire       [15:0]   _zz_addrb_26;
  wire       [0:0]    _zz_ena_26;
  wire       [15:0]   _zz_addra_27;
  wire       [15:0]   _zz_addrb_27;
  wire       [0:0]    _zz_ena_27;
  wire       [15:0]   _zz_addra_28;
  wire       [15:0]   _zz_addrb_28;
  wire       [0:0]    _zz_ena_28;
  wire       [15:0]   _zz_addra_29;
  wire       [15:0]   _zz_addrb_29;
  wire       [0:0]    _zz_ena_29;
  wire       [15:0]   _zz_addra_30;
  wire       [15:0]   _zz_addrb_30;
  wire       [0:0]    _zz_ena_30;
  wire       [15:0]   _zz_addra_31;
  wire       [15:0]   _zz_addrb_31;
  wire       [0:0]    _zz_ena_31;
  wire       [15:0]   _zz_addra_32;
  wire       [15:0]   _zz_addrb_32;
  wire       [0:0]    _zz_ena_32;
  wire       [15:0]   _zz_addra_33;
  wire       [15:0]   _zz_addrb_33;
  wire       [0:0]    _zz_ena_33;
  wire       [15:0]   _zz_addra_34;
  wire       [15:0]   _zz_addrb_34;
  wire       [0:0]    _zz_ena_34;
  wire       [15:0]   _zz_addra_35;
  wire       [15:0]   _zz_addrb_35;
  wire       [0:0]    _zz_ena_35;
  wire       [15:0]   _zz_addra_36;
  wire       [15:0]   _zz_addrb_36;
  wire       [0:0]    _zz_ena_36;
  wire       [15:0]   _zz_addra_37;
  wire       [15:0]   _zz_addrb_37;
  wire       [0:0]    _zz_ena_37;
  wire       [15:0]   _zz_addra_38;
  wire       [15:0]   _zz_addrb_38;
  wire       [0:0]    _zz_ena_38;
  wire       [15:0]   _zz_addra_39;
  wire       [15:0]   _zz_addrb_39;
  wire       [0:0]    _zz_ena_39;
  wire       [15:0]   _zz_addra_40;
  wire       [15:0]   _zz_addrb_40;
  wire       [0:0]    _zz_ena_40;
  wire       [15:0]   _zz_addra_41;
  wire       [15:0]   _zz_addrb_41;
  wire       [0:0]    _zz_ena_41;
  wire       [15:0]   _zz_addra_42;
  wire       [15:0]   _zz_addrb_42;
  wire       [0:0]    _zz_ena_42;
  wire       [15:0]   _zz_addra_43;
  wire       [15:0]   _zz_addrb_43;
  wire       [0:0]    _zz_ena_43;
  wire       [15:0]   _zz_addra_44;
  wire       [15:0]   _zz_addrb_44;
  wire       [0:0]    _zz_ena_44;
  wire       [15:0]   _zz_addra_45;
  wire       [15:0]   _zz_addrb_45;
  wire       [0:0]    _zz_ena_45;
  wire       [15:0]   _zz_addra_46;
  wire       [15:0]   _zz_addrb_46;
  wire       [0:0]    _zz_ena_46;
  wire       [15:0]   _zz_addra_47;
  wire       [15:0]   _zz_addrb_47;
  wire       [0:0]    _zz_ena_47;
  wire       [15:0]   _zz_addra_48;
  wire       [15:0]   _zz_addrb_48;
  wire       [0:0]    _zz_ena_48;
  wire       [15:0]   _zz_addra_49;
  wire       [15:0]   _zz_addrb_49;
  wire       [0:0]    _zz_ena_49;
  wire       [15:0]   _zz_addra_50;
  wire       [15:0]   _zz_addrb_50;
  wire       [0:0]    _zz_ena_50;
  wire       [15:0]   _zz_addra_51;
  wire       [15:0]   _zz_addrb_51;
  wire       [0:0]    _zz_ena_51;
  wire       [15:0]   _zz_addra_52;
  wire       [15:0]   _zz_addrb_52;
  wire       [0:0]    _zz_ena_52;
  wire       [15:0]   _zz_addra_53;
  wire       [15:0]   _zz_addrb_53;
  wire       [0:0]    _zz_ena_53;
  wire       [15:0]   _zz_addra_54;
  wire       [15:0]   _zz_addrb_54;
  wire       [0:0]    _zz_ena_54;
  wire       [15:0]   _zz_addra_55;
  wire       [15:0]   _zz_addrb_55;
  wire       [0:0]    _zz_ena_55;
  wire       [15:0]   _zz_addra_56;
  wire       [15:0]   _zz_addrb_56;
  wire       [0:0]    _zz_ena_56;
  wire       [15:0]   _zz_addra_57;
  wire       [15:0]   _zz_addrb_57;
  wire       [0:0]    _zz_ena_57;
  wire       [15:0]   _zz_addra_58;
  wire       [15:0]   _zz_addrb_58;
  wire       [0:0]    _zz_ena_58;
  wire       [15:0]   _zz_addra_59;
  wire       [15:0]   _zz_addrb_59;
  wire       [0:0]    _zz_ena_59;
  wire       [15:0]   _zz_addra_60;
  wire       [15:0]   _zz_addrb_60;
  wire       [0:0]    _zz_ena_60;
  wire       [15:0]   _zz_addra_61;
  wire       [15:0]   _zz_addrb_61;
  wire       [0:0]    _zz_ena_61;
  wire       [15:0]   _zz_addra_62;
  wire       [15:0]   _zz_addrb_62;
  wire       [0:0]    _zz_ena_62;
  wire       [15:0]   _zz_addra_63;
  wire       [15:0]   _zz_addrb_63;
  wire       [0:0]    _zz_ena_63;
  reg                 start_regNext;
  wire                when_SA3D_WeightCache_l33;
  reg        [3:0]    Fsm_currentState;
  reg        [3:0]    Fsm_nextState;
  wire                Fsm_Init_End;
  wire                Fsm_Weight_All_Cached;
  wire                Fsm_SA_Computed;
  wire                when_WaCounter_l19;
  reg        [2:0]    Init_Count_count;
  reg                 Init_Count_valid;
  wire                when_WaCounter_l14;
  reg        [63:0]   InData_Switch;
  wire       [12:0]   Matrix_In_MaxCnt;
  wire                sData_fire;
  reg        [15:0]   In_Row_Cnt_count;
  wire                In_Row_Cnt_valid;
  reg        [15:0]   In_Col_Cnt_count;
  wire                In_Col_Cnt_valid;
  reg        [15:0]   Read_Row_Base_Addr;
  reg        [15:0]   Write_Row_Base_Addr;
  wire                when_WaCounter_l40;
  reg        [15:0]   OutRow_Cnt_count;
  wire                OutRow_Cnt_valid;
  wire       [3:0]    _zz_OutCol_Cnt_count;
  reg        [15:0]   OutCol_Cnt_count;
  reg                 OutCol_Cnt_valid;
  reg        [5:0]    Col_In_8_Cnt_count;
  reg                 Col_In_8_Cnt_valid;
  wire                when_SA3D_WeightCache_l129;
  wire                when_SA3D_WeightCache_l134;
  wire                sData_fire_1;
  wire                sData_fire_2;
  wire                sData_fire_3;
  wire                sData_fire_4;
  wire                sData_fire_5;
  wire                sData_fire_6;
  wire                sData_fire_7;
  wire                sData_fire_8;
  wire                sData_fire_9;
  wire                sData_fire_10;
  wire                sData_fire_11;
  wire                sData_fire_12;
  wire                sData_fire_13;
  wire                sData_fire_14;
  wire                sData_fire_15;
  wire                sData_fire_16;
  wire                sData_fire_17;
  wire                sData_fire_18;
  wire                sData_fire_19;
  wire                sData_fire_20;
  wire                sData_fire_21;
  wire                sData_fire_22;
  wire                sData_fire_23;
  wire                sData_fire_24;
  wire                sData_fire_25;
  wire                sData_fire_26;
  wire                sData_fire_27;
  wire                sData_fire_28;
  wire                sData_fire_29;
  wire                sData_fire_30;
  wire                sData_fire_31;
  wire                sData_fire_32;
  wire                sData_fire_33;
  wire                sData_fire_34;
  wire                sData_fire_35;
  wire                sData_fire_36;
  wire                sData_fire_37;
  wire                sData_fire_38;
  wire                sData_fire_39;
  wire                sData_fire_40;
  wire                sData_fire_41;
  wire                sData_fire_42;
  wire                sData_fire_43;
  wire                sData_fire_44;
  wire                sData_fire_45;
  wire                sData_fire_46;
  wire                sData_fire_47;
  wire                sData_fire_48;
  wire                sData_fire_49;
  wire                sData_fire_50;
  wire                sData_fire_51;
  wire                sData_fire_52;
  wire                sData_fire_53;
  wire                sData_fire_54;
  wire                sData_fire_55;
  wire                sData_fire_56;
  wire                sData_fire_57;
  wire                sData_fire_58;
  wire                sData_fire_59;
  wire                sData_fire_60;
  wire                sData_fire_61;
  wire                sData_fire_62;
  wire                sData_fire_63;
  wire                sData_fire_64;
  reg        [7:0]    MatrixCol_Switch_1;
  reg        [7:0]    MatrixCol_Switch_1_regNext;
  `ifndef SYNTHESIS
  reg [95:0] Fsm_currentState_string;
  reg [95:0] Fsm_nextState_string;
  `endif


  assign _zz_In_Row_Cnt_valid_1 = (Matrix_In_MaxCnt - 13'h0001);
  assign _zz_In_Row_Cnt_valid = {3'd0, _zz_In_Row_Cnt_valid_1};
  assign _zz_In_Col_Cnt_valid = (Matrix_Col - 16'h0001);
  assign _zz_OutRow_Cnt_valid = (Matrix_Row - 16'h0001);
  assign _zz_OutCol_Cnt_valid = {12'd0, _zz_OutCol_Cnt_count};
  assign _zz_OutCol_Cnt_count_1 = {12'd0, _zz_OutCol_Cnt_count};
  assign _zz_Write_Row_Base_Addr = {3'd0, Matrix_In_MaxCnt};
  assign _zz_addra = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena = InData_Switch[0 : 0];
  assign _zz_addra_1 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_1 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_1 = InData_Switch[1 : 1];
  assign _zz_addra_2 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_2 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_2 = InData_Switch[2 : 2];
  assign _zz_addra_3 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_3 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_3 = InData_Switch[3 : 3];
  assign _zz_addra_4 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_4 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_4 = InData_Switch[4 : 4];
  assign _zz_addra_5 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_5 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_5 = InData_Switch[5 : 5];
  assign _zz_addra_6 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_6 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_6 = InData_Switch[6 : 6];
  assign _zz_addra_7 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_7 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_7 = InData_Switch[7 : 7];
  assign _zz_addra_8 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_8 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_8 = InData_Switch[8 : 8];
  assign _zz_addra_9 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_9 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_9 = InData_Switch[9 : 9];
  assign _zz_addra_10 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_10 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_10 = InData_Switch[10 : 10];
  assign _zz_addra_11 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_11 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_11 = InData_Switch[11 : 11];
  assign _zz_addra_12 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_12 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_12 = InData_Switch[12 : 12];
  assign _zz_addra_13 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_13 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_13 = InData_Switch[13 : 13];
  assign _zz_addra_14 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_14 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_14 = InData_Switch[14 : 14];
  assign _zz_addra_15 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_15 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_15 = InData_Switch[15 : 15];
  assign _zz_addra_16 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_16 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_16 = InData_Switch[16 : 16];
  assign _zz_addra_17 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_17 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_17 = InData_Switch[17 : 17];
  assign _zz_addra_18 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_18 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_18 = InData_Switch[18 : 18];
  assign _zz_addra_19 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_19 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_19 = InData_Switch[19 : 19];
  assign _zz_addra_20 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_20 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_20 = InData_Switch[20 : 20];
  assign _zz_addra_21 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_21 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_21 = InData_Switch[21 : 21];
  assign _zz_addra_22 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_22 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_22 = InData_Switch[22 : 22];
  assign _zz_addra_23 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_23 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_23 = InData_Switch[23 : 23];
  assign _zz_addra_24 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_24 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_24 = InData_Switch[24 : 24];
  assign _zz_addra_25 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_25 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_25 = InData_Switch[25 : 25];
  assign _zz_addra_26 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_26 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_26 = InData_Switch[26 : 26];
  assign _zz_addra_27 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_27 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_27 = InData_Switch[27 : 27];
  assign _zz_addra_28 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_28 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_28 = InData_Switch[28 : 28];
  assign _zz_addra_29 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_29 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_29 = InData_Switch[29 : 29];
  assign _zz_addra_30 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_30 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_30 = InData_Switch[30 : 30];
  assign _zz_addra_31 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_31 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_31 = InData_Switch[31 : 31];
  assign _zz_addra_32 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_32 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_32 = InData_Switch[32 : 32];
  assign _zz_addra_33 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_33 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_33 = InData_Switch[33 : 33];
  assign _zz_addra_34 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_34 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_34 = InData_Switch[34 : 34];
  assign _zz_addra_35 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_35 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_35 = InData_Switch[35 : 35];
  assign _zz_addra_36 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_36 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_36 = InData_Switch[36 : 36];
  assign _zz_addra_37 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_37 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_37 = InData_Switch[37 : 37];
  assign _zz_addra_38 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_38 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_38 = InData_Switch[38 : 38];
  assign _zz_addra_39 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_39 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_39 = InData_Switch[39 : 39];
  assign _zz_addra_40 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_40 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_40 = InData_Switch[40 : 40];
  assign _zz_addra_41 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_41 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_41 = InData_Switch[41 : 41];
  assign _zz_addra_42 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_42 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_42 = InData_Switch[42 : 42];
  assign _zz_addra_43 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_43 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_43 = InData_Switch[43 : 43];
  assign _zz_addra_44 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_44 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_44 = InData_Switch[44 : 44];
  assign _zz_addra_45 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_45 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_45 = InData_Switch[45 : 45];
  assign _zz_addra_46 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_46 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_46 = InData_Switch[46 : 46];
  assign _zz_addra_47 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_47 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_47 = InData_Switch[47 : 47];
  assign _zz_addra_48 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_48 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_48 = InData_Switch[48 : 48];
  assign _zz_addra_49 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_49 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_49 = InData_Switch[49 : 49];
  assign _zz_addra_50 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_50 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_50 = InData_Switch[50 : 50];
  assign _zz_addra_51 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_51 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_51 = InData_Switch[51 : 51];
  assign _zz_addra_52 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_52 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_52 = InData_Switch[52 : 52];
  assign _zz_addra_53 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_53 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_53 = InData_Switch[53 : 53];
  assign _zz_addra_54 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_54 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_54 = InData_Switch[54 : 54];
  assign _zz_addra_55 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_55 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_55 = InData_Switch[55 : 55];
  assign _zz_addra_56 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_56 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_56 = InData_Switch[56 : 56];
  assign _zz_addra_57 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_57 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_57 = InData_Switch[57 : 57];
  assign _zz_addra_58 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_58 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_58 = InData_Switch[58 : 58];
  assign _zz_addra_59 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_59 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_59 = InData_Switch[59 : 59];
  assign _zz_addra_60 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_60 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_60 = InData_Switch[60 : 60];
  assign _zz_addra_61 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_61 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_61 = InData_Switch[61 : 61];
  assign _zz_addra_62 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_62 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_62 = InData_Switch[62 : 62];
  assign _zz_addra_63 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_63 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_63 = InData_Switch[63 : 63];
  Weight_Bram xil_SimpleDualBram (
    .clka  (clk                           ), //i
    .addra (xil_SimpleDualBram_addra[10:0]), //i
    .dina  (sData_payload[63:0]           ), //i
    .ena   (xil_SimpleDualBram_ena        ), //i
    .wea   (1'b1                          ), //i
    .addrb (xil_SimpleDualBram_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_doutb[7:0] ), //o
    .clkb  (clk                           )  //i
  );
  Weight_Bram xil_SimpleDualBram_1 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_1_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_1_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_1_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_1_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_2 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_2_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_2_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_2_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_2_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_3 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_3_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_3_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_3_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_3_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_4 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_4_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_4_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_4_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_4_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_5 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_5_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_5_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_5_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_5_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_6 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_6_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_6_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_6_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_6_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_7 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_7_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_7_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_7_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_7_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_8 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_8_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_8_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_8_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_8_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_9 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_9_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_9_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_9_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_9_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_10 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_10_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_10_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_10_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_10_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_11 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_11_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_11_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_11_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_11_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_12 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_12_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_12_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_12_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_12_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_13 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_13_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_13_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_13_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_13_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_14 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_14_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_14_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_14_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_14_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_15 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_15_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_15_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_15_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_15_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_16 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_16_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_16_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_16_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_16_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_17 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_17_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_17_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_17_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_17_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_18 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_18_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_18_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_18_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_18_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_19 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_19_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_19_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_19_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_19_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_20 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_20_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_20_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_20_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_20_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_21 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_21_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_21_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_21_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_21_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_22 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_22_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_22_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_22_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_22_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_23 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_23_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_23_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_23_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_23_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_24 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_24_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_24_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_24_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_24_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_25 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_25_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_25_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_25_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_25_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_26 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_26_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_26_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_26_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_26_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_27 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_27_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_27_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_27_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_27_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_28 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_28_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_28_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_28_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_28_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_29 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_29_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_29_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_29_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_29_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_30 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_30_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_30_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_30_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_30_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_31 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_31_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_31_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_31_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_31_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_32 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_32_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_32_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_32_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_32_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_33 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_33_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_33_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_33_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_33_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_34 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_34_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_34_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_34_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_34_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_35 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_35_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_35_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_35_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_35_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_36 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_36_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_36_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_36_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_36_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_37 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_37_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_37_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_37_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_37_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_38 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_38_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_38_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_38_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_38_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_39 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_39_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_39_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_39_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_39_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_40 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_40_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_40_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_40_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_40_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_41 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_41_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_41_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_41_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_41_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_42 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_42_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_42_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_42_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_42_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_43 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_43_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_43_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_43_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_43_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_44 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_44_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_44_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_44_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_44_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_45 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_45_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_45_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_45_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_45_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_46 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_46_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_46_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_46_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_46_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_47 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_47_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_47_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_47_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_47_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_48 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_48_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_48_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_48_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_48_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_49 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_49_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_49_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_49_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_49_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_50 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_50_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_50_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_50_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_50_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_51 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_51_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_51_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_51_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_51_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_52 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_52_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_52_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_52_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_52_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_53 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_53_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_53_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_53_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_53_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_54 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_54_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_54_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_54_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_54_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_55 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_55_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_55_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_55_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_55_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_56 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_56_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_56_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_56_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_56_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_57 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_57_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_57_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_57_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_57_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_58 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_58_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_58_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_58_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_58_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_59 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_59_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_59_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_59_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_59_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_60 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_60_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_60_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_60_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_60_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_61 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_61_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_61_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_61_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_61_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_62 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_62_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_62_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_62_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_62_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_63 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_63_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_63_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_63_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_63_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      WEIGHT_CACHE_STATUS_IDLE : Fsm_currentState_string = "IDLE        ";
      WEIGHT_CACHE_STATUS_INIT : Fsm_currentState_string = "INIT        ";
      WEIGHT_CACHE_STATUS_CACHE_WEIGHT : Fsm_currentState_string = "CACHE_WEIGHT";
      WEIGHT_CACHE_STATUS_SA_COMPUTE : Fsm_currentState_string = "SA_COMPUTE  ";
      default : Fsm_currentState_string = "????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      WEIGHT_CACHE_STATUS_IDLE : Fsm_nextState_string = "IDLE        ";
      WEIGHT_CACHE_STATUS_INIT : Fsm_nextState_string = "INIT        ";
      WEIGHT_CACHE_STATUS_CACHE_WEIGHT : Fsm_nextState_string = "CACHE_WEIGHT";
      WEIGHT_CACHE_STATUS_SA_COMPUTE : Fsm_nextState_string = "SA_COMPUTE  ";
      default : Fsm_nextState_string = "????????????";
    endcase
  end
  `endif

  assign when_SA3D_WeightCache_l33 = (start && (! start_regNext));
  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & WEIGHT_CACHE_STATUS_IDLE) == WEIGHT_CACHE_STATUS_IDLE) : begin
        if(when_SA3D_WeightCache_l33) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_INIT;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_IDLE;
        end
      end
      (((Fsm_currentState) & WEIGHT_CACHE_STATUS_INIT) == WEIGHT_CACHE_STATUS_INIT) : begin
        if(Fsm_Init_End) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_CACHE_WEIGHT;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_INIT;
        end
      end
      (((Fsm_currentState) & WEIGHT_CACHE_STATUS_CACHE_WEIGHT) == WEIGHT_CACHE_STATUS_CACHE_WEIGHT) : begin
        if(Fsm_Weight_All_Cached) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_SA_COMPUTE;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_CACHE_WEIGHT;
        end
      end
      default : begin
        if(Fsm_SA_Computed) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_IDLE;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_SA_COMPUTE;
        end
      end
    endcase
  end

  assign when_WaCounter_l19 = ((Fsm_currentState & WEIGHT_CACHE_STATUS_INIT) != 4'b0000);
  assign when_WaCounter_l14 = (Init_Count_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l14) begin
      Init_Count_valid = 1'b1;
    end else begin
      Init_Count_valid = 1'b0;
    end
  end

  assign Fsm_Init_End = Init_Count_valid;
  assign Matrix_In_MaxCnt = (Matrix_Row >>> 3);
  assign sData_fire = (sData_valid && sData_ready);
  assign In_Row_Cnt_valid = ((In_Row_Cnt_count == _zz_In_Row_Cnt_valid) && sData_fire);
  assign In_Col_Cnt_valid = ((In_Col_Cnt_count == _zz_In_Col_Cnt_valid) && In_Row_Cnt_valid);
  assign when_WaCounter_l40 = (Raddr_Valid && ((Fsm_currentState & WEIGHT_CACHE_STATUS_SA_COMPUTE) != 4'b0000));
  assign OutRow_Cnt_valid = ((OutRow_Cnt_count == _zz_OutRow_Cnt_valid) && when_WaCounter_l40);
  assign _zz_OutCol_Cnt_count = 4'b1000;
  always @(*) begin
    OutCol_Cnt_valid = ((OutCol_Cnt_count <= _zz_OutCol_Cnt_valid) && OutRow_Cnt_valid);
    if(start) begin
      OutCol_Cnt_valid = 1'b0;
    end
  end

  always @(*) begin
    Col_In_8_Cnt_valid = ((Col_In_8_Cnt_count == 6'h3f) && In_Row_Cnt_valid);
    if(OutCol_Cnt_valid) begin
      Col_In_8_Cnt_valid = 1'b0;
    end
  end

  assign when_SA3D_WeightCache_l129 = ((Fsm_currentState & WEIGHT_CACHE_STATUS_INIT) != 4'b0000);
  assign when_SA3D_WeightCache_l134 = ((Fsm_currentState & WEIGHT_CACHE_STATUS_INIT) != 4'b0000);
  assign Fsm_Weight_All_Cached = In_Col_Cnt_valid;
  assign Weight_Cached = In_Col_Cnt_valid;
  assign xil_SimpleDualBram_addra = _zz_addra[10:0];
  assign xil_SimpleDualBram_addrb = _zz_addrb[13:0];
  assign sData_fire_1 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_ena = (_zz_ena[0] && sData_fire_1);
  assign mData_0 = xil_SimpleDualBram_doutb;
  assign xil_SimpleDualBram_1_addra = _zz_addra_1[10:0];
  assign xil_SimpleDualBram_1_addrb = _zz_addrb_1[13:0];
  assign sData_fire_2 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_1_ena = (_zz_ena_1[0] && sData_fire_2);
  assign mData_1 = xil_SimpleDualBram_1_doutb;
  assign xil_SimpleDualBram_2_addra = _zz_addra_2[10:0];
  assign xil_SimpleDualBram_2_addrb = _zz_addrb_2[13:0];
  assign sData_fire_3 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_2_ena = (_zz_ena_2[0] && sData_fire_3);
  assign mData_2 = xil_SimpleDualBram_2_doutb;
  assign xil_SimpleDualBram_3_addra = _zz_addra_3[10:0];
  assign xil_SimpleDualBram_3_addrb = _zz_addrb_3[13:0];
  assign sData_fire_4 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_3_ena = (_zz_ena_3[0] && sData_fire_4);
  assign mData_3 = xil_SimpleDualBram_3_doutb;
  assign xil_SimpleDualBram_4_addra = _zz_addra_4[10:0];
  assign xil_SimpleDualBram_4_addrb = _zz_addrb_4[13:0];
  assign sData_fire_5 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_4_ena = (_zz_ena_4[0] && sData_fire_5);
  assign mData_4 = xil_SimpleDualBram_4_doutb;
  assign xil_SimpleDualBram_5_addra = _zz_addra_5[10:0];
  assign xil_SimpleDualBram_5_addrb = _zz_addrb_5[13:0];
  assign sData_fire_6 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_5_ena = (_zz_ena_5[0] && sData_fire_6);
  assign mData_5 = xil_SimpleDualBram_5_doutb;
  assign xil_SimpleDualBram_6_addra = _zz_addra_6[10:0];
  assign xil_SimpleDualBram_6_addrb = _zz_addrb_6[13:0];
  assign sData_fire_7 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_6_ena = (_zz_ena_6[0] && sData_fire_7);
  assign mData_6 = xil_SimpleDualBram_6_doutb;
  assign xil_SimpleDualBram_7_addra = _zz_addra_7[10:0];
  assign xil_SimpleDualBram_7_addrb = _zz_addrb_7[13:0];
  assign sData_fire_8 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_7_ena = (_zz_ena_7[0] && sData_fire_8);
  assign mData_7 = xil_SimpleDualBram_7_doutb;
  assign xil_SimpleDualBram_8_addra = _zz_addra_8[10:0];
  assign xil_SimpleDualBram_8_addrb = _zz_addrb_8[13:0];
  assign sData_fire_9 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_8_ena = (_zz_ena_8[0] && sData_fire_9);
  assign mData_8 = xil_SimpleDualBram_8_doutb;
  assign xil_SimpleDualBram_9_addra = _zz_addra_9[10:0];
  assign xil_SimpleDualBram_9_addrb = _zz_addrb_9[13:0];
  assign sData_fire_10 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_9_ena = (_zz_ena_9[0] && sData_fire_10);
  assign mData_9 = xil_SimpleDualBram_9_doutb;
  assign xil_SimpleDualBram_10_addra = _zz_addra_10[10:0];
  assign xil_SimpleDualBram_10_addrb = _zz_addrb_10[13:0];
  assign sData_fire_11 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_10_ena = (_zz_ena_10[0] && sData_fire_11);
  assign mData_10 = xil_SimpleDualBram_10_doutb;
  assign xil_SimpleDualBram_11_addra = _zz_addra_11[10:0];
  assign xil_SimpleDualBram_11_addrb = _zz_addrb_11[13:0];
  assign sData_fire_12 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_11_ena = (_zz_ena_11[0] && sData_fire_12);
  assign mData_11 = xil_SimpleDualBram_11_doutb;
  assign xil_SimpleDualBram_12_addra = _zz_addra_12[10:0];
  assign xil_SimpleDualBram_12_addrb = _zz_addrb_12[13:0];
  assign sData_fire_13 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_12_ena = (_zz_ena_12[0] && sData_fire_13);
  assign mData_12 = xil_SimpleDualBram_12_doutb;
  assign xil_SimpleDualBram_13_addra = _zz_addra_13[10:0];
  assign xil_SimpleDualBram_13_addrb = _zz_addrb_13[13:0];
  assign sData_fire_14 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_13_ena = (_zz_ena_13[0] && sData_fire_14);
  assign mData_13 = xil_SimpleDualBram_13_doutb;
  assign xil_SimpleDualBram_14_addra = _zz_addra_14[10:0];
  assign xil_SimpleDualBram_14_addrb = _zz_addrb_14[13:0];
  assign sData_fire_15 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_14_ena = (_zz_ena_14[0] && sData_fire_15);
  assign mData_14 = xil_SimpleDualBram_14_doutb;
  assign xil_SimpleDualBram_15_addra = _zz_addra_15[10:0];
  assign xil_SimpleDualBram_15_addrb = _zz_addrb_15[13:0];
  assign sData_fire_16 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_15_ena = (_zz_ena_15[0] && sData_fire_16);
  assign mData_15 = xil_SimpleDualBram_15_doutb;
  assign xil_SimpleDualBram_16_addra = _zz_addra_16[10:0];
  assign xil_SimpleDualBram_16_addrb = _zz_addrb_16[13:0];
  assign sData_fire_17 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_16_ena = (_zz_ena_16[0] && sData_fire_17);
  assign mData_16 = xil_SimpleDualBram_16_doutb;
  assign xil_SimpleDualBram_17_addra = _zz_addra_17[10:0];
  assign xil_SimpleDualBram_17_addrb = _zz_addrb_17[13:0];
  assign sData_fire_18 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_17_ena = (_zz_ena_17[0] && sData_fire_18);
  assign mData_17 = xil_SimpleDualBram_17_doutb;
  assign xil_SimpleDualBram_18_addra = _zz_addra_18[10:0];
  assign xil_SimpleDualBram_18_addrb = _zz_addrb_18[13:0];
  assign sData_fire_19 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_18_ena = (_zz_ena_18[0] && sData_fire_19);
  assign mData_18 = xil_SimpleDualBram_18_doutb;
  assign xil_SimpleDualBram_19_addra = _zz_addra_19[10:0];
  assign xil_SimpleDualBram_19_addrb = _zz_addrb_19[13:0];
  assign sData_fire_20 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_19_ena = (_zz_ena_19[0] && sData_fire_20);
  assign mData_19 = xil_SimpleDualBram_19_doutb;
  assign xil_SimpleDualBram_20_addra = _zz_addra_20[10:0];
  assign xil_SimpleDualBram_20_addrb = _zz_addrb_20[13:0];
  assign sData_fire_21 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_20_ena = (_zz_ena_20[0] && sData_fire_21);
  assign mData_20 = xil_SimpleDualBram_20_doutb;
  assign xil_SimpleDualBram_21_addra = _zz_addra_21[10:0];
  assign xil_SimpleDualBram_21_addrb = _zz_addrb_21[13:0];
  assign sData_fire_22 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_21_ena = (_zz_ena_21[0] && sData_fire_22);
  assign mData_21 = xil_SimpleDualBram_21_doutb;
  assign xil_SimpleDualBram_22_addra = _zz_addra_22[10:0];
  assign xil_SimpleDualBram_22_addrb = _zz_addrb_22[13:0];
  assign sData_fire_23 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_22_ena = (_zz_ena_22[0] && sData_fire_23);
  assign mData_22 = xil_SimpleDualBram_22_doutb;
  assign xil_SimpleDualBram_23_addra = _zz_addra_23[10:0];
  assign xil_SimpleDualBram_23_addrb = _zz_addrb_23[13:0];
  assign sData_fire_24 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_23_ena = (_zz_ena_23[0] && sData_fire_24);
  assign mData_23 = xil_SimpleDualBram_23_doutb;
  assign xil_SimpleDualBram_24_addra = _zz_addra_24[10:0];
  assign xil_SimpleDualBram_24_addrb = _zz_addrb_24[13:0];
  assign sData_fire_25 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_24_ena = (_zz_ena_24[0] && sData_fire_25);
  assign mData_24 = xil_SimpleDualBram_24_doutb;
  assign xil_SimpleDualBram_25_addra = _zz_addra_25[10:0];
  assign xil_SimpleDualBram_25_addrb = _zz_addrb_25[13:0];
  assign sData_fire_26 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_25_ena = (_zz_ena_25[0] && sData_fire_26);
  assign mData_25 = xil_SimpleDualBram_25_doutb;
  assign xil_SimpleDualBram_26_addra = _zz_addra_26[10:0];
  assign xil_SimpleDualBram_26_addrb = _zz_addrb_26[13:0];
  assign sData_fire_27 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_26_ena = (_zz_ena_26[0] && sData_fire_27);
  assign mData_26 = xil_SimpleDualBram_26_doutb;
  assign xil_SimpleDualBram_27_addra = _zz_addra_27[10:0];
  assign xil_SimpleDualBram_27_addrb = _zz_addrb_27[13:0];
  assign sData_fire_28 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_27_ena = (_zz_ena_27[0] && sData_fire_28);
  assign mData_27 = xil_SimpleDualBram_27_doutb;
  assign xil_SimpleDualBram_28_addra = _zz_addra_28[10:0];
  assign xil_SimpleDualBram_28_addrb = _zz_addrb_28[13:0];
  assign sData_fire_29 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_28_ena = (_zz_ena_28[0] && sData_fire_29);
  assign mData_28 = xil_SimpleDualBram_28_doutb;
  assign xil_SimpleDualBram_29_addra = _zz_addra_29[10:0];
  assign xil_SimpleDualBram_29_addrb = _zz_addrb_29[13:0];
  assign sData_fire_30 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_29_ena = (_zz_ena_29[0] && sData_fire_30);
  assign mData_29 = xil_SimpleDualBram_29_doutb;
  assign xil_SimpleDualBram_30_addra = _zz_addra_30[10:0];
  assign xil_SimpleDualBram_30_addrb = _zz_addrb_30[13:0];
  assign sData_fire_31 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_30_ena = (_zz_ena_30[0] && sData_fire_31);
  assign mData_30 = xil_SimpleDualBram_30_doutb;
  assign xil_SimpleDualBram_31_addra = _zz_addra_31[10:0];
  assign xil_SimpleDualBram_31_addrb = _zz_addrb_31[13:0];
  assign sData_fire_32 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_31_ena = (_zz_ena_31[0] && sData_fire_32);
  assign mData_31 = xil_SimpleDualBram_31_doutb;
  assign xil_SimpleDualBram_32_addra = _zz_addra_32[10:0];
  assign xil_SimpleDualBram_32_addrb = _zz_addrb_32[13:0];
  assign sData_fire_33 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_32_ena = (_zz_ena_32[0] && sData_fire_33);
  assign mData_32 = xil_SimpleDualBram_32_doutb;
  assign xil_SimpleDualBram_33_addra = _zz_addra_33[10:0];
  assign xil_SimpleDualBram_33_addrb = _zz_addrb_33[13:0];
  assign sData_fire_34 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_33_ena = (_zz_ena_33[0] && sData_fire_34);
  assign mData_33 = xil_SimpleDualBram_33_doutb;
  assign xil_SimpleDualBram_34_addra = _zz_addra_34[10:0];
  assign xil_SimpleDualBram_34_addrb = _zz_addrb_34[13:0];
  assign sData_fire_35 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_34_ena = (_zz_ena_34[0] && sData_fire_35);
  assign mData_34 = xil_SimpleDualBram_34_doutb;
  assign xil_SimpleDualBram_35_addra = _zz_addra_35[10:0];
  assign xil_SimpleDualBram_35_addrb = _zz_addrb_35[13:0];
  assign sData_fire_36 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_35_ena = (_zz_ena_35[0] && sData_fire_36);
  assign mData_35 = xil_SimpleDualBram_35_doutb;
  assign xil_SimpleDualBram_36_addra = _zz_addra_36[10:0];
  assign xil_SimpleDualBram_36_addrb = _zz_addrb_36[13:0];
  assign sData_fire_37 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_36_ena = (_zz_ena_36[0] && sData_fire_37);
  assign mData_36 = xil_SimpleDualBram_36_doutb;
  assign xil_SimpleDualBram_37_addra = _zz_addra_37[10:0];
  assign xil_SimpleDualBram_37_addrb = _zz_addrb_37[13:0];
  assign sData_fire_38 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_37_ena = (_zz_ena_37[0] && sData_fire_38);
  assign mData_37 = xil_SimpleDualBram_37_doutb;
  assign xil_SimpleDualBram_38_addra = _zz_addra_38[10:0];
  assign xil_SimpleDualBram_38_addrb = _zz_addrb_38[13:0];
  assign sData_fire_39 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_38_ena = (_zz_ena_38[0] && sData_fire_39);
  assign mData_38 = xil_SimpleDualBram_38_doutb;
  assign xil_SimpleDualBram_39_addra = _zz_addra_39[10:0];
  assign xil_SimpleDualBram_39_addrb = _zz_addrb_39[13:0];
  assign sData_fire_40 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_39_ena = (_zz_ena_39[0] && sData_fire_40);
  assign mData_39 = xil_SimpleDualBram_39_doutb;
  assign xil_SimpleDualBram_40_addra = _zz_addra_40[10:0];
  assign xil_SimpleDualBram_40_addrb = _zz_addrb_40[13:0];
  assign sData_fire_41 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_40_ena = (_zz_ena_40[0] && sData_fire_41);
  assign mData_40 = xil_SimpleDualBram_40_doutb;
  assign xil_SimpleDualBram_41_addra = _zz_addra_41[10:0];
  assign xil_SimpleDualBram_41_addrb = _zz_addrb_41[13:0];
  assign sData_fire_42 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_41_ena = (_zz_ena_41[0] && sData_fire_42);
  assign mData_41 = xil_SimpleDualBram_41_doutb;
  assign xil_SimpleDualBram_42_addra = _zz_addra_42[10:0];
  assign xil_SimpleDualBram_42_addrb = _zz_addrb_42[13:0];
  assign sData_fire_43 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_42_ena = (_zz_ena_42[0] && sData_fire_43);
  assign mData_42 = xil_SimpleDualBram_42_doutb;
  assign xil_SimpleDualBram_43_addra = _zz_addra_43[10:0];
  assign xil_SimpleDualBram_43_addrb = _zz_addrb_43[13:0];
  assign sData_fire_44 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_43_ena = (_zz_ena_43[0] && sData_fire_44);
  assign mData_43 = xil_SimpleDualBram_43_doutb;
  assign xil_SimpleDualBram_44_addra = _zz_addra_44[10:0];
  assign xil_SimpleDualBram_44_addrb = _zz_addrb_44[13:0];
  assign sData_fire_45 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_44_ena = (_zz_ena_44[0] && sData_fire_45);
  assign mData_44 = xil_SimpleDualBram_44_doutb;
  assign xil_SimpleDualBram_45_addra = _zz_addra_45[10:0];
  assign xil_SimpleDualBram_45_addrb = _zz_addrb_45[13:0];
  assign sData_fire_46 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_45_ena = (_zz_ena_45[0] && sData_fire_46);
  assign mData_45 = xil_SimpleDualBram_45_doutb;
  assign xil_SimpleDualBram_46_addra = _zz_addra_46[10:0];
  assign xil_SimpleDualBram_46_addrb = _zz_addrb_46[13:0];
  assign sData_fire_47 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_46_ena = (_zz_ena_46[0] && sData_fire_47);
  assign mData_46 = xil_SimpleDualBram_46_doutb;
  assign xil_SimpleDualBram_47_addra = _zz_addra_47[10:0];
  assign xil_SimpleDualBram_47_addrb = _zz_addrb_47[13:0];
  assign sData_fire_48 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_47_ena = (_zz_ena_47[0] && sData_fire_48);
  assign mData_47 = xil_SimpleDualBram_47_doutb;
  assign xil_SimpleDualBram_48_addra = _zz_addra_48[10:0];
  assign xil_SimpleDualBram_48_addrb = _zz_addrb_48[13:0];
  assign sData_fire_49 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_48_ena = (_zz_ena_48[0] && sData_fire_49);
  assign mData_48 = xil_SimpleDualBram_48_doutb;
  assign xil_SimpleDualBram_49_addra = _zz_addra_49[10:0];
  assign xil_SimpleDualBram_49_addrb = _zz_addrb_49[13:0];
  assign sData_fire_50 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_49_ena = (_zz_ena_49[0] && sData_fire_50);
  assign mData_49 = xil_SimpleDualBram_49_doutb;
  assign xil_SimpleDualBram_50_addra = _zz_addra_50[10:0];
  assign xil_SimpleDualBram_50_addrb = _zz_addrb_50[13:0];
  assign sData_fire_51 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_50_ena = (_zz_ena_50[0] && sData_fire_51);
  assign mData_50 = xil_SimpleDualBram_50_doutb;
  assign xil_SimpleDualBram_51_addra = _zz_addra_51[10:0];
  assign xil_SimpleDualBram_51_addrb = _zz_addrb_51[13:0];
  assign sData_fire_52 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_51_ena = (_zz_ena_51[0] && sData_fire_52);
  assign mData_51 = xil_SimpleDualBram_51_doutb;
  assign xil_SimpleDualBram_52_addra = _zz_addra_52[10:0];
  assign xil_SimpleDualBram_52_addrb = _zz_addrb_52[13:0];
  assign sData_fire_53 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_52_ena = (_zz_ena_52[0] && sData_fire_53);
  assign mData_52 = xil_SimpleDualBram_52_doutb;
  assign xil_SimpleDualBram_53_addra = _zz_addra_53[10:0];
  assign xil_SimpleDualBram_53_addrb = _zz_addrb_53[13:0];
  assign sData_fire_54 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_53_ena = (_zz_ena_53[0] && sData_fire_54);
  assign mData_53 = xil_SimpleDualBram_53_doutb;
  assign xil_SimpleDualBram_54_addra = _zz_addra_54[10:0];
  assign xil_SimpleDualBram_54_addrb = _zz_addrb_54[13:0];
  assign sData_fire_55 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_54_ena = (_zz_ena_54[0] && sData_fire_55);
  assign mData_54 = xil_SimpleDualBram_54_doutb;
  assign xil_SimpleDualBram_55_addra = _zz_addra_55[10:0];
  assign xil_SimpleDualBram_55_addrb = _zz_addrb_55[13:0];
  assign sData_fire_56 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_55_ena = (_zz_ena_55[0] && sData_fire_56);
  assign mData_55 = xil_SimpleDualBram_55_doutb;
  assign xil_SimpleDualBram_56_addra = _zz_addra_56[10:0];
  assign xil_SimpleDualBram_56_addrb = _zz_addrb_56[13:0];
  assign sData_fire_57 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_56_ena = (_zz_ena_56[0] && sData_fire_57);
  assign mData_56 = xil_SimpleDualBram_56_doutb;
  assign xil_SimpleDualBram_57_addra = _zz_addra_57[10:0];
  assign xil_SimpleDualBram_57_addrb = _zz_addrb_57[13:0];
  assign sData_fire_58 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_57_ena = (_zz_ena_57[0] && sData_fire_58);
  assign mData_57 = xil_SimpleDualBram_57_doutb;
  assign xil_SimpleDualBram_58_addra = _zz_addra_58[10:0];
  assign xil_SimpleDualBram_58_addrb = _zz_addrb_58[13:0];
  assign sData_fire_59 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_58_ena = (_zz_ena_58[0] && sData_fire_59);
  assign mData_58 = xil_SimpleDualBram_58_doutb;
  assign xil_SimpleDualBram_59_addra = _zz_addra_59[10:0];
  assign xil_SimpleDualBram_59_addrb = _zz_addrb_59[13:0];
  assign sData_fire_60 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_59_ena = (_zz_ena_59[0] && sData_fire_60);
  assign mData_59 = xil_SimpleDualBram_59_doutb;
  assign xil_SimpleDualBram_60_addra = _zz_addra_60[10:0];
  assign xil_SimpleDualBram_60_addrb = _zz_addrb_60[13:0];
  assign sData_fire_61 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_60_ena = (_zz_ena_60[0] && sData_fire_61);
  assign mData_60 = xil_SimpleDualBram_60_doutb;
  assign xil_SimpleDualBram_61_addra = _zz_addra_61[10:0];
  assign xil_SimpleDualBram_61_addrb = _zz_addrb_61[13:0];
  assign sData_fire_62 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_61_ena = (_zz_ena_61[0] && sData_fire_62);
  assign mData_61 = xil_SimpleDualBram_61_doutb;
  assign xil_SimpleDualBram_62_addra = _zz_addra_62[10:0];
  assign xil_SimpleDualBram_62_addrb = _zz_addrb_62[13:0];
  assign sData_fire_63 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_62_ena = (_zz_ena_62[0] && sData_fire_63);
  assign mData_62 = xil_SimpleDualBram_62_doutb;
  assign xil_SimpleDualBram_63_addra = _zz_addra_63[10:0];
  assign xil_SimpleDualBram_63_addrb = _zz_addrb_63[13:0];
  assign sData_fire_64 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_63_ena = (_zz_ena_63[0] && sData_fire_64);
  assign mData_63 = xil_SimpleDualBram_63_doutb;
  assign sData_ready = ((Fsm_currentState & WEIGHT_CACHE_STATUS_CACHE_WEIGHT) != 4'b0000);
  assign Fsm_SA_Computed = LayerEnd;
  always @(*) begin
    case(OutCol_Cnt_count)
      16'h0001 : begin
        MatrixCol_Switch_1[0 : 0] = 1'b1;
        MatrixCol_Switch_1[7 : 1] = 7'h0;
      end
      16'h0002 : begin
        MatrixCol_Switch_1[1 : 0] = 2'b11;
        MatrixCol_Switch_1[7 : 2] = 6'h0;
      end
      16'h0003 : begin
        MatrixCol_Switch_1[2 : 0] = 3'b111;
        MatrixCol_Switch_1[7 : 3] = 5'h0;
      end
      16'h0004 : begin
        MatrixCol_Switch_1[3 : 0] = 4'b1111;
        MatrixCol_Switch_1[7 : 4] = 4'b0000;
      end
      16'h0005 : begin
        MatrixCol_Switch_1[4 : 0] = 5'h1f;
        MatrixCol_Switch_1[7 : 5] = 3'b000;
      end
      16'h0006 : begin
        MatrixCol_Switch_1[5 : 0] = 6'h3f;
        MatrixCol_Switch_1[7 : 6] = 2'b00;
      end
      16'h0007 : begin
        MatrixCol_Switch_1[6 : 0] = 7'h7f;
        MatrixCol_Switch_1[7 : 7] = 1'b0;
      end
      default : begin
        MatrixCol_Switch_1 = 8'hff;
      end
    endcase
  end

  assign MatrixCol_Switch = MatrixCol_Switch_1_regNext;
  always @(posedge clk) begin
    start_regNext <= start;
    MatrixCol_Switch_1_regNext <= MatrixCol_Switch_1;
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= WEIGHT_CACHE_STATUS_IDLE;
      Init_Count_count <= 3'b000;
      InData_Switch <= 64'h0000000000000001;
      In_Row_Cnt_count <= 16'h0;
      In_Col_Cnt_count <= 16'h0;
      Read_Row_Base_Addr <= 16'h0;
      Write_Row_Base_Addr <= 16'h0;
      OutRow_Cnt_count <= 16'h0;
      OutCol_Cnt_count <= Matrix_Col;
      Col_In_8_Cnt_count <= 6'h0;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l19) begin
        Init_Count_count <= (Init_Count_count + 3'b001);
        if(Init_Count_valid) begin
          Init_Count_count <= 3'b000;
        end
      end
      if(sData_fire) begin
        if(In_Row_Cnt_valid) begin
          In_Row_Cnt_count <= 16'h0;
        end else begin
          In_Row_Cnt_count <= (In_Row_Cnt_count + 16'h0001);
        end
      end
      if(In_Row_Cnt_valid) begin
        if(In_Col_Cnt_valid) begin
          In_Col_Cnt_count <= 16'h0;
        end else begin
          In_Col_Cnt_count <= (In_Col_Cnt_count + 16'h0001);
        end
      end
      if(when_WaCounter_l40) begin
        if(OutRow_Cnt_valid) begin
          OutRow_Cnt_count <= 16'h0;
        end else begin
          OutRow_Cnt_count <= (OutRow_Cnt_count + 16'h0001);
        end
      end
      if(OutRow_Cnt_valid) begin
        if(OutCol_Cnt_valid) begin
          OutCol_Cnt_count <= Matrix_Col;
        end else begin
          OutCol_Cnt_count <= (OutCol_Cnt_count - _zz_OutCol_Cnt_count_1);
        end
      end
      if(start) begin
        OutCol_Cnt_count <= Matrix_Col;
      end
      if(In_Row_Cnt_valid) begin
        if(Col_In_8_Cnt_valid) begin
          Col_In_8_Cnt_count <= 6'h0;
        end else begin
          Col_In_8_Cnt_count <= (Col_In_8_Cnt_count + 6'h01);
        end
      end
      if(OutCol_Cnt_valid) begin
        Col_In_8_Cnt_count <= 6'h0;
        Read_Row_Base_Addr <= 16'h0;
      end else begin
        if(OutRow_Cnt_valid) begin
          Read_Row_Base_Addr <= (Read_Row_Base_Addr + Matrix_Row);
        end
      end
      if(when_SA3D_WeightCache_l129) begin
        InData_Switch <= 64'h0000000000000001;
      end else begin
        if(In_Row_Cnt_valid) begin
          InData_Switch <= {InData_Switch[62 : 0],InData_Switch[63 : 63]};
        end
      end
      if(when_SA3D_WeightCache_l134) begin
        Write_Row_Base_Addr <= 16'h0;
      end else begin
        if(Col_In_8_Cnt_valid) begin
          Write_Row_Base_Addr <= (Write_Row_Base_Addr + _zz_Write_Row_Base_Addr);
        end
      end
    end
  end


endmodule
