// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : MyModule
// Git hash  : cbb23ce93bb580394fd976a943de961953f507e8

`timescale 1ns/1ps

module MyModule (
  output     [0:0]    io_PEZ_0_0,
  output     [0:0]    io_PEZ_0_1,
  output     [0:0]    io_PEZ_0_2,
  output     [0:0]    io_PEZ_0_3,
  output     [0:0]    io_PEZ_0_4,
  output     [0:0]    io_PEZ_0_5,
  output     [0:0]    io_PEZ_0_6,
  output     [0:0]    io_PEZ_0_7,
  output     [0:0]    io_PEZ_1_0,
  output     [0:0]    io_PEZ_1_1,
  output     [0:0]    io_PEZ_1_2,
  output     [0:0]    io_PEZ_1_3,
  output     [0:0]    io_PEZ_1_4,
  output     [0:0]    io_PEZ_1_5,
  output     [0:0]    io_PEZ_1_6,
  output     [0:0]    io_PEZ_1_7,
  output     [0:0]    io_PEZ_2_0,
  output     [0:0]    io_PEZ_2_1,
  output     [0:0]    io_PEZ_2_2,
  output     [0:0]    io_PEZ_2_3,
  output     [0:0]    io_PEZ_2_4,
  output     [0:0]    io_PEZ_2_5,
  output     [0:0]    io_PEZ_2_6,
  output     [0:0]    io_PEZ_2_7,
  output     [0:0]    io_PEZ_3_0,
  output     [0:0]    io_PEZ_3_1,
  output     [0:0]    io_PEZ_3_2,
  output     [0:0]    io_PEZ_3_3,
  output     [0:0]    io_PEZ_3_4,
  output     [0:0]    io_PEZ_3_5,
  output     [0:0]    io_PEZ_3_6,
  output     [0:0]    io_PEZ_3_7,
  output     [0:0]    io_PEZ_4_0,
  output     [0:0]    io_PEZ_4_1,
  output     [0:0]    io_PEZ_4_2,
  output     [0:0]    io_PEZ_4_3,
  output     [0:0]    io_PEZ_4_4,
  output     [0:0]    io_PEZ_4_5,
  output     [0:0]    io_PEZ_4_6,
  output     [0:0]    io_PEZ_4_7,
  output     [0:0]    io_PEZ_5_0,
  output     [0:0]    io_PEZ_5_1,
  output     [0:0]    io_PEZ_5_2,
  output     [0:0]    io_PEZ_5_3,
  output     [0:0]    io_PEZ_5_4,
  output     [0:0]    io_PEZ_5_5,
  output     [0:0]    io_PEZ_5_6,
  output     [0:0]    io_PEZ_5_7,
  output     [0:0]    io_PEZ_6_0,
  output     [0:0]    io_PEZ_6_1,
  output     [0:0]    io_PEZ_6_2,
  output     [0:0]    io_PEZ_6_3,
  output     [0:0]    io_PEZ_6_4,
  output     [0:0]    io_PEZ_6_5,
  output     [0:0]    io_PEZ_6_6,
  output     [0:0]    io_PEZ_6_7,
  output     [0:0]    io_PEZ_7_0,
  output     [0:0]    io_PEZ_7_1,
  output     [0:0]    io_PEZ_7_2,
  output     [0:0]    io_PEZ_7_3,
  output     [0:0]    io_PEZ_7_4,
  output     [0:0]    io_PEZ_7_5,
  output     [0:0]    io_PEZ_7_6,
  output     [0:0]    io_PEZ_7_7
);

  wire       [0:0]    vecArray_0_0;
  wire       [0:0]    vecArray_0_1;
  wire       [0:0]    vecArray_0_2;
  wire       [0:0]    vecArray_0_3;
  wire       [0:0]    vecArray_0_4;
  wire       [0:0]    vecArray_0_5;
  wire       [0:0]    vecArray_0_6;
  wire       [0:0]    vecArray_0_7;
  wire       [0:0]    vecArray_1_0;
  wire       [0:0]    vecArray_1_1;
  wire       [0:0]    vecArray_1_2;
  wire       [0:0]    vecArray_1_3;
  wire       [0:0]    vecArray_1_4;
  wire       [0:0]    vecArray_1_5;
  wire       [0:0]    vecArray_1_6;
  wire       [0:0]    vecArray_1_7;
  wire       [0:0]    vecArray_2_0;
  wire       [0:0]    vecArray_2_1;
  wire       [0:0]    vecArray_2_2;
  wire       [0:0]    vecArray_2_3;
  wire       [0:0]    vecArray_2_4;
  wire       [0:0]    vecArray_2_5;
  wire       [0:0]    vecArray_2_6;
  wire       [0:0]    vecArray_2_7;
  wire       [0:0]    vecArray_3_0;
  wire       [0:0]    vecArray_3_1;
  wire       [0:0]    vecArray_3_2;
  wire       [0:0]    vecArray_3_3;
  wire       [0:0]    vecArray_3_4;
  wire       [0:0]    vecArray_3_5;
  wire       [0:0]    vecArray_3_6;
  wire       [0:0]    vecArray_3_7;
  wire       [0:0]    vecArray_4_0;
  wire       [0:0]    vecArray_4_1;
  wire       [0:0]    vecArray_4_2;
  wire       [0:0]    vecArray_4_3;
  wire       [0:0]    vecArray_4_4;
  wire       [0:0]    vecArray_4_5;
  wire       [0:0]    vecArray_4_6;
  wire       [0:0]    vecArray_4_7;
  wire       [0:0]    vecArray_5_0;
  wire       [0:0]    vecArray_5_1;
  wire       [0:0]    vecArray_5_2;
  wire       [0:0]    vecArray_5_3;
  wire       [0:0]    vecArray_5_4;
  wire       [0:0]    vecArray_5_5;
  wire       [0:0]    vecArray_5_6;
  wire       [0:0]    vecArray_5_7;
  wire       [0:0]    vecArray_6_0;
  wire       [0:0]    vecArray_6_1;
  wire       [0:0]    vecArray_6_2;
  wire       [0:0]    vecArray_6_3;
  wire       [0:0]    vecArray_6_4;
  wire       [0:0]    vecArray_6_5;
  wire       [0:0]    vecArray_6_6;
  wire       [0:0]    vecArray_6_7;
  wire       [0:0]    vecArray_7_0;
  wire       [0:0]    vecArray_7_1;
  wire       [0:0]    vecArray_7_2;
  wire       [0:0]    vecArray_7_3;
  wire       [0:0]    vecArray_7_4;
  wire       [0:0]    vecArray_7_5;
  wire       [0:0]    vecArray_7_6;
  wire       [0:0]    vecArray_7_7;

  assign vecArray_0_0 = 1'b0;
  assign vecArray_0_1 = 1'b0;
  assign vecArray_0_2 = 1'b0;
  assign vecArray_0_3 = 1'b0;
  assign vecArray_0_4 = 1'b0;
  assign vecArray_0_5 = 1'b0;
  assign vecArray_0_6 = 1'b0;
  assign vecArray_0_7 = 1'b0;
  assign vecArray_1_0 = 1'b0;
  assign vecArray_1_1 = 1'b0;
  assign vecArray_1_2 = 1'b0;
  assign vecArray_1_3 = 1'b0;
  assign vecArray_1_4 = 1'b0;
  assign vecArray_1_5 = 1'b0;
  assign vecArray_1_6 = 1'b0;
  assign vecArray_1_7 = 1'b0;
  assign vecArray_2_0 = 1'b0;
  assign vecArray_2_1 = 1'b0;
  assign vecArray_2_2 = 1'b0;
  assign vecArray_2_3 = 1'b0;
  assign vecArray_2_4 = 1'b0;
  assign vecArray_2_5 = 1'b0;
  assign vecArray_2_6 = 1'b0;
  assign vecArray_2_7 = 1'b0;
  assign vecArray_3_0 = 1'b0;
  assign vecArray_3_1 = 1'b0;
  assign vecArray_3_2 = 1'b0;
  assign vecArray_3_3 = 1'b0;
  assign vecArray_3_4 = 1'b0;
  assign vecArray_3_5 = 1'b0;
  assign vecArray_3_6 = 1'b0;
  assign vecArray_3_7 = 1'b0;
  assign vecArray_4_0 = 1'b0;
  assign vecArray_4_1 = 1'b0;
  assign vecArray_4_2 = 1'b0;
  assign vecArray_4_3 = 1'b0;
  assign vecArray_4_4 = 1'b0;
  assign vecArray_4_5 = 1'b0;
  assign vecArray_4_6 = 1'b0;
  assign vecArray_4_7 = 1'b0;
  assign vecArray_5_0 = 1'b0;
  assign vecArray_5_1 = 1'b0;
  assign vecArray_5_2 = 1'b0;
  assign vecArray_5_3 = 1'b0;
  assign vecArray_5_4 = 1'b0;
  assign vecArray_5_5 = 1'b0;
  assign vecArray_5_6 = 1'b0;
  assign vecArray_5_7 = 1'b0;
  assign vecArray_6_0 = 1'b0;
  assign vecArray_6_1 = 1'b0;
  assign vecArray_6_2 = 1'b0;
  assign vecArray_6_3 = 1'b0;
  assign vecArray_6_4 = 1'b0;
  assign vecArray_6_5 = 1'b0;
  assign vecArray_6_6 = 1'b0;
  assign vecArray_6_7 = 1'b0;
  assign vecArray_7_0 = 1'b0;
  assign vecArray_7_1 = 1'b0;
  assign vecArray_7_2 = 1'b0;
  assign vecArray_7_3 = 1'b0;
  assign vecArray_7_4 = 1'b0;
  assign vecArray_7_5 = 1'b0;
  assign vecArray_7_6 = 1'b0;
  assign vecArray_7_7 = 1'b0;
  assign io_PEZ_0_0 = vecArray_0_0;
  assign io_PEZ_0_1 = vecArray_0_1;
  assign io_PEZ_0_2 = vecArray_0_2;
  assign io_PEZ_0_3 = vecArray_0_3;
  assign io_PEZ_0_4 = vecArray_0_4;
  assign io_PEZ_0_5 = vecArray_0_5;
  assign io_PEZ_0_6 = vecArray_0_6;
  assign io_PEZ_0_7 = vecArray_0_7;
  assign io_PEZ_1_0 = vecArray_1_0;
  assign io_PEZ_1_1 = vecArray_1_1;
  assign io_PEZ_1_2 = vecArray_1_2;
  assign io_PEZ_1_3 = vecArray_1_3;
  assign io_PEZ_1_4 = vecArray_1_4;
  assign io_PEZ_1_5 = vecArray_1_5;
  assign io_PEZ_1_6 = vecArray_1_6;
  assign io_PEZ_1_7 = vecArray_1_7;
  assign io_PEZ_2_0 = vecArray_2_0;
  assign io_PEZ_2_1 = vecArray_2_1;
  assign io_PEZ_2_2 = vecArray_2_2;
  assign io_PEZ_2_3 = vecArray_2_3;
  assign io_PEZ_2_4 = vecArray_2_4;
  assign io_PEZ_2_5 = vecArray_2_5;
  assign io_PEZ_2_6 = vecArray_2_6;
  assign io_PEZ_2_7 = vecArray_2_7;
  assign io_PEZ_3_0 = vecArray_3_0;
  assign io_PEZ_3_1 = vecArray_3_1;
  assign io_PEZ_3_2 = vecArray_3_2;
  assign io_PEZ_3_3 = vecArray_3_3;
  assign io_PEZ_3_4 = vecArray_3_4;
  assign io_PEZ_3_5 = vecArray_3_5;
  assign io_PEZ_3_6 = vecArray_3_6;
  assign io_PEZ_3_7 = vecArray_3_7;
  assign io_PEZ_4_0 = vecArray_4_0;
  assign io_PEZ_4_1 = vecArray_4_1;
  assign io_PEZ_4_2 = vecArray_4_2;
  assign io_PEZ_4_3 = vecArray_4_3;
  assign io_PEZ_4_4 = vecArray_4_4;
  assign io_PEZ_4_5 = vecArray_4_5;
  assign io_PEZ_4_6 = vecArray_4_6;
  assign io_PEZ_4_7 = vecArray_4_7;
  assign io_PEZ_5_0 = vecArray_5_0;
  assign io_PEZ_5_1 = vecArray_5_1;
  assign io_PEZ_5_2 = vecArray_5_2;
  assign io_PEZ_5_3 = vecArray_5_3;
  assign io_PEZ_5_4 = vecArray_5_4;
  assign io_PEZ_5_5 = vecArray_5_5;
  assign io_PEZ_5_6 = vecArray_5_6;
  assign io_PEZ_5_7 = vecArray_5_7;
  assign io_PEZ_6_0 = vecArray_6_0;
  assign io_PEZ_6_1 = vecArray_6_1;
  assign io_PEZ_6_2 = vecArray_6_2;
  assign io_PEZ_6_3 = vecArray_6_3;
  assign io_PEZ_6_4 = vecArray_6_4;
  assign io_PEZ_6_5 = vecArray_6_5;
  assign io_PEZ_6_6 = vecArray_6_6;
  assign io_PEZ_6_7 = vecArray_6_7;
  assign io_PEZ_7_0 = vecArray_7_0;
  assign io_PEZ_7_1 = vecArray_7_1;
  assign io_PEZ_7_2 = vecArray_7_2;
  assign io_PEZ_7_3 = vecArray_7_3;
  assign io_PEZ_7_4 = vecArray_7_4;
  assign io_PEZ_7_5 = vecArray_7_5;
  assign io_PEZ_7_6 = vecArray_7_6;
  assign io_PEZ_7_7 = vecArray_7_7;

endmodule
