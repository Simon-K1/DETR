// Generator : SpinalHDL v1.7.0    git head : eca519e78d4e6022e34911ec300a432ed9db8220
// Component : ConvOutput
// Git hash  : 33f9b9ad8900612c58d00d8143aee24055ba8f37

`timescale 1ns/1ps

module ConvOutput (
  input               sData_0_valid,
  output              sData_0_ready,
  input      [7:0]    sData_0_payload,
  input               sData_1_valid,
  output              sData_1_ready,
  input      [7:0]    sData_1_payload,
  input               sData_2_valid,
  output              sData_2_ready,
  input      [7:0]    sData_2_payload,
  input               sData_3_valid,
  output              sData_3_ready,
  input      [7:0]    sData_3_payload,
  input               sData_4_valid,
  output              sData_4_ready,
  input      [7:0]    sData_4_payload,
  input               sData_5_valid,
  output              sData_5_ready,
  input      [7:0]    sData_5_payload,
  input               sData_6_valid,
  output              sData_6_ready,
  input      [7:0]    sData_6_payload,
  input               sData_7_valid,
  output              sData_7_ready,
  input      [7:0]    sData_7_payload
);


  assign sData_0_ready = 1'b0;
  assign sData_1_ready = 1'b0;
  assign sData_2_ready = 1'b0;
  assign sData_3_ready = 1'b0;
  assign sData_4_ready = 1'b0;
  assign sData_5_ready = 1'b0;
  assign sData_6_ready = 1'b0;
  assign sData_7_ready = 1'b0;

endmodule
