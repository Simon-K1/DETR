// Generator : SpinalHDL v1.7.0    git head : eca519e78d4e6022e34911ec300a432ed9db8220
// Component : Img2ColStreamV2
// Git hash  : 3f47e2272714eaadc4903fce7d57faff55e9534d

`timescale 1ns/1ps

module Img2ColStreamV2 (
  output reg [63:0]   mData,
  input               mReady,
  output              mValid,
  input      [63:0]   s_axis_s2mm_tdata,
  input      [7:0]    s_axis_s2mm_tkeep,
  input               s_axis_s2mm_tlast,
  output              s_axis_s2mm_tready,
  input               s_axis_s2mm_tvalid,
  input               start,
  output              Raddr_Valid,
  output              LayerEnd,
  input               clk,
  input               reset
);

  wire       [15:0]   SubModule_Test_Generate_Period;
  wire                streamFifo_io_push_valid;
  wire                streamFifo_1_io_push_valid;
  wire                streamFifo_2_io_push_valid;
  wire                streamFifo_3_io_push_valid;
  wire                streamFifo_4_io_push_valid;
  wire                streamFifo_5_io_push_valid;
  wire                streamFifo_6_io_push_valid;
  wire                streamFifo_7_io_push_valid;
  wire                SubModule_sData_ready;
  wire       [63:0]   SubModule_mData;
  wire                SubModule_mValid;
  wire                SubModule_mLast;
  wire                SubModule_Test_Signal;
  wire                SubModule_Test_End;
  wire                SubModule_Raddr_Valid;
  wire                SubModule_LayerEnd;
  wire                streamFifo_io_push_ready;
  wire                streamFifo_io_pop_valid;
  wire       [63:0]   streamFifo_io_pop_payload;
  wire       [4:0]    streamFifo_io_occupancy;
  wire       [4:0]    streamFifo_io_availability;
  wire                axisDataConverter_8_inStream_ready;
  wire                axisDataConverter_8_outStream_valid;
  wire       [7:0]    axisDataConverter_8_outStream_payload;
  wire                streamFifo_1_io_push_ready;
  wire                streamFifo_1_io_pop_valid;
  wire       [63:0]   streamFifo_1_io_pop_payload;
  wire       [4:0]    streamFifo_1_io_occupancy;
  wire       [4:0]    streamFifo_1_io_availability;
  wire                axisDataConverter_9_inStream_ready;
  wire                axisDataConverter_9_outStream_valid;
  wire       [7:0]    axisDataConverter_9_outStream_payload;
  wire                streamFifo_2_io_push_ready;
  wire                streamFifo_2_io_pop_valid;
  wire       [63:0]   streamFifo_2_io_pop_payload;
  wire       [4:0]    streamFifo_2_io_occupancy;
  wire       [4:0]    streamFifo_2_io_availability;
  wire                axisDataConverter_10_inStream_ready;
  wire                axisDataConverter_10_outStream_valid;
  wire       [7:0]    axisDataConverter_10_outStream_payload;
  wire                streamFifo_3_io_push_ready;
  wire                streamFifo_3_io_pop_valid;
  wire       [63:0]   streamFifo_3_io_pop_payload;
  wire       [4:0]    streamFifo_3_io_occupancy;
  wire       [4:0]    streamFifo_3_io_availability;
  wire                axisDataConverter_11_inStream_ready;
  wire                axisDataConverter_11_outStream_valid;
  wire       [7:0]    axisDataConverter_11_outStream_payload;
  wire                streamFifo_4_io_push_ready;
  wire                streamFifo_4_io_pop_valid;
  wire       [63:0]   streamFifo_4_io_pop_payload;
  wire       [4:0]    streamFifo_4_io_occupancy;
  wire       [4:0]    streamFifo_4_io_availability;
  wire                axisDataConverter_12_inStream_ready;
  wire                axisDataConverter_12_outStream_valid;
  wire       [7:0]    axisDataConverter_12_outStream_payload;
  wire                streamFifo_5_io_push_ready;
  wire                streamFifo_5_io_pop_valid;
  wire       [63:0]   streamFifo_5_io_pop_payload;
  wire       [4:0]    streamFifo_5_io_occupancy;
  wire       [4:0]    streamFifo_5_io_availability;
  wire                axisDataConverter_13_inStream_ready;
  wire                axisDataConverter_13_outStream_valid;
  wire       [7:0]    axisDataConverter_13_outStream_payload;
  wire                streamFifo_6_io_push_ready;
  wire                streamFifo_6_io_pop_valid;
  wire       [63:0]   streamFifo_6_io_pop_payload;
  wire       [4:0]    streamFifo_6_io_occupancy;
  wire       [4:0]    streamFifo_6_io_availability;
  wire                axisDataConverter_14_inStream_ready;
  wire                axisDataConverter_14_outStream_valid;
  wire       [7:0]    axisDataConverter_14_outStream_payload;
  wire                streamFifo_7_io_push_ready;
  wire                streamFifo_7_io_pop_valid;
  wire       [63:0]   streamFifo_7_io_pop_payload;
  wire       [4:0]    streamFifo_7_io_occupancy;
  wire       [4:0]    streamFifo_7_io_availability;
  wire                axisDataConverter_15_inStream_ready;
  wire                axisDataConverter_15_outStream_valid;
  wire       [7:0]    axisDataConverter_15_outStream_payload;
  reg        [7:0]    OutData_Switch;
  wire                TestValid_Signal_0;
  wire                TestValid_Signal_1;
  wire                TestValid_Signal_2;
  wire                TestValid_Signal_3;
  wire                TestValid_Signal_4;
  wire                TestValid_Signal_5;
  wire                TestValid_Signal_6;
  wire                TestValid_Signal_7;
  reg        [7:0]    axisDataConverter_8_outStream_payload_regNext;
  reg        [7:0]    axisDataConverter_9_outStream_payload_regNext;
  reg        [7:0]    axisDataConverter_10_outStream_payload_regNext;
  reg        [7:0]    axisDataConverter_11_outStream_payload_regNext;
  reg        [7:0]    axisDataConverter_12_outStream_payload_regNext;
  reg        [7:0]    axisDataConverter_13_outStream_payload_regNext;
  reg        [7:0]    axisDataConverter_14_outStream_payload_regNext;
  reg        [7:0]    axisDataConverter_15_outStream_payload_regNext;
  reg                 axisDataConverter_8_outStream_valid_regNext;
  reg                 SubModule_LayerEnd_delay_1;
  reg                 SubModule_LayerEnd_delay_2;
  reg                 SubModule_LayerEnd_delay_3;
  wire                when_WaCounter_l18;
  reg        [31:0]   Out_Data_Counter_count;
  reg                 Out_Data_Counter_valid;
  wire                when_WaCounter_l13;
  wire                when_WaCounter_l18_1;
  reg        [31:0]   In_Data_Counter_count;
  reg                 In_Data_Counter_valid;
  wire                when_WaCounter_l13_1;

  Img2Col_Top SubModule (
    .start                          (start                               ), //i
    .sData_valid                    (s_axis_s2mm_tvalid                  ), //i
    .sData_ready                    (SubModule_sData_ready               ), //o
    .sData_payload                  (s_axis_s2mm_tdata[63:0]             ), //i
    .mData                          (SubModule_mData[63:0]               ), //o
    .mReady                         (streamFifo_io_push_ready            ), //i
    .mValid                         (SubModule_mValid                    ), //o
    .mLast                          (SubModule_mLast                     ), //o
    .Stride                         (5'h02                               ), //i
    .Kernel_Size                    (5'h04                               ), //i
    .Window_Size                    (16'h0010                            ), //i
    .InFeature_Size                 (16'h00e2                            ), //i
    .InFeature_Channel              (16'h0020                            ), //i
    .OutFeature_Channel             (16'h0020                            ), //i
    .OutFeature_Size                (16'h0070                            ), //i
    .OutCol_Count_Times             (16'h000e                            ), //i
    .InCol_Count_Times              (16'h0388                            ), //i
    .OutRow_Count_Times             (16'h0070                            ), //i
    .OutFeature_Channel_Count_Times (16'h0004                            ), //i
    .Test_Signal                    (SubModule_Test_Signal               ), //o
    .Test_Generate_Period           (SubModule_Test_Generate_Period[15:0]), //i
    .Test_End                       (SubModule_Test_End                  ), //o
    .Sliding_Size                   (13'h0008                            ), //i
    .Raddr_Valid                    (SubModule_Raddr_Valid               ), //o
    .LayerEnd                       (SubModule_LayerEnd                  ), //o
    .clk                            (clk                                 ), //i
    .reset                          (reset                               )  //i
  );
  WidthConverter_Fifo streamFifo (
    .io_push_valid   (streamFifo_io_push_valid          ), //i
    .io_push_ready   (streamFifo_io_push_ready          ), //o
    .io_push_payload (SubModule_mData[63:0]             ), //i
    .io_pop_valid    (streamFifo_io_pop_valid           ), //o
    .io_pop_ready    (axisDataConverter_8_inStream_ready), //i
    .io_pop_payload  (streamFifo_io_pop_payload[63:0]   ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (streamFifo_io_occupancy[4:0]      ), //o
    .io_availability (streamFifo_io_availability[4:0]   ), //o
    .clk             (clk                               ), //i
    .reset           (reset                             )  //i
  );
  AxisDataConverter axisDataConverter_8 (
    .inStream_valid    (streamFifo_io_pop_valid                   ), //i
    .inStream_ready    (axisDataConverter_8_inStream_ready        ), //o
    .inStream_payload  (streamFifo_io_pop_payload[63:0]           ), //i
    .outStream_valid   (axisDataConverter_8_outStream_valid       ), //o
    .outStream_ready   (1'b1                                      ), //i
    .outStream_payload (axisDataConverter_8_outStream_payload[7:0]), //o
    .clk               (clk                                       ), //i
    .reset             (reset                                     )  //i
  );
  WidthConverter_Fifo streamFifo_1 (
    .io_push_valid   (streamFifo_1_io_push_valid        ), //i
    .io_push_ready   (streamFifo_1_io_push_ready        ), //o
    .io_push_payload (SubModule_mData[63:0]             ), //i
    .io_pop_valid    (streamFifo_1_io_pop_valid         ), //o
    .io_pop_ready    (axisDataConverter_9_inStream_ready), //i
    .io_pop_payload  (streamFifo_1_io_pop_payload[63:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (streamFifo_1_io_occupancy[4:0]    ), //o
    .io_availability (streamFifo_1_io_availability[4:0] ), //o
    .clk             (clk                               ), //i
    .reset           (reset                             )  //i
  );
  AxisDataConverter axisDataConverter_9 (
    .inStream_valid    (streamFifo_1_io_pop_valid                 ), //i
    .inStream_ready    (axisDataConverter_9_inStream_ready        ), //o
    .inStream_payload  (streamFifo_1_io_pop_payload[63:0]         ), //i
    .outStream_valid   (axisDataConverter_9_outStream_valid       ), //o
    .outStream_ready   (1'b1                                      ), //i
    .outStream_payload (axisDataConverter_9_outStream_payload[7:0]), //o
    .clk               (clk                                       ), //i
    .reset             (reset                                     )  //i
  );
  WidthConverter_Fifo streamFifo_2 (
    .io_push_valid   (streamFifo_2_io_push_valid         ), //i
    .io_push_ready   (streamFifo_2_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_2_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_10_inStream_ready), //i
    .io_pop_payload  (streamFifo_2_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_2_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_2_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_10 (
    .inStream_valid    (streamFifo_2_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_10_inStream_ready        ), //o
    .inStream_payload  (streamFifo_2_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_10_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_10_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  WidthConverter_Fifo streamFifo_3 (
    .io_push_valid   (streamFifo_3_io_push_valid         ), //i
    .io_push_ready   (streamFifo_3_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_3_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_11_inStream_ready), //i
    .io_pop_payload  (streamFifo_3_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_3_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_3_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_11 (
    .inStream_valid    (streamFifo_3_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_11_inStream_ready        ), //o
    .inStream_payload  (streamFifo_3_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_11_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_11_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  WidthConverter_Fifo streamFifo_4 (
    .io_push_valid   (streamFifo_4_io_push_valid         ), //i
    .io_push_ready   (streamFifo_4_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_4_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_12_inStream_ready), //i
    .io_pop_payload  (streamFifo_4_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_4_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_4_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_12 (
    .inStream_valid    (streamFifo_4_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_12_inStream_ready        ), //o
    .inStream_payload  (streamFifo_4_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_12_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_12_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  WidthConverter_Fifo streamFifo_5 (
    .io_push_valid   (streamFifo_5_io_push_valid         ), //i
    .io_push_ready   (streamFifo_5_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_5_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_13_inStream_ready), //i
    .io_pop_payload  (streamFifo_5_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_5_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_5_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_13 (
    .inStream_valid    (streamFifo_5_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_13_inStream_ready        ), //o
    .inStream_payload  (streamFifo_5_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_13_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_13_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  WidthConverter_Fifo streamFifo_6 (
    .io_push_valid   (streamFifo_6_io_push_valid         ), //i
    .io_push_ready   (streamFifo_6_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_6_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_14_inStream_ready), //i
    .io_pop_payload  (streamFifo_6_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_6_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_6_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_14 (
    .inStream_valid    (streamFifo_6_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_14_inStream_ready        ), //o
    .inStream_payload  (streamFifo_6_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_14_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_14_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  WidthConverter_Fifo streamFifo_7 (
    .io_push_valid   (streamFifo_7_io_push_valid         ), //i
    .io_push_ready   (streamFifo_7_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_7_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_15_inStream_ready), //i
    .io_pop_payload  (streamFifo_7_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_7_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_7_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_15 (
    .inStream_valid    (streamFifo_7_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_15_inStream_ready        ), //o
    .inStream_payload  (streamFifo_7_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_15_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_15_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  assign streamFifo_io_push_valid = (OutData_Switch[0] && SubModule_mValid);
  always @(*) begin
    mData[7 : 0] = axisDataConverter_8_outStream_payload_regNext;
    mData[15 : 8] = axisDataConverter_9_outStream_payload_regNext;
    mData[23 : 16] = axisDataConverter_10_outStream_payload_regNext;
    mData[31 : 24] = axisDataConverter_11_outStream_payload_regNext;
    mData[39 : 32] = axisDataConverter_12_outStream_payload_regNext;
    mData[47 : 40] = axisDataConverter_13_outStream_payload_regNext;
    mData[55 : 48] = axisDataConverter_14_outStream_payload_regNext;
    mData[63 : 56] = axisDataConverter_15_outStream_payload_regNext;
  end

  assign streamFifo_1_io_push_valid = (OutData_Switch[1] && SubModule_mValid);
  assign streamFifo_2_io_push_valid = (OutData_Switch[2] && SubModule_mValid);
  assign streamFifo_3_io_push_valid = (OutData_Switch[3] && SubModule_mValid);
  assign streamFifo_4_io_push_valid = (OutData_Switch[4] && SubModule_mValid);
  assign streamFifo_5_io_push_valid = (OutData_Switch[5] && SubModule_mValid);
  assign streamFifo_6_io_push_valid = (OutData_Switch[6] && SubModule_mValid);
  assign streamFifo_7_io_push_valid = (OutData_Switch[7] && SubModule_mValid);
  assign mValid = axisDataConverter_8_outStream_valid_regNext;
  assign Raddr_Valid = axisDataConverter_8_outStream_valid;
  assign s_axis_s2mm_tready = SubModule_sData_ready;
  assign LayerEnd = SubModule_LayerEnd_delay_3;
  assign when_WaCounter_l18 = (mReady && mValid);
  assign when_WaCounter_l13 = (Out_Data_Counter_count == 32'hffffffff);
  always @(*) begin
    if(when_WaCounter_l13) begin
      Out_Data_Counter_valid = 1'b1;
    end else begin
      Out_Data_Counter_valid = 1'b0;
    end
    if(start) begin
      Out_Data_Counter_valid = 1'b0;
    end
  end

  assign when_WaCounter_l18_1 = (s_axis_s2mm_tvalid && s_axis_s2mm_tready);
  assign when_WaCounter_l13_1 = (In_Data_Counter_count == 32'hffffffff);
  always @(*) begin
    if(when_WaCounter_l13_1) begin
      In_Data_Counter_valid = 1'b1;
    end else begin
      In_Data_Counter_valid = 1'b0;
    end
    if(start) begin
      In_Data_Counter_valid = 1'b0;
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      OutData_Switch <= 8'h01;
      Out_Data_Counter_count <= 32'h0;
      In_Data_Counter_count <= 32'h0;
    end else begin
      if(SubModule_mValid) begin
        OutData_Switch <= {OutData_Switch[6 : 0],OutData_Switch[7 : 7]};
      end
      if(when_WaCounter_l18) begin
        Out_Data_Counter_count <= (Out_Data_Counter_count + 32'h00000001);
        if(Out_Data_Counter_valid) begin
          Out_Data_Counter_count <= 32'h0;
        end
      end
      if(when_WaCounter_l18_1) begin
        In_Data_Counter_count <= (In_Data_Counter_count + 32'h00000001);
        if(In_Data_Counter_valid) begin
          In_Data_Counter_count <= 32'h0;
        end
      end
      if(start) begin
        Out_Data_Counter_count <= 32'h0;
        In_Data_Counter_count <= 32'h0;
      end
    end
  end

  always @(posedge clk) begin
    axisDataConverter_8_outStream_payload_regNext <= axisDataConverter_8_outStream_payload;
    axisDataConverter_9_outStream_payload_regNext <= axisDataConverter_9_outStream_payload;
    axisDataConverter_10_outStream_payload_regNext <= axisDataConverter_10_outStream_payload;
    axisDataConverter_11_outStream_payload_regNext <= axisDataConverter_11_outStream_payload;
    axisDataConverter_12_outStream_payload_regNext <= axisDataConverter_12_outStream_payload;
    axisDataConverter_13_outStream_payload_regNext <= axisDataConverter_13_outStream_payload;
    axisDataConverter_14_outStream_payload_regNext <= axisDataConverter_14_outStream_payload;
    axisDataConverter_15_outStream_payload_regNext <= axisDataConverter_15_outStream_payload;
    axisDataConverter_8_outStream_valid_regNext <= axisDataConverter_8_outStream_valid;
    SubModule_LayerEnd_delay_1 <= SubModule_LayerEnd;
    SubModule_LayerEnd_delay_2 <= SubModule_LayerEnd_delay_1;
    SubModule_LayerEnd_delay_3 <= SubModule_LayerEnd_delay_2;
  end


endmodule

//AxisDataConverter replaced by AxisDataConverter

//WidthConverter_Fifo replaced by WidthConverter_Fifo

//AxisDataConverter replaced by AxisDataConverter

//WidthConverter_Fifo replaced by WidthConverter_Fifo

//AxisDataConverter replaced by AxisDataConverter

//WidthConverter_Fifo replaced by WidthConverter_Fifo

//AxisDataConverter replaced by AxisDataConverter

//WidthConverter_Fifo replaced by WidthConverter_Fifo

//AxisDataConverter replaced by AxisDataConverter

//WidthConverter_Fifo replaced by WidthConverter_Fifo

//AxisDataConverter replaced by AxisDataConverter

//WidthConverter_Fifo replaced by WidthConverter_Fifo

//AxisDataConverter replaced by AxisDataConverter

//WidthConverter_Fifo replaced by WidthConverter_Fifo

module AxisDataConverter (
  input               inStream_valid,
  output              inStream_ready,
  input      [63:0]   inStream_payload,
  output              outStream_valid,
  input               outStream_ready,
  output     [7:0]    outStream_payload,
  input               clk,
  input               reset
);

  wire       [2:0]    _zz__zz_inStream_ready_1;
  wire       [0:0]    _zz__zz_inStream_ready_1_1;
  wire       [63:0]   _zz__zz_outStream_payload;
  reg        [7:0]    _zz_outStream_payload_1;
  wire                outStream_fire;
  reg                 _zz_inStream_ready;
  reg        [2:0]    _zz_inStream_ready_1;
  reg        [2:0]    _zz_inStream_ready_2;
  wire                _zz_inStream_ready_3;
  wire       [63:0]   _zz_outStream_payload;

  assign _zz__zz_inStream_ready_1_1 = _zz_inStream_ready;
  assign _zz__zz_inStream_ready_1 = {2'd0, _zz__zz_inStream_ready_1_1};
  assign _zz__zz_outStream_payload = inStream_payload;
  always @(*) begin
    case(_zz_inStream_ready_2)
      3'b000 : _zz_outStream_payload_1 = _zz_outStream_payload[7 : 0];
      3'b001 : _zz_outStream_payload_1 = _zz_outStream_payload[15 : 8];
      3'b010 : _zz_outStream_payload_1 = _zz_outStream_payload[23 : 16];
      3'b011 : _zz_outStream_payload_1 = _zz_outStream_payload[31 : 24];
      3'b100 : _zz_outStream_payload_1 = _zz_outStream_payload[39 : 32];
      3'b101 : _zz_outStream_payload_1 = _zz_outStream_payload[47 : 40];
      3'b110 : _zz_outStream_payload_1 = _zz_outStream_payload[55 : 48];
      default : _zz_outStream_payload_1 = _zz_outStream_payload[63 : 56];
    endcase
  end

  assign outStream_fire = (outStream_valid && outStream_ready);
  always @(*) begin
    _zz_inStream_ready = 1'b0;
    if(outStream_fire) begin
      _zz_inStream_ready = 1'b1;
    end
  end

  assign _zz_inStream_ready_3 = (_zz_inStream_ready_2 == 3'b111);
  always @(*) begin
    _zz_inStream_ready_1 = (_zz_inStream_ready_2 + _zz__zz_inStream_ready_1);
    if(1'b0) begin
      _zz_inStream_ready_1 = 3'b000;
    end
  end

  assign outStream_valid = inStream_valid;
  assign _zz_outStream_payload = _zz__zz_outStream_payload;
  assign outStream_payload = _zz_outStream_payload_1;
  assign inStream_ready = (outStream_ready && _zz_inStream_ready_3);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _zz_inStream_ready_2 <= 3'b000;
    end else begin
      _zz_inStream_ready_2 <= _zz_inStream_ready_1;
    end
  end


endmodule

module WidthConverter_Fifo (
  input               io_push_valid,
  output              io_push_ready,
  input      [63:0]   io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [63:0]   io_pop_payload,
  input               io_flush,
  output     [4:0]    io_occupancy,
  output     [4:0]    io_availability,
  input               clk,
  input               reset
);

  reg        [63:0]   _zz_logic_ram_port0;
  wire       [3:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [3:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [63:0]   _zz_logic_ram_port_1;
  wire       [3:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [3:0]    logic_pushPtr_valueNext;
  reg        [3:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [3:0]    logic_popPtr_valueNext;
  reg        [3:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1021;
  wire       [3:0]    logic_ptrDif;
  reg [63:0] logic_ram [0:15];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {3'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {3'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  assign _zz_logic_ram_port_1 = io_push_payload;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 4'b1111);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 4'b0000;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 4'b1111);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 4'b0000;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1021 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_pushPtr_value <= 4'b0000;
      logic_popPtr_value <= 4'b0000;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1021) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module Img2Col_Top (
  input               start,
  input               sData_valid,
  output              sData_ready,
  input      [63:0]   sData_payload,
  output     [63:0]   mData,
  input               mReady,
  output              mValid,
  output              mLast,
  input      [4:0]    Stride,
  input      [4:0]    Kernel_Size,
  input      [15:0]   Window_Size,
  input      [15:0]   InFeature_Size,
  input      [15:0]   InFeature_Channel,
  input      [15:0]   OutFeature_Channel,
  input      [15:0]   OutFeature_Size,
  input      [15:0]   OutCol_Count_Times,
  input      [15:0]   InCol_Count_Times,
  input      [15:0]   OutRow_Count_Times,
  input      [15:0]   OutFeature_Channel_Count_Times,
  output              Test_Signal,
  input      [15:0]   Test_Generate_Period,
  output              Test_End,
  input      [12:0]   Sliding_Size,
  output              Raddr_Valid,
  output              LayerEnd,
  input               clk,
  input               reset
);
  localparam IMG2COL_ENUM_IDLE = 7'd1;
  localparam IMG2COL_ENUM_INIT = 7'd2;
  localparam IMG2COL_ENUM_INIT_ADDR = 7'd4;
  localparam IMG2COL_ENUM_DATA_CACHE = 7'd8;
  localparam IMG2COL_ENUM_WAIT_COMPUTE = 7'd16;
  localparam IMG2COL_ENUM_UPDATE_ADDR = 7'd32;
  localparam IMG2COL_ENUM_START_COMPUTE = 7'd64;

  reg                 AddrFifo_io_push_valid;
  reg                 AddrFifo_io_pop_ready;
  wire                AddrFifo_io_flush;
  reg                 RaddrFifo0_io_push_valid;
  reg        [15:0]   RaddrFifo0_io_push_payload;
  reg                 RaddrFifo0_io_pop_ready;
  wire                RaddrFifo0_io_flush;
  wire                Img2Col_SubModule_start;
  wire                Img2Col_SubModule_NewAddrIn_valid;
  wire       [14:0]   DGB_addra;
  wire       [14:0]   DGB_addrb;
  wire                AddrFifo_io_push_ready;
  wire                AddrFifo_io_pop_valid;
  wire       [15:0]   AddrFifo_io_pop_payload;
  wire       [5:0]    AddrFifo_io_occupancy;
  wire       [5:0]    AddrFifo_io_availability;
  wire                RaddrFifo0_io_push_ready;
  wire                RaddrFifo0_io_pop_valid;
  wire       [15:0]   RaddrFifo0_io_pop_payload;
  wire       [5:0]    RaddrFifo0_io_occupancy;
  wire       [5:0]    RaddrFifo0_io_availability;
  wire                Img2Col_SubModule_NewAddrIn_ready;
  wire                Img2Col_SubModule_SA_Idle;
  wire       [15:0]   Img2Col_SubModule_Raddr;
  wire                Img2Col_SubModule_Raddr_Valid;
  wire                Img2Col_SubModule_SA_End;
  wire                Img2Col_SubModule_AddrReceived;
  wire       [63:0]   DGB_doutb;
  wire       [4:0]    _zz_Addr_Init_Cnt_valid;
  wire       [4:0]    _zz_Addr_Init_Cnt_valid_1;
  wire       [15:0]   _zz_In_Col_Cnt_valid;
  wire       [4:0]    _zz_Row_Cache_Cnt_valid;
  wire       [15:0]   _zz_In_Row_Cnt_valid;
  wire       [15:0]   _zz_when_Data_Generate_V2_l183;
  wire       [4:0]    _zz_when_Data_Generate_V2_l183_1;
  wire       [15:0]   _zz_Out_Row_Cnt_valid;
  wire       [15:0]   _zz_Test_Valid;
  reg                 start_regNext;
  wire                when_Data_Generate_V2_l35;
  reg        [6:0]    Fsm_currentState;
  reg        [6:0]    Fsm_nextState;
  wire                Fsm_Init_End;
  wire                Fsm_Addr_Inited;
  wire                Fsm_Data_Cached;
  wire                Fsm_Addr_Updated;
  wire                Fsm_SA_Ready;
  wire                Fsm_Cache_End;
  wire                Fsm_Layer_End;
  wire                when_Data_Generate_V2_l56;
  wire                when_WaCounter_l18;
  reg        [2:0]    Init_Count_count;
  reg                 Init_Count_valid;
  wire                when_WaCounter_l13;
  wire                when_WaCounter_l37;
  reg        [4:0]    Addr_Init_Cnt_count;
  wire                Addr_Init_Cnt_valid;
  reg        [15:0]   WaddrOffset;
  wire                when_Data_Generate_V2_l138;
  wire                AddrFifo_io_pop_fire;
  wire                when_Data_Generate_V2_l145;
  wire                when_Data_Generate_V2_l149;
  reg        [15:0]   Raddr_Initialization;
  wire                when_Data_Generate_V2_l159;
  wire                when_Data_Generate_V2_l163;
  reg        [4:0]    Cache_Row_Num;
  reg        [4:0]    Raddr_Updata_Cnt_Num;
  wire                sData_fire;
  reg        [15:0]   In_Col_Cnt_count;
  wire                In_Col_Cnt_valid;
  reg        [4:0]    Row_Cache_Cnt_count;
  wire                Row_Cache_Cnt_valid;
  reg        [15:0]   In_Row_Cnt_count;
  wire                In_Row_Cnt_valid;
  wire                when_Data_Generate_V2_l183;
  reg                 CacheEnd_Flag;
  wire                when_Data_Generate_V2_l194;
  wire                Img2ColOutput_Module_Ready_Receive_Addr;
  wire                when_Data_Generate_V2_l211;
  wire                RaddrFifo0_io_pop_fire;
  reg        [15:0]   Out_Row_Cnt_count;
  wire                Out_Row_Cnt_valid;
  wire       [15:0]   Waddr;
  wire                sData_fire_1;
  reg                 Img2Col_SubModule_Raddr_Valid_regNext;
  reg                 Out_Row_Cnt_valid_regNext;
  reg        [15:0]   Out_Row_Cnt_count_regNext;
  wire                Test_Valid;
  reg                 Test_Valid_regNext;
  `ifndef SYNTHESIS
  reg [103:0] Fsm_currentState_string;
  reg [103:0] Fsm_nextState_string;
  `endif


  assign _zz_Addr_Init_Cnt_valid = (_zz_Addr_Init_Cnt_valid_1 - 5'h01);
  assign _zz_Addr_Init_Cnt_valid_1 = (Kernel_Size + Stride);
  assign _zz_In_Col_Cnt_valid = (InCol_Count_Times - 16'h0001);
  assign _zz_Row_Cache_Cnt_valid = (Cache_Row_Num - 5'h01);
  assign _zz_In_Row_Cnt_valid = (InFeature_Size - 16'h0001);
  assign _zz_when_Data_Generate_V2_l183_1 = (Kernel_Size - 5'h01);
  assign _zz_when_Data_Generate_V2_l183 = {11'd0, _zz_when_Data_Generate_V2_l183_1};
  assign _zz_Out_Row_Cnt_valid = (OutRow_Count_Times - 16'h0001);
  assign _zz_Test_Valid = (Test_Generate_Period - 16'h0001);
  WaddrOffset_Fifo AddrFifo (
    .io_push_valid   (AddrFifo_io_push_valid       ), //i
    .io_push_ready   (AddrFifo_io_push_ready       ), //o
    .io_push_payload (WaddrOffset[15:0]            ), //i
    .io_pop_valid    (AddrFifo_io_pop_valid        ), //o
    .io_pop_ready    (AddrFifo_io_pop_ready        ), //i
    .io_pop_payload  (AddrFifo_io_pop_payload[15:0]), //o
    .io_flush        (AddrFifo_io_flush            ), //i
    .io_occupancy    (AddrFifo_io_occupancy[5:0]   ), //o
    .io_availability (AddrFifo_io_availability[5:0]), //o
    .clk             (clk                          ), //i
    .reset           (reset                        )  //i
  );
  WaddrOffset_Fifo RaddrFifo0 (
    .io_push_valid   (RaddrFifo0_io_push_valid        ), //i
    .io_push_ready   (RaddrFifo0_io_push_ready        ), //o
    .io_push_payload (RaddrFifo0_io_push_payload[15:0]), //i
    .io_pop_valid    (RaddrFifo0_io_pop_valid         ), //o
    .io_pop_ready    (RaddrFifo0_io_pop_ready         ), //i
    .io_pop_payload  (RaddrFifo0_io_pop_payload[15:0] ), //o
    .io_flush        (RaddrFifo0_io_flush             ), //i
    .io_occupancy    (RaddrFifo0_io_occupancy[5:0]    ), //o
    .io_availability (RaddrFifo0_io_availability[5:0] ), //o
    .clk             (clk                             ), //i
    .reset           (reset                           )  //i
  );
  Img2Col_OutPut Img2Col_SubModule (
    .start                          (Img2Col_SubModule_start             ), //i
    .NewAddrIn_valid                (Img2Col_SubModule_NewAddrIn_valid   ), //i
    .NewAddrIn_ready                (Img2Col_SubModule_NewAddrIn_ready   ), //o
    .NewAddrIn_payload              (RaddrFifo0_io_pop_payload[15:0]     ), //i
    .SA_Idle                        (Img2Col_SubModule_SA_Idle           ), //o
    .Raddr                          (Img2Col_SubModule_Raddr[15:0]       ), //o
    .Raddr_Valid                    (Img2Col_SubModule_Raddr_Valid       ), //o
    .SA_End                         (Img2Col_SubModule_SA_End            ), //o
    .Stride                         (Stride[4:0]                         ), //i
    .Kernel_Size                    (Kernel_Size[4:0]                    ), //i
    .Window_Size                    (Window_Size[15:0]                   ), //i
    .InFeature_Size                 (InFeature_Size[15:0]                ), //i
    .InFeature_Channel              (InFeature_Channel[15:0]             ), //i
    .OutFeature_Channel             (OutFeature_Channel[15:0]            ), //i
    .OutFeature_Size                (OutFeature_Size[15:0]               ), //i
    .OutCol_Count_Times             (OutCol_Count_Times[15:0]            ), //i
    .InCol_Count_Times              (InCol_Count_Times[15:0]             ), //i
    .OutFeature_Channel_Count_Times (OutFeature_Channel_Count_Times[15:0]), //i
    .Sliding_Size                   (Sliding_Size[12:0]                  ), //i
    .mReady                         (mReady                              ), //i
    .AddrReceived                   (Img2Col_SubModule_AddrReceived      ), //o
    .LayerEnd                       (Fsm_Layer_End                       ), //i
    .clk                            (clk                                 ), //i
    .reset                          (reset                               )  //i
  );
  DataGen_Bram DGB (
    .clka  (clk                ), //i
    .addra (DGB_addra[14:0]    ), //i
    .dina  (sData_payload[63:0]), //i
    .ena   (sData_fire_1       ), //i
    .wea   (1'b1               ), //i
    .addrb (DGB_addrb[14:0]    ), //i
    .doutb (DGB_doutb[63:0]    ), //o
    .clkb  (clk                )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      IMG2COL_ENUM_IDLE : Fsm_currentState_string = "IDLE         ";
      IMG2COL_ENUM_INIT : Fsm_currentState_string = "INIT         ";
      IMG2COL_ENUM_INIT_ADDR : Fsm_currentState_string = "INIT_ADDR    ";
      IMG2COL_ENUM_DATA_CACHE : Fsm_currentState_string = "DATA_CACHE   ";
      IMG2COL_ENUM_WAIT_COMPUTE : Fsm_currentState_string = "WAIT_COMPUTE ";
      IMG2COL_ENUM_UPDATE_ADDR : Fsm_currentState_string = "UPDATE_ADDR  ";
      IMG2COL_ENUM_START_COMPUTE : Fsm_currentState_string = "START_COMPUTE";
      default : Fsm_currentState_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      IMG2COL_ENUM_IDLE : Fsm_nextState_string = "IDLE         ";
      IMG2COL_ENUM_INIT : Fsm_nextState_string = "INIT         ";
      IMG2COL_ENUM_INIT_ADDR : Fsm_nextState_string = "INIT_ADDR    ";
      IMG2COL_ENUM_DATA_CACHE : Fsm_nextState_string = "DATA_CACHE   ";
      IMG2COL_ENUM_WAIT_COMPUTE : Fsm_nextState_string = "WAIT_COMPUTE ";
      IMG2COL_ENUM_UPDATE_ADDR : Fsm_nextState_string = "UPDATE_ADDR  ";
      IMG2COL_ENUM_START_COMPUTE : Fsm_nextState_string = "START_COMPUTE";
      default : Fsm_nextState_string = "?????????????";
    endcase
  end
  `endif

  assign when_Data_Generate_V2_l35 = (start && (! start_regNext));
  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & IMG2COL_ENUM_IDLE) == IMG2COL_ENUM_IDLE) : begin
        if(when_Data_Generate_V2_l35) begin
          Fsm_nextState = IMG2COL_ENUM_INIT;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_IDLE;
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_INIT) == IMG2COL_ENUM_INIT) : begin
        if(Fsm_Init_End) begin
          Fsm_nextState = IMG2COL_ENUM_INIT_ADDR;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_INIT;
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_INIT_ADDR) == IMG2COL_ENUM_INIT_ADDR) : begin
        if(Fsm_Addr_Inited) begin
          Fsm_nextState = IMG2COL_ENUM_DATA_CACHE;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_INIT_ADDR;
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_DATA_CACHE) == IMG2COL_ENUM_DATA_CACHE) : begin
        if(when_Data_Generate_V2_l56) begin
          Fsm_nextState = IMG2COL_ENUM_WAIT_COMPUTE;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_DATA_CACHE;
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_WAIT_COMPUTE) == IMG2COL_ENUM_WAIT_COMPUTE) : begin
        if(Fsm_Layer_End) begin
          Fsm_nextState = IMG2COL_ENUM_IDLE;
        end else begin
          if(Fsm_SA_Ready) begin
            Fsm_nextState = IMG2COL_ENUM_UPDATE_ADDR;
          end else begin
            Fsm_nextState = IMG2COL_ENUM_WAIT_COMPUTE;
          end
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_UPDATE_ADDR) == IMG2COL_ENUM_UPDATE_ADDR) : begin
        if(Fsm_Addr_Updated) begin
          Fsm_nextState = IMG2COL_ENUM_START_COMPUTE;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_UPDATE_ADDR;
        end
      end
      default : begin
        if(Fsm_Layer_End) begin
          Fsm_nextState = IMG2COL_ENUM_IDLE;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_DATA_CACHE;
        end
      end
    endcase
  end

  assign when_Data_Generate_V2_l56 = (Fsm_Data_Cached || Fsm_Cache_End);
  assign when_WaCounter_l18 = ((Fsm_currentState & IMG2COL_ENUM_INIT) != 7'b0000000);
  assign when_WaCounter_l13 = (Init_Count_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l13) begin
      Init_Count_valid = 1'b1;
    end else begin
      Init_Count_valid = 1'b0;
    end
  end

  assign Fsm_Init_End = Init_Count_valid;
  assign when_WaCounter_l37 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign Addr_Init_Cnt_valid = ((Addr_Init_Cnt_count == _zz_Addr_Init_Cnt_valid) && when_WaCounter_l37);
  assign Fsm_Addr_Inited = Addr_Init_Cnt_valid;
  always @(*) begin
    AddrFifo_io_push_valid = 1'b0;
    if(when_Data_Generate_V2_l138) begin
      AddrFifo_io_push_valid = 1'b1;
    end
    if(In_Col_Cnt_valid) begin
      AddrFifo_io_push_valid = 1'b1;
    end
  end

  always @(*) begin
    AddrFifo_io_pop_ready = 1'b0;
    if(when_Data_Generate_V2_l149) begin
      AddrFifo_io_pop_ready = 1'b1;
    end
    if(In_Col_Cnt_valid) begin
      AddrFifo_io_pop_ready = 1'b1;
    end
  end

  assign when_Data_Generate_V2_l138 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign AddrFifo_io_pop_fire = (AddrFifo_io_pop_valid && AddrFifo_io_pop_ready);
  assign when_Data_Generate_V2_l145 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign when_Data_Generate_V2_l149 = (((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000) && ((Fsm_nextState & IMG2COL_ENUM_DATA_CACHE) != 7'b0000000));
  always @(*) begin
    RaddrFifo0_io_push_valid = 1'b0;
    if(when_Data_Generate_V2_l159) begin
      RaddrFifo0_io_push_valid = 1'b1;
    end
    if(when_Data_Generate_V2_l211) begin
      RaddrFifo0_io_push_valid = RaddrFifo0_io_pop_fire;
    end
  end

  always @(*) begin
    RaddrFifo0_io_pop_ready = 1'b0;
    if(when_Data_Generate_V2_l211) begin
      RaddrFifo0_io_pop_ready = Img2ColOutput_Module_Ready_Receive_Addr;
    end
  end

  always @(*) begin
    RaddrFifo0_io_push_payload = RaddrFifo0_io_pop_payload;
    if(when_Data_Generate_V2_l159) begin
      RaddrFifo0_io_push_payload = Raddr_Initialization;
    end
    if(when_Data_Generate_V2_l211) begin
      RaddrFifo0_io_push_payload = RaddrFifo0_io_pop_payload;
    end
  end

  assign when_Data_Generate_V2_l159 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign when_Data_Generate_V2_l163 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign sData_fire = (sData_valid && sData_ready);
  assign In_Col_Cnt_valid = ((In_Col_Cnt_count == _zz_In_Col_Cnt_valid) && sData_fire);
  assign Row_Cache_Cnt_valid = ((Row_Cache_Cnt_count == _zz_Row_Cache_Cnt_valid) && In_Col_Cnt_valid);
  assign In_Row_Cnt_valid = ((In_Row_Cnt_count == _zz_In_Row_Cnt_valid) && In_Col_Cnt_valid);
  assign when_Data_Generate_V2_l183 = (_zz_when_Data_Generate_V2_l183 < In_Row_Cnt_count);
  always @(*) begin
    if(when_Data_Generate_V2_l183) begin
      Cache_Row_Num = Stride;
    end else begin
      Cache_Row_Num = Kernel_Size;
    end
  end

  always @(*) begin
    if(when_Data_Generate_V2_l183) begin
      Raddr_Updata_Cnt_Num = Stride;
    end else begin
      Raddr_Updata_Cnt_Num = Kernel_Size;
    end
  end

  assign Fsm_Data_Cached = Row_Cache_Cnt_valid;
  assign when_Data_Generate_V2_l194 = ((Fsm_currentState & IMG2COL_ENUM_IDLE) != 7'b0000000);
  assign Fsm_Cache_End = CacheEnd_Flag;
  assign sData_ready = ((Fsm_currentState & IMG2COL_ENUM_DATA_CACHE) != 7'b0000000);
  assign when_Data_Generate_V2_l211 = ((Fsm_currentState & IMG2COL_ENUM_UPDATE_ADDR) != 7'b0000000);
  assign RaddrFifo0_io_pop_fire = (RaddrFifo0_io_pop_valid && RaddrFifo0_io_pop_ready);
  assign Img2Col_SubModule_start = ((Fsm_currentState & IMG2COL_ENUM_UPDATE_ADDR) != 7'b0000000);
  assign Fsm_SA_Ready = Img2Col_SubModule_SA_Idle;
  assign Img2ColOutput_Module_Ready_Receive_Addr = Img2Col_SubModule_NewAddrIn_ready;
  assign Img2Col_SubModule_NewAddrIn_valid = ((Fsm_currentState & IMG2COL_ENUM_UPDATE_ADDR) != 7'b0000000);
  assign LayerEnd = Fsm_Layer_End;
  assign Fsm_Addr_Updated = Img2Col_SubModule_AddrReceived;
  assign Out_Row_Cnt_valid = ((Out_Row_Cnt_count == _zz_Out_Row_Cnt_valid) && Img2Col_SubModule_SA_End);
  assign Fsm_Layer_End = Out_Row_Cnt_valid;
  assign Waddr = (WaddrOffset + In_Col_Cnt_count);
  assign DGB_addra = Waddr[14:0];
  assign sData_fire_1 = (sData_valid && sData_ready);
  assign DGB_addrb = Img2Col_SubModule_Raddr[14:0];
  assign mData = DGB_doutb;
  assign mValid = Img2Col_SubModule_Raddr_Valid_regNext;
  assign mLast = Out_Row_Cnt_valid_regNext;
  assign Test_Valid = (_zz_Test_Valid == Out_Row_Cnt_count_regNext);
  assign Test_Signal = Test_Valid;
  assign Test_End = ((! Test_Valid) && Test_Valid_regNext);
  assign AddrFifo_io_flush = ((Fsm_nextState & IMG2COL_ENUM_IDLE) != 7'b0000000);
  assign RaddrFifo0_io_flush = ((Fsm_nextState & IMG2COL_ENUM_IDLE) != 7'b0000000);
  assign Raddr_Valid = Img2Col_SubModule_Raddr_Valid;
  always @(posedge clk) begin
    start_regNext <= start;
    Img2Col_SubModule_Raddr_Valid_regNext <= Img2Col_SubModule_Raddr_Valid;
    Out_Row_Cnt_valid_regNext <= Out_Row_Cnt_valid;
    Out_Row_Cnt_count_regNext <= Out_Row_Cnt_count;
    Test_Valid_regNext <= Test_Valid;
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= IMG2COL_ENUM_IDLE;
      Init_Count_count <= 3'b000;
      Addr_Init_Cnt_count <= 5'h0;
      WaddrOffset <= 16'h0;
      Raddr_Initialization <= 16'h0;
      In_Col_Cnt_count <= 16'h0;
      Row_Cache_Cnt_count <= 5'h0;
      In_Row_Cnt_count <= 16'h0;
      CacheEnd_Flag <= 1'b0;
      Out_Row_Cnt_count <= 16'h0;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l18) begin
        Init_Count_count <= (Init_Count_count + 3'b001);
        if(Init_Count_valid) begin
          Init_Count_count <= 3'b000;
        end
      end
      if(when_WaCounter_l37) begin
        if(Addr_Init_Cnt_valid) begin
          Addr_Init_Cnt_count <= 5'h0;
        end else begin
          Addr_Init_Cnt_count <= (Addr_Init_Cnt_count + 5'h01);
        end
      end
      if(AddrFifo_io_pop_fire) begin
        WaddrOffset <= AddrFifo_io_pop_payload;
      end else begin
        if(when_Data_Generate_V2_l145) begin
          WaddrOffset <= (WaddrOffset + InCol_Count_Times);
        end
      end
      if(when_Data_Generate_V2_l163) begin
        Raddr_Initialization <= (Raddr_Initialization + InCol_Count_Times);
      end else begin
        Raddr_Initialization <= 16'h0;
      end
      if(sData_fire) begin
        if(In_Col_Cnt_valid) begin
          In_Col_Cnt_count <= 16'h0;
        end else begin
          In_Col_Cnt_count <= (In_Col_Cnt_count + 16'h0001);
        end
      end
      if(In_Col_Cnt_valid) begin
        if(Row_Cache_Cnt_valid) begin
          Row_Cache_Cnt_count <= 5'h0;
        end else begin
          Row_Cache_Cnt_count <= (Row_Cache_Cnt_count + 5'h01);
        end
      end
      if(In_Col_Cnt_valid) begin
        if(In_Row_Cnt_valid) begin
          In_Row_Cnt_count <= 16'h0;
        end else begin
          In_Row_Cnt_count <= (In_Row_Cnt_count + 16'h0001);
        end
      end
      if(In_Row_Cnt_valid) begin
        CacheEnd_Flag <= 1'b1;
      end else begin
        if(when_Data_Generate_V2_l194) begin
          CacheEnd_Flag <= 1'b0;
        end
      end
      if(Img2Col_SubModule_SA_End) begin
        if(Out_Row_Cnt_valid) begin
          Out_Row_Cnt_count <= 16'h0;
        end else begin
          Out_Row_Cnt_count <= (Out_Row_Cnt_count + 16'h0001);
        end
      end
    end
  end


endmodule

module Img2Col_OutPut (
  input               start,
  input               NewAddrIn_valid,
  output              NewAddrIn_ready,
  input      [15:0]   NewAddrIn_payload,
  output              SA_Idle,
  output     [15:0]   Raddr,
  output              Raddr_Valid,
  output              SA_End,
  input      [4:0]    Stride,
  input      [4:0]    Kernel_Size,
  input      [15:0]   Window_Size,
  input      [15:0]   InFeature_Size,
  input      [15:0]   InFeature_Channel,
  input      [15:0]   OutFeature_Channel,
  input      [15:0]   OutFeature_Size,
  input      [15:0]   OutCol_Count_Times,
  input      [15:0]   InCol_Count_Times,
  input      [15:0]   OutFeature_Channel_Count_Times,
  input      [12:0]   Sliding_Size,
  input               mReady,
  output reg          AddrReceived,
  input               LayerEnd,
  input               clk,
  input               reset
);
  localparam IMG2COL_OUTPUT_ENUM_IDLE = 6'd1;
  localparam IMG2COL_OUTPUT_ENUM_INIT = 6'd2;
  localparam IMG2COL_OUTPUT_ENUM_INIT_ADDR = 6'd4;
  localparam IMG2COL_OUTPUT_ENUM_SA_COMPUTE = 6'd8;
  localparam IMG2COL_OUTPUT_ENUM_UPDATE_ADDR = 6'd16;
  localparam IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY = 6'd32;

  reg                 RaddrFifo1_io_push_valid;
  reg        [15:0]   RaddrFifo1_io_push_payload;
  reg                 RaddrFifo1_io_pop_ready;
  wire                RaddrFifo1_io_flush;
  wire                RaddrFifo1_io_push_ready;
  wire                RaddrFifo1_io_pop_valid;
  wire       [15:0]   RaddrFifo1_io_pop_payload;
  wire       [5:0]    RaddrFifo1_io_occupancy;
  wire       [5:0]    RaddrFifo1_io_availability;
  wire       [4:0]    _zz_Raddr_Init_Cnt_valid;
  wire       [4:0]    _zz_Raddr_Update_Cnt_valid;
  wire       [12:0]   _zz_In_Channel_Process_Cnt_valid;
  wire       [12:0]   _zz_In_Channel_Process_Cnt_valid_1;
  wire       [15:0]   _zz_Window_Col_Cnt_valid;
  wire       [4:0]    _zz_Window_Col_Cnt_valid_1;
  wire       [15:0]   _zz_Window_Row_Cnt_valid;
  wire       [4:0]    _zz_Window_Row_Cnt_valid_1;
  wire       [15:0]   _zz_Out_Channel_Cnt_valid;
  wire       [15:0]   _zz_Out_Col_Cnt_valid;
  wire       [15:0]   _zz_when_Data_Generate_V2_l446;
  wire       [15:0]   _zz_when_Data_Generate_V2_l446_1;
  wire       [15:0]   _zz_WindowSize_Cnt_valid;
  wire       [15:0]   _zz_WindowSize_Cnt_valid_1;
  wire       [31:0]   _zz_Kernel_Base_Addr;
  wire       [15:0]   _zz_Kernel_Base_Addr_1;
  wire       [31:0]   _zz_Kernel_Addr;
  wire       [15:0]   _zz_Kernel_Addr_1;
  wire       [31:0]   _zz_Kernel_Addr_2;
  wire       [31:0]   _zz_Kernel_Addr_3;
  wire       [31:0]   _zz_Kernel_Addr_4;
  wire       [31:0]   _zz_Raddr;
  wire       [31:0]   _zz_Raddr_1;
  reg                 start_regNext;
  wire                when_Data_Generate_V2_l303;
  reg        [5:0]    Fsm_currentState;
  reg        [5:0]    Fsm_nextState;
  wire                Fsm_Init_End;
  wire                Fsm_Addr_Inited;
  wire                Fsm_SA_Computed;
  wire                Fsm_Addr_Updated;
  wire                Fsm_LayerEnd;
  wire                Fsm_NextReady;
  wire                when_Data_Generate_V2_l335;
  wire                when_WaCounter_l18;
  reg        [2:0]    Init_Count_count;
  reg                 Init_Count_valid;
  wire                when_WaCounter_l13;
  reg        [15:0]   Row_Base_Addr;
  wire                RaddrFifo1_io_pop_fire;
  wire                RaddrFifo1_io_push_fire;
  wire                when_WaCounter_l37;
  reg        [4:0]    Raddr_Init_Cnt_count;
  wire                Raddr_Init_Cnt_valid;
  wire                RaddrFifo1_io_push_fire_1;
  wire                when_WaCounter_l37_1;
  reg        [4:0]    Raddr_Update_Cnt_count;
  wire                Raddr_Update_Cnt_valid;
  wire                when_Data_Generate_V2_l412;
  wire                when_WaCounter_l37_2;
  reg        [2:0]    SA_Row_Cnt_count;
  reg                 SA_Row_Cnt_valid;
  reg        [12:0]   In_Channel_Process_Cnt_count;
  wire                In_Channel_Process_Cnt_valid;
  reg        [15:0]   Window_Col_Cnt_count;
  wire                Window_Col_Cnt_valid;
  reg        [15:0]   Window_Row_Cnt_count;
  wire                Window_Row_Cnt_valid;
  reg        [15:0]   Out_Channel_Cnt_count;
  wire                Out_Channel_Cnt_valid;
  reg        [15:0]   Out_Col_Cnt_count;
  wire                Out_Col_Cnt_valid;
  reg        [15:0]   OutFeature_Col_Lefted;
  wire                when_Data_Generate_V2_l443;
  wire                when_Data_Generate_V2_l446;
  reg        [12:0]   WindowSize_Cnt_count;
  wire                WindowSize_Cnt_valid;
  reg        [31:0]   Kernel_Addr;
  reg        [31:0]   Kernel_Base_Addr;
  wire                when_Data_Generate_V2_l471;
  wire                when_Data_Generate_V2_l481;
  wire                RaddrFifo1_io_push_fire_2;
  wire                when_Data_Generate_V2_l485;
  `ifndef SYNTHESIS
  reg [119:0] Fsm_currentState_string;
  reg [119:0] Fsm_nextState_string;
  `endif


  assign _zz_Raddr_Init_Cnt_valid = (Kernel_Size - 5'h01);
  assign _zz_Raddr_Update_Cnt_valid = (Stride - 5'h01);
  assign _zz_In_Channel_Process_Cnt_valid = (_zz_In_Channel_Process_Cnt_valid_1 - 13'h0001);
  assign _zz_In_Channel_Process_Cnt_valid_1 = (InFeature_Channel >>> 3);
  assign _zz_Window_Col_Cnt_valid_1 = (Kernel_Size - 5'h01);
  assign _zz_Window_Col_Cnt_valid = {11'd0, _zz_Window_Col_Cnt_valid_1};
  assign _zz_Window_Row_Cnt_valid_1 = (Kernel_Size - 5'h01);
  assign _zz_Window_Row_Cnt_valid = {11'd0, _zz_Window_Row_Cnt_valid_1};
  assign _zz_Out_Channel_Cnt_valid = (OutFeature_Channel_Count_Times - 16'h0001);
  assign _zz_Out_Col_Cnt_valid = (OutCol_Count_Times - 16'h0001);
  assign _zz_when_Data_Generate_V2_l446 = {13'd0, SA_Row_Cnt_count};
  assign _zz_when_Data_Generate_V2_l446_1 = (OutFeature_Col_Lefted - 16'h0001);
  assign _zz_WindowSize_Cnt_valid = {3'd0, WindowSize_Cnt_count};
  assign _zz_WindowSize_Cnt_valid_1 = (Window_Size - 16'h0001);
  assign _zz_Kernel_Base_Addr_1 = ({3'd0,Sliding_Size} <<< 3);
  assign _zz_Kernel_Base_Addr = {16'd0, _zz_Kernel_Base_Addr_1};
  assign _zz_Kernel_Addr_1 = ({3'd0,Sliding_Size} <<< 3);
  assign _zz_Kernel_Addr = {16'd0, _zz_Kernel_Addr_1};
  assign _zz_Kernel_Addr_2 = (Kernel_Base_Addr + _zz_Kernel_Addr_3);
  assign _zz_Kernel_Addr_3 = {19'd0, WindowSize_Cnt_count};
  assign _zz_Kernel_Addr_4 = {19'd0, Sliding_Size};
  assign _zz_Raddr = (Kernel_Addr + _zz_Raddr_1);
  assign _zz_Raddr_1 = {16'd0, Row_Base_Addr};
  WaddrOffset_Fifo RaddrFifo1 (
    .io_push_valid   (RaddrFifo1_io_push_valid        ), //i
    .io_push_ready   (RaddrFifo1_io_push_ready        ), //o
    .io_push_payload (RaddrFifo1_io_push_payload[15:0]), //i
    .io_pop_valid    (RaddrFifo1_io_pop_valid         ), //o
    .io_pop_ready    (RaddrFifo1_io_pop_ready         ), //i
    .io_pop_payload  (RaddrFifo1_io_pop_payload[15:0] ), //o
    .io_flush        (RaddrFifo1_io_flush             ), //i
    .io_occupancy    (RaddrFifo1_io_occupancy[5:0]    ), //o
    .io_availability (RaddrFifo1_io_availability[5:0] ), //o
    .clk             (clk                             ), //i
    .reset           (reset                           )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      IMG2COL_OUTPUT_ENUM_IDLE : Fsm_currentState_string = "IDLE           ";
      IMG2COL_OUTPUT_ENUM_INIT : Fsm_currentState_string = "INIT           ";
      IMG2COL_OUTPUT_ENUM_INIT_ADDR : Fsm_currentState_string = "INIT_ADDR      ";
      IMG2COL_OUTPUT_ENUM_SA_COMPUTE : Fsm_currentState_string = "SA_COMPUTE     ";
      IMG2COL_OUTPUT_ENUM_UPDATE_ADDR : Fsm_currentState_string = "UPDATE_ADDR    ";
      IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY : Fsm_currentState_string = "WAIT_NEXT_READY";
      default : Fsm_currentState_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      IMG2COL_OUTPUT_ENUM_IDLE : Fsm_nextState_string = "IDLE           ";
      IMG2COL_OUTPUT_ENUM_INIT : Fsm_nextState_string = "INIT           ";
      IMG2COL_OUTPUT_ENUM_INIT_ADDR : Fsm_nextState_string = "INIT_ADDR      ";
      IMG2COL_OUTPUT_ENUM_SA_COMPUTE : Fsm_nextState_string = "SA_COMPUTE     ";
      IMG2COL_OUTPUT_ENUM_UPDATE_ADDR : Fsm_nextState_string = "UPDATE_ADDR    ";
      IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY : Fsm_nextState_string = "WAIT_NEXT_READY";
      default : Fsm_nextState_string = "???????????????";
    endcase
  end
  `endif

  assign when_Data_Generate_V2_l303 = (start && (! start_regNext));
  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_IDLE) == IMG2COL_OUTPUT_ENUM_IDLE) : begin
        if(when_Data_Generate_V2_l303) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_INIT;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_IDLE;
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_INIT) == IMG2COL_OUTPUT_ENUM_INIT) : begin
        if(Fsm_Init_End) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_INIT_ADDR;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_INIT;
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_INIT_ADDR) == IMG2COL_OUTPUT_ENUM_INIT_ADDR) : begin
        if(Fsm_Addr_Inited) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_INIT_ADDR;
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY) == IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY) : begin
        if(Fsm_NextReady) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_SA_COMPUTE;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY;
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) == IMG2COL_OUTPUT_ENUM_SA_COMPUTE) : begin
        if(Fsm_LayerEnd) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_IDLE;
        end else begin
          if(Fsm_SA_Computed) begin
            Fsm_nextState = IMG2COL_OUTPUT_ENUM_UPDATE_ADDR;
          end else begin
            if(when_Data_Generate_V2_l335) begin
              Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY;
            end else begin
              Fsm_nextState = IMG2COL_OUTPUT_ENUM_SA_COMPUTE;
            end
          end
        end
      end
      default : begin
        if(Fsm_Addr_Updated) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_UPDATE_ADDR;
        end
      end
    endcase
  end

  assign when_Data_Generate_V2_l335 = (! Fsm_NextReady);
  assign when_WaCounter_l18 = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT) != 6'b000000);
  assign when_WaCounter_l13 = (Init_Count_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l13) begin
      Init_Count_valid = 1'b1;
    end else begin
      Init_Count_valid = 1'b0;
    end
  end

  assign Fsm_Init_End = Init_Count_valid;
  assign NewAddrIn_ready = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT_ADDR) != 6'b000000) || ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 6'b000000));
  always @(*) begin
    RaddrFifo1_io_push_valid = 1'b0;
    if(when_Data_Generate_V2_l481) begin
      RaddrFifo1_io_push_valid = NewAddrIn_valid;
    end else begin
      if(when_Data_Generate_V2_l485) begin
        RaddrFifo1_io_push_valid = NewAddrIn_valid;
      end else begin
        RaddrFifo1_io_push_valid = Window_Col_Cnt_valid;
      end
    end
  end

  always @(*) begin
    RaddrFifo1_io_pop_ready = 1'b0;
    if(when_Data_Generate_V2_l412) begin
      RaddrFifo1_io_pop_ready = 1'b1;
    end
    if(!when_Data_Generate_V2_l481) begin
      if(when_Data_Generate_V2_l485) begin
        RaddrFifo1_io_pop_ready = RaddrFifo1_io_push_fire_2;
      end
    end
    if(Window_Col_Cnt_valid) begin
      RaddrFifo1_io_pop_ready = 1'b1;
    end
  end

  assign RaddrFifo1_io_pop_fire = (RaddrFifo1_io_pop_valid && RaddrFifo1_io_pop_ready);
  assign RaddrFifo1_io_push_fire = (RaddrFifo1_io_push_valid && RaddrFifo1_io_push_ready);
  assign when_WaCounter_l37 = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT_ADDR) != 6'b000000) && RaddrFifo1_io_push_fire);
  assign Raddr_Init_Cnt_valid = ((Raddr_Init_Cnt_count == _zz_Raddr_Init_Cnt_valid) && when_WaCounter_l37);
  assign Fsm_Addr_Inited = Raddr_Init_Cnt_valid;
  assign RaddrFifo1_io_push_fire_1 = (RaddrFifo1_io_push_valid && RaddrFifo1_io_push_ready);
  assign when_WaCounter_l37_1 = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 6'b000000) && RaddrFifo1_io_push_fire_1);
  assign Raddr_Update_Cnt_valid = ((Raddr_Update_Cnt_count == _zz_Raddr_Update_Cnt_valid) && when_WaCounter_l37_1);
  assign Fsm_Addr_Updated = Raddr_Update_Cnt_valid;
  assign Fsm_NextReady = mReady;
  always @(*) begin
    AddrReceived = 1'b0;
    if(when_Data_Generate_V2_l412) begin
      AddrReceived = 1'b1;
    end
  end

  assign when_Data_Generate_V2_l412 = ((((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT_ADDR) != 6'b000000) && ((Fsm_nextState & IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY) != 6'b000000)) || (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 6'b000000) && ((Fsm_nextState & IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY) != 6'b000000)));
  assign when_WaCounter_l37_2 = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) != 6'b000000) && mReady);
  always @(*) begin
    SA_Row_Cnt_valid = ((SA_Row_Cnt_count == 3'b111) && when_WaCounter_l37_2);
    if(when_Data_Generate_V2_l446) begin
      SA_Row_Cnt_valid = 1'b1;
    end
  end

  assign In_Channel_Process_Cnt_valid = ((In_Channel_Process_Cnt_count == _zz_In_Channel_Process_Cnt_valid) && SA_Row_Cnt_valid);
  assign Window_Col_Cnt_valid = ((Window_Col_Cnt_count == _zz_Window_Col_Cnt_valid) && In_Channel_Process_Cnt_valid);
  assign Window_Row_Cnt_valid = ((Window_Row_Cnt_count == _zz_Window_Row_Cnt_valid) && Window_Col_Cnt_valid);
  assign Out_Channel_Cnt_valid = ((Out_Channel_Cnt_count == _zz_Out_Channel_Cnt_valid) && Window_Row_Cnt_valid);
  assign Out_Col_Cnt_valid = ((Out_Col_Cnt_count == _zz_Out_Col_Cnt_valid) && Out_Channel_Cnt_valid);
  assign SA_End = Out_Col_Cnt_valid;
  assign when_Data_Generate_V2_l443 = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT) != 6'b000000);
  assign when_Data_Generate_V2_l446 = (((_zz_when_Data_Generate_V2_l446 == _zz_when_Data_Generate_V2_l446_1) && mReady) && ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) != 6'b000000));
  assign WindowSize_Cnt_valid = ((_zz_WindowSize_Cnt_valid == _zz_WindowSize_Cnt_valid_1) && SA_Row_Cnt_valid);
  assign when_Data_Generate_V2_l471 = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) != 6'b000000) && mReady);
  assign Raddr = _zz_Raddr[15:0];
  assign Fsm_SA_Computed = Out_Col_Cnt_valid;
  assign SA_Idle = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_IDLE) != 6'b000000) || ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 6'b000000));
  assign when_Data_Generate_V2_l481 = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT_ADDR) != 6'b000000);
  always @(*) begin
    if(when_Data_Generate_V2_l481) begin
      RaddrFifo1_io_push_payload = NewAddrIn_payload;
    end else begin
      if(when_Data_Generate_V2_l485) begin
        RaddrFifo1_io_push_payload = NewAddrIn_payload;
      end else begin
        RaddrFifo1_io_push_payload = Row_Base_Addr;
      end
    end
  end

  assign RaddrFifo1_io_push_fire_2 = (RaddrFifo1_io_push_valid && RaddrFifo1_io_push_ready);
  assign when_Data_Generate_V2_l485 = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 6'b000000);
  assign Raddr_Valid = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) != 6'b000000) && mReady);
  assign Fsm_LayerEnd = LayerEnd;
  assign RaddrFifo1_io_flush = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_IDLE) != 6'b000000);
  always @(posedge clk) begin
    start_regNext <= start;
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= IMG2COL_OUTPUT_ENUM_IDLE;
      Init_Count_count <= 3'b000;
      Row_Base_Addr <= 16'h0;
      Raddr_Init_Cnt_count <= 5'h0;
      Raddr_Update_Cnt_count <= 5'h0;
      SA_Row_Cnt_count <= 3'b000;
      In_Channel_Process_Cnt_count <= 13'h0;
      Window_Col_Cnt_count <= 16'h0;
      Window_Row_Cnt_count <= 16'h0;
      Out_Channel_Cnt_count <= 16'h0;
      Out_Col_Cnt_count <= 16'h0;
      OutFeature_Col_Lefted <= 16'h0;
      WindowSize_Cnt_count <= 13'h0;
      Kernel_Addr <= 32'h0;
      Kernel_Base_Addr <= 32'h0;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l18) begin
        Init_Count_count <= (Init_Count_count + 3'b001);
        if(Init_Count_valid) begin
          Init_Count_count <= 3'b000;
        end
      end
      if(RaddrFifo1_io_pop_fire) begin
        Row_Base_Addr <= RaddrFifo1_io_pop_payload;
      end
      if(when_WaCounter_l37) begin
        if(Raddr_Init_Cnt_valid) begin
          Raddr_Init_Cnt_count <= 5'h0;
        end else begin
          Raddr_Init_Cnt_count <= (Raddr_Init_Cnt_count + 5'h01);
        end
      end
      if(when_WaCounter_l37_1) begin
        if(Raddr_Update_Cnt_valid) begin
          Raddr_Update_Cnt_count <= 5'h0;
        end else begin
          Raddr_Update_Cnt_count <= (Raddr_Update_Cnt_count + 5'h01);
        end
      end
      if(when_WaCounter_l37_2) begin
        if(SA_Row_Cnt_valid) begin
          SA_Row_Cnt_count <= 3'b000;
        end else begin
          SA_Row_Cnt_count <= (SA_Row_Cnt_count + 3'b001);
        end
      end
      if(SA_Row_Cnt_valid) begin
        if(In_Channel_Process_Cnt_valid) begin
          In_Channel_Process_Cnt_count <= 13'h0;
        end else begin
          In_Channel_Process_Cnt_count <= (In_Channel_Process_Cnt_count + 13'h0001);
        end
      end
      if(In_Channel_Process_Cnt_valid) begin
        if(Window_Col_Cnt_valid) begin
          Window_Col_Cnt_count <= 16'h0;
        end else begin
          Window_Col_Cnt_count <= (Window_Col_Cnt_count + 16'h0001);
        end
      end
      if(Window_Col_Cnt_valid) begin
        if(Window_Row_Cnt_valid) begin
          Window_Row_Cnt_count <= 16'h0;
        end else begin
          Window_Row_Cnt_count <= (Window_Row_Cnt_count + 16'h0001);
        end
      end
      if(Window_Row_Cnt_valid) begin
        if(Out_Channel_Cnt_valid) begin
          Out_Channel_Cnt_count <= 16'h0;
        end else begin
          Out_Channel_Cnt_count <= (Out_Channel_Cnt_count + 16'h0001);
        end
      end
      if(Out_Channel_Cnt_valid) begin
        if(Out_Col_Cnt_valid) begin
          Out_Col_Cnt_count <= 16'h0;
        end else begin
          Out_Col_Cnt_count <= (Out_Col_Cnt_count + 16'h0001);
        end
      end
      if(Out_Col_Cnt_valid) begin
        OutFeature_Col_Lefted <= OutFeature_Size;
      end else begin
        if(Out_Channel_Cnt_valid) begin
          OutFeature_Col_Lefted <= (OutFeature_Col_Lefted - 16'h0008);
        end else begin
          if(when_Data_Generate_V2_l443) begin
            OutFeature_Col_Lefted <= OutFeature_Size;
          end
        end
      end
      if(when_Data_Generate_V2_l446) begin
        SA_Row_Cnt_count <= 3'b000;
      end
      if(SA_Row_Cnt_valid) begin
        if(WindowSize_Cnt_valid) begin
          WindowSize_Cnt_count <= 13'h0;
        end else begin
          WindowSize_Cnt_count <= (WindowSize_Cnt_count + 13'h0001);
        end
      end
      if(Out_Col_Cnt_valid) begin
        Kernel_Base_Addr <= 32'h0;
      end else begin
        if(Out_Channel_Cnt_valid) begin
          Kernel_Base_Addr <= (Kernel_Base_Addr + _zz_Kernel_Base_Addr);
        end
      end
      if(Out_Col_Cnt_valid) begin
        Kernel_Addr <= 32'h0;
      end else begin
        if(Out_Channel_Cnt_valid) begin
          Kernel_Addr <= (Kernel_Base_Addr + _zz_Kernel_Addr);
        end else begin
          if(Window_Row_Cnt_valid) begin
            Kernel_Addr <= Kernel_Base_Addr;
          end else begin
            if(WindowSize_Cnt_valid) begin
              Kernel_Addr <= Kernel_Base_Addr;
            end else begin
              if(SA_Row_Cnt_valid) begin
                Kernel_Addr <= (_zz_Kernel_Addr_2 + 32'h00000001);
              end else begin
                if(when_Data_Generate_V2_l471) begin
                  Kernel_Addr <= (Kernel_Addr + _zz_Kernel_Addr_4);
                end
              end
            end
          end
        end
      end
    end
  end


endmodule

//WaddrOffset_Fifo replaced by WaddrOffset_Fifo

//WaddrOffset_Fifo replaced by WaddrOffset_Fifo

module WaddrOffset_Fifo (
  input               io_push_valid,
  output              io_push_ready,
  input      [15:0]   io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [15:0]   io_pop_payload,
  input               io_flush,
  output reg [5:0]    io_occupancy,
  output reg [5:0]    io_availability,
  input               clk,
  input               reset
);

  reg        [15:0]   _zz_logic_ram_port0;
  wire       [5:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [5:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [15:0]   _zz_logic_ram_port_1;
  wire       [5:0]    _zz_io_occupancy;
  wire       [5:0]    _zz_io_availability;
  wire       [5:0]    _zz_io_availability_1;
  wire       [5:0]    _zz_io_availability_2;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [5:0]    logic_pushPtr_valueNext;
  reg        [5:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [5:0]    logic_popPtr_valueNext;
  reg        [5:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1021;
  wire       [5:0]    logic_ptrDif;
  reg [15:0] logic_ram [0:32];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {5'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {5'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_occupancy = (6'h21 + logic_ptrDif);
  assign _zz_io_availability = (6'h21 + _zz_io_availability_1);
  assign _zz_io_availability_1 = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_availability_2 = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  assign _zz_logic_ram_port_1 = io_push_payload;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 6'h20);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    if(logic_pushPtr_willOverflow) begin
      logic_pushPtr_valueNext = 6'h0;
    end else begin
      logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    end
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 6'h0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 6'h20);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    if(logic_popPtr_willOverflow) begin
      logic_popPtr_valueNext = 6'h0;
    end else begin
      logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    end
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 6'h0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1021 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  always @(*) begin
    if(logic_ptrMatch) begin
      io_occupancy = (logic_risingOccupancy ? 6'h21 : 6'h0);
    end else begin
      io_occupancy = ((logic_popPtr_value < logic_pushPtr_value) ? logic_ptrDif : _zz_io_occupancy);
    end
  end

  always @(*) begin
    if(logic_ptrMatch) begin
      io_availability = (logic_risingOccupancy ? 6'h0 : 6'h21);
    end else begin
      io_availability = ((logic_popPtr_value < logic_pushPtr_value) ? _zz_io_availability : _zz_io_availability_2);
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_pushPtr_value <= 6'h0;
      logic_popPtr_value <= 6'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1021) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule
