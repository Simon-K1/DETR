// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : SA_2D
// Git hash  : ae0794446f1a331f88fb3854541dace15ffb33b0

`timescale 1ns/1ps

module SA_2D (
  input      [7:0]    io_MatrixA_0,
  input      [7:0]    io_MatrixA_1,
  input      [7:0]    io_MatrixA_2,
  input      [7:0]    io_MatrixA_3,
  input      [7:0]    io_MatrixA_4,
  input      [7:0]    io_MatrixA_5,
  input      [7:0]    io_MatrixA_6,
  input      [7:0]    io_MatrixA_7,
  input      [7:0]    io_MatrixB_0,
  input      [7:0]    io_MatrixB_1,
  input      [7:0]    io_MatrixB_2,
  input      [7:0]    io_MatrixB_3,
  input      [7:0]    io_MatrixB_4,
  input      [7:0]    io_MatrixB_5,
  input      [7:0]    io_MatrixB_6,
  input      [7:0]    io_MatrixB_7,
  input               io_A_Valid_0,
  input               io_A_Valid_1,
  input               io_A_Valid_2,
  input               io_A_Valid_3,
  input               io_A_Valid_4,
  input               io_A_Valid_5,
  input               io_A_Valid_6,
  input               io_A_Valid_7,
  input               io_B_Valid_0,
  input               io_B_Valid_1,
  input               io_B_Valid_2,
  input               io_B_Valid_3,
  input               io_B_Valid_4,
  input               io_B_Valid_5,
  input               io_B_Valid_6,
  input               io_B_Valid_7,
  input      [15:0]   io_signCount,
  output reg [31:0]   MatrixC_0,
  output reg [31:0]   MatrixC_1,
  output reg [31:0]   MatrixC_2,
  output reg [31:0]   MatrixC_3,
  output reg [31:0]   MatrixC_4,
  output reg [31:0]   MatrixC_5,
  output reg [31:0]   MatrixC_6,
  output reg [31:0]   MatrixC_7,
  input               start,
  input               clk,
  input               reset
);

  wire                PE00_valid;
  wire                PE01_valid;
  wire                PE02_valid;
  wire                PE03_valid;
  wire                PE04_valid;
  wire                PE05_valid;
  wire                PE06_valid;
  wire                PE07_valid;
  wire                PE10_valid;
  wire                PE11_valid;
  wire                PE12_valid;
  wire                PE13_valid;
  wire                PE14_valid;
  wire                PE15_valid;
  wire                PE16_valid;
  wire                PE17_valid;
  wire                PE20_valid;
  wire                PE21_valid;
  wire                PE22_valid;
  wire                PE23_valid;
  wire                PE24_valid;
  wire                PE25_valid;
  wire                PE26_valid;
  wire                PE27_valid;
  wire                PE30_valid;
  wire                PE31_valid;
  wire                PE32_valid;
  wire                PE33_valid;
  wire                PE34_valid;
  wire                PE35_valid;
  wire                PE36_valid;
  wire                PE37_valid;
  wire                PE40_valid;
  wire                PE41_valid;
  wire                PE42_valid;
  wire                PE43_valid;
  wire                PE44_valid;
  wire                PE45_valid;
  wire                PE46_valid;
  wire                PE47_valid;
  wire                PE50_valid;
  wire                PE51_valid;
  wire                PE52_valid;
  wire                PE53_valid;
  wire                PE54_valid;
  wire                PE55_valid;
  wire                PE56_valid;
  wire                PE57_valid;
  wire                PE60_valid;
  wire                PE61_valid;
  wire                PE62_valid;
  wire                PE63_valid;
  wire                PE64_valid;
  wire                PE65_valid;
  wire                PE66_valid;
  wire                PE67_valid;
  wire                PE70_valid;
  wire                PE71_valid;
  wire                PE72_valid;
  wire                PE73_valid;
  wire                PE74_valid;
  wire                PE75_valid;
  wire                PE76_valid;
  wire                PE77_valid;
  wire       [7:0]    PE00_acount;
  wire       [7:0]    PE00_bcount;
  wire       [31:0]   PE00_PE_OUT;
  wire                PE00_finish;
  wire       [7:0]    PE01_acount;
  wire       [7:0]    PE01_bcount;
  wire       [31:0]   PE01_PE_OUT;
  wire                PE01_finish;
  wire       [7:0]    PE02_acount;
  wire       [7:0]    PE02_bcount;
  wire       [31:0]   PE02_PE_OUT;
  wire                PE02_finish;
  wire       [7:0]    PE03_acount;
  wire       [7:0]    PE03_bcount;
  wire       [31:0]   PE03_PE_OUT;
  wire                PE03_finish;
  wire       [7:0]    PE04_acount;
  wire       [7:0]    PE04_bcount;
  wire       [31:0]   PE04_PE_OUT;
  wire                PE04_finish;
  wire       [7:0]    PE05_acount;
  wire       [7:0]    PE05_bcount;
  wire       [31:0]   PE05_PE_OUT;
  wire                PE05_finish;
  wire       [7:0]    PE06_acount;
  wire       [7:0]    PE06_bcount;
  wire       [31:0]   PE06_PE_OUT;
  wire                PE06_finish;
  wire       [7:0]    PE07_acount;
  wire       [7:0]    PE07_bcount;
  wire       [31:0]   PE07_PE_OUT;
  wire                PE07_finish;
  wire       [7:0]    PE10_acount;
  wire       [7:0]    PE10_bcount;
  wire       [31:0]   PE10_PE_OUT;
  wire                PE10_finish;
  wire       [7:0]    PE11_acount;
  wire       [7:0]    PE11_bcount;
  wire       [31:0]   PE11_PE_OUT;
  wire                PE11_finish;
  wire       [7:0]    PE12_acount;
  wire       [7:0]    PE12_bcount;
  wire       [31:0]   PE12_PE_OUT;
  wire                PE12_finish;
  wire       [7:0]    PE13_acount;
  wire       [7:0]    PE13_bcount;
  wire       [31:0]   PE13_PE_OUT;
  wire                PE13_finish;
  wire       [7:0]    PE14_acount;
  wire       [7:0]    PE14_bcount;
  wire       [31:0]   PE14_PE_OUT;
  wire                PE14_finish;
  wire       [7:0]    PE15_acount;
  wire       [7:0]    PE15_bcount;
  wire       [31:0]   PE15_PE_OUT;
  wire                PE15_finish;
  wire       [7:0]    PE16_acount;
  wire       [7:0]    PE16_bcount;
  wire       [31:0]   PE16_PE_OUT;
  wire                PE16_finish;
  wire       [7:0]    PE17_acount;
  wire       [7:0]    PE17_bcount;
  wire       [31:0]   PE17_PE_OUT;
  wire                PE17_finish;
  wire       [7:0]    PE20_acount;
  wire       [7:0]    PE20_bcount;
  wire       [31:0]   PE20_PE_OUT;
  wire                PE20_finish;
  wire       [7:0]    PE21_acount;
  wire       [7:0]    PE21_bcount;
  wire       [31:0]   PE21_PE_OUT;
  wire                PE21_finish;
  wire       [7:0]    PE22_acount;
  wire       [7:0]    PE22_bcount;
  wire       [31:0]   PE22_PE_OUT;
  wire                PE22_finish;
  wire       [7:0]    PE23_acount;
  wire       [7:0]    PE23_bcount;
  wire       [31:0]   PE23_PE_OUT;
  wire                PE23_finish;
  wire       [7:0]    PE24_acount;
  wire       [7:0]    PE24_bcount;
  wire       [31:0]   PE24_PE_OUT;
  wire                PE24_finish;
  wire       [7:0]    PE25_acount;
  wire       [7:0]    PE25_bcount;
  wire       [31:0]   PE25_PE_OUT;
  wire                PE25_finish;
  wire       [7:0]    PE26_acount;
  wire       [7:0]    PE26_bcount;
  wire       [31:0]   PE26_PE_OUT;
  wire                PE26_finish;
  wire       [7:0]    PE27_acount;
  wire       [7:0]    PE27_bcount;
  wire       [31:0]   PE27_PE_OUT;
  wire                PE27_finish;
  wire       [7:0]    PE30_acount;
  wire       [7:0]    PE30_bcount;
  wire       [31:0]   PE30_PE_OUT;
  wire                PE30_finish;
  wire       [7:0]    PE31_acount;
  wire       [7:0]    PE31_bcount;
  wire       [31:0]   PE31_PE_OUT;
  wire                PE31_finish;
  wire       [7:0]    PE32_acount;
  wire       [7:0]    PE32_bcount;
  wire       [31:0]   PE32_PE_OUT;
  wire                PE32_finish;
  wire       [7:0]    PE33_acount;
  wire       [7:0]    PE33_bcount;
  wire       [31:0]   PE33_PE_OUT;
  wire                PE33_finish;
  wire       [7:0]    PE34_acount;
  wire       [7:0]    PE34_bcount;
  wire       [31:0]   PE34_PE_OUT;
  wire                PE34_finish;
  wire       [7:0]    PE35_acount;
  wire       [7:0]    PE35_bcount;
  wire       [31:0]   PE35_PE_OUT;
  wire                PE35_finish;
  wire       [7:0]    PE36_acount;
  wire       [7:0]    PE36_bcount;
  wire       [31:0]   PE36_PE_OUT;
  wire                PE36_finish;
  wire       [7:0]    PE37_acount;
  wire       [7:0]    PE37_bcount;
  wire       [31:0]   PE37_PE_OUT;
  wire                PE37_finish;
  wire       [7:0]    PE40_acount;
  wire       [7:0]    PE40_bcount;
  wire       [31:0]   PE40_PE_OUT;
  wire                PE40_finish;
  wire       [7:0]    PE41_acount;
  wire       [7:0]    PE41_bcount;
  wire       [31:0]   PE41_PE_OUT;
  wire                PE41_finish;
  wire       [7:0]    PE42_acount;
  wire       [7:0]    PE42_bcount;
  wire       [31:0]   PE42_PE_OUT;
  wire                PE42_finish;
  wire       [7:0]    PE43_acount;
  wire       [7:0]    PE43_bcount;
  wire       [31:0]   PE43_PE_OUT;
  wire                PE43_finish;
  wire       [7:0]    PE44_acount;
  wire       [7:0]    PE44_bcount;
  wire       [31:0]   PE44_PE_OUT;
  wire                PE44_finish;
  wire       [7:0]    PE45_acount;
  wire       [7:0]    PE45_bcount;
  wire       [31:0]   PE45_PE_OUT;
  wire                PE45_finish;
  wire       [7:0]    PE46_acount;
  wire       [7:0]    PE46_bcount;
  wire       [31:0]   PE46_PE_OUT;
  wire                PE46_finish;
  wire       [7:0]    PE47_acount;
  wire       [7:0]    PE47_bcount;
  wire       [31:0]   PE47_PE_OUT;
  wire                PE47_finish;
  wire       [7:0]    PE50_acount;
  wire       [7:0]    PE50_bcount;
  wire       [31:0]   PE50_PE_OUT;
  wire                PE50_finish;
  wire       [7:0]    PE51_acount;
  wire       [7:0]    PE51_bcount;
  wire       [31:0]   PE51_PE_OUT;
  wire                PE51_finish;
  wire       [7:0]    PE52_acount;
  wire       [7:0]    PE52_bcount;
  wire       [31:0]   PE52_PE_OUT;
  wire                PE52_finish;
  wire       [7:0]    PE53_acount;
  wire       [7:0]    PE53_bcount;
  wire       [31:0]   PE53_PE_OUT;
  wire                PE53_finish;
  wire       [7:0]    PE54_acount;
  wire       [7:0]    PE54_bcount;
  wire       [31:0]   PE54_PE_OUT;
  wire                PE54_finish;
  wire       [7:0]    PE55_acount;
  wire       [7:0]    PE55_bcount;
  wire       [31:0]   PE55_PE_OUT;
  wire                PE55_finish;
  wire       [7:0]    PE56_acount;
  wire       [7:0]    PE56_bcount;
  wire       [31:0]   PE56_PE_OUT;
  wire                PE56_finish;
  wire       [7:0]    PE57_acount;
  wire       [7:0]    PE57_bcount;
  wire       [31:0]   PE57_PE_OUT;
  wire                PE57_finish;
  wire       [7:0]    PE60_acount;
  wire       [7:0]    PE60_bcount;
  wire       [31:0]   PE60_PE_OUT;
  wire                PE60_finish;
  wire       [7:0]    PE61_acount;
  wire       [7:0]    PE61_bcount;
  wire       [31:0]   PE61_PE_OUT;
  wire                PE61_finish;
  wire       [7:0]    PE62_acount;
  wire       [7:0]    PE62_bcount;
  wire       [31:0]   PE62_PE_OUT;
  wire                PE62_finish;
  wire       [7:0]    PE63_acount;
  wire       [7:0]    PE63_bcount;
  wire       [31:0]   PE63_PE_OUT;
  wire                PE63_finish;
  wire       [7:0]    PE64_acount;
  wire       [7:0]    PE64_bcount;
  wire       [31:0]   PE64_PE_OUT;
  wire                PE64_finish;
  wire       [7:0]    PE65_acount;
  wire       [7:0]    PE65_bcount;
  wire       [31:0]   PE65_PE_OUT;
  wire                PE65_finish;
  wire       [7:0]    PE66_acount;
  wire       [7:0]    PE66_bcount;
  wire       [31:0]   PE66_PE_OUT;
  wire                PE66_finish;
  wire       [7:0]    PE67_acount;
  wire       [7:0]    PE67_bcount;
  wire       [31:0]   PE67_PE_OUT;
  wire                PE67_finish;
  wire       [7:0]    PE70_acount;
  wire       [7:0]    PE70_bcount;
  wire       [31:0]   PE70_PE_OUT;
  wire                PE70_finish;
  wire       [7:0]    PE71_acount;
  wire       [7:0]    PE71_bcount;
  wire       [31:0]   PE71_PE_OUT;
  wire                PE71_finish;
  wire       [7:0]    PE72_acount;
  wire       [7:0]    PE72_bcount;
  wire       [31:0]   PE72_PE_OUT;
  wire                PE72_finish;
  wire       [7:0]    PE73_acount;
  wire       [7:0]    PE73_bcount;
  wire       [31:0]   PE73_PE_OUT;
  wire                PE73_finish;
  wire       [7:0]    PE74_acount;
  wire       [7:0]    PE74_bcount;
  wire       [31:0]   PE74_PE_OUT;
  wire                PE74_finish;
  wire       [7:0]    PE75_acount;
  wire       [7:0]    PE75_bcount;
  wire       [31:0]   PE75_PE_OUT;
  wire                PE75_finish;
  wire       [7:0]    PE76_acount;
  wire       [7:0]    PE76_bcount;
  wire       [31:0]   PE76_PE_OUT;
  wire                PE76_finish;
  wire       [7:0]    PE77_acount;
  wire       [7:0]    PE77_bcount;
  wire       [31:0]   PE77_PE_OUT;
  wire                PE77_finish;
  reg        [15:0]   io_signCount_regNextWhen;
  reg                 io_A_Valid_0_delay_1;
  reg                 io_A_Valid_0_delay_1_1;
  reg                 io_A_Valid_0_delay_2;
  reg                 io_A_Valid_0_delay_1_2;
  reg                 io_A_Valid_0_delay_2_1;
  reg                 io_A_Valid_0_delay_3;
  reg                 io_A_Valid_0_delay_1_3;
  reg                 io_A_Valid_0_delay_2_2;
  reg                 io_A_Valid_0_delay_3_1;
  reg                 io_A_Valid_0_delay_4;
  reg                 io_A_Valid_0_delay_1_4;
  reg                 io_A_Valid_0_delay_2_3;
  reg                 io_A_Valid_0_delay_3_2;
  reg                 io_A_Valid_0_delay_4_1;
  reg                 io_A_Valid_0_delay_5;
  reg                 io_A_Valid_0_delay_1_5;
  reg                 io_A_Valid_0_delay_2_4;
  reg                 io_A_Valid_0_delay_3_3;
  reg                 io_A_Valid_0_delay_4_2;
  reg                 io_A_Valid_0_delay_5_1;
  reg                 io_A_Valid_0_delay_6;
  reg                 io_A_Valid_0_delay_1_6;
  reg                 io_A_Valid_0_delay_2_5;
  reg                 io_A_Valid_0_delay_3_4;
  reg                 io_A_Valid_0_delay_4_3;
  reg                 io_A_Valid_0_delay_5_2;
  reg                 io_A_Valid_0_delay_6_1;
  reg                 io_A_Valid_0_delay_7;
  reg        [15:0]   io_signCount_regNextWhen_1;
  reg                 io_B_Valid_0_delay_1;
  reg                 io_A_Valid_1_delay_1;
  reg                 io_B_Valid_1_delay_1;
  reg                 io_A_Valid_1_delay_1_1;
  reg                 io_A_Valid_1_delay_2;
  reg                 io_B_Valid_2_delay_1;
  reg                 io_A_Valid_1_delay_1_2;
  reg                 io_A_Valid_1_delay_2_1;
  reg                 io_A_Valid_1_delay_3;
  reg                 io_B_Valid_3_delay_1;
  reg                 io_A_Valid_1_delay_1_3;
  reg                 io_A_Valid_1_delay_2_2;
  reg                 io_A_Valid_1_delay_3_1;
  reg                 io_A_Valid_1_delay_4;
  reg                 io_B_Valid_4_delay_1;
  reg                 io_A_Valid_1_delay_1_4;
  reg                 io_A_Valid_1_delay_2_3;
  reg                 io_A_Valid_1_delay_3_2;
  reg                 io_A_Valid_1_delay_4_1;
  reg                 io_A_Valid_1_delay_5;
  reg                 io_B_Valid_5_delay_1;
  reg                 io_A_Valid_1_delay_1_5;
  reg                 io_A_Valid_1_delay_2_4;
  reg                 io_A_Valid_1_delay_3_3;
  reg                 io_A_Valid_1_delay_4_2;
  reg                 io_A_Valid_1_delay_5_1;
  reg                 io_A_Valid_1_delay_6;
  reg                 io_B_Valid_6_delay_1;
  reg                 io_A_Valid_1_delay_1_6;
  reg                 io_A_Valid_1_delay_2_5;
  reg                 io_A_Valid_1_delay_3_4;
  reg                 io_A_Valid_1_delay_4_3;
  reg                 io_A_Valid_1_delay_5_2;
  reg                 io_A_Valid_1_delay_6_1;
  reg                 io_A_Valid_1_delay_7;
  reg                 io_B_Valid_7_delay_1;
  reg        [15:0]   io_signCount_regNextWhen_2;
  reg                 io_B_Valid_0_delay_1_1;
  reg                 io_B_Valid_0_delay_2;
  reg                 io_A_Valid_2_delay_1;
  reg                 io_B_Valid_1_delay_1_1;
  reg                 io_B_Valid_1_delay_2;
  reg                 io_A_Valid_2_delay_1_1;
  reg                 io_A_Valid_2_delay_2;
  reg                 io_B_Valid_2_delay_1_1;
  reg                 io_B_Valid_2_delay_2;
  reg                 io_A_Valid_2_delay_1_2;
  reg                 io_A_Valid_2_delay_2_1;
  reg                 io_A_Valid_2_delay_3;
  reg                 io_B_Valid_3_delay_1_1;
  reg                 io_B_Valid_3_delay_2;
  reg                 io_A_Valid_2_delay_1_3;
  reg                 io_A_Valid_2_delay_2_2;
  reg                 io_A_Valid_2_delay_3_1;
  reg                 io_A_Valid_2_delay_4;
  reg                 io_B_Valid_4_delay_1_1;
  reg                 io_B_Valid_4_delay_2;
  reg                 io_A_Valid_2_delay_1_4;
  reg                 io_A_Valid_2_delay_2_3;
  reg                 io_A_Valid_2_delay_3_2;
  reg                 io_A_Valid_2_delay_4_1;
  reg                 io_A_Valid_2_delay_5;
  reg                 io_B_Valid_5_delay_1_1;
  reg                 io_B_Valid_5_delay_2;
  reg                 io_A_Valid_2_delay_1_5;
  reg                 io_A_Valid_2_delay_2_4;
  reg                 io_A_Valid_2_delay_3_3;
  reg                 io_A_Valid_2_delay_4_2;
  reg                 io_A_Valid_2_delay_5_1;
  reg                 io_A_Valid_2_delay_6;
  reg                 io_B_Valid_6_delay_1_1;
  reg                 io_B_Valid_6_delay_2;
  reg                 io_A_Valid_2_delay_1_6;
  reg                 io_A_Valid_2_delay_2_5;
  reg                 io_A_Valid_2_delay_3_4;
  reg                 io_A_Valid_2_delay_4_3;
  reg                 io_A_Valid_2_delay_5_2;
  reg                 io_A_Valid_2_delay_6_1;
  reg                 io_A_Valid_2_delay_7;
  reg                 io_B_Valid_7_delay_1_1;
  reg                 io_B_Valid_7_delay_2;
  reg        [15:0]   io_signCount_regNextWhen_3;
  reg                 io_B_Valid_0_delay_1_2;
  reg                 io_B_Valid_0_delay_2_1;
  reg                 io_B_Valid_0_delay_3;
  reg                 io_A_Valid_3_delay_1;
  reg                 io_B_Valid_1_delay_1_2;
  reg                 io_B_Valid_1_delay_2_1;
  reg                 io_B_Valid_1_delay_3;
  reg                 io_A_Valid_3_delay_1_1;
  reg                 io_A_Valid_3_delay_2;
  reg                 io_B_Valid_2_delay_1_2;
  reg                 io_B_Valid_2_delay_2_1;
  reg                 io_B_Valid_2_delay_3;
  reg                 io_A_Valid_3_delay_1_2;
  reg                 io_A_Valid_3_delay_2_1;
  reg                 io_A_Valid_3_delay_3;
  reg                 io_B_Valid_3_delay_1_2;
  reg                 io_B_Valid_3_delay_2_1;
  reg                 io_B_Valid_3_delay_3;
  reg                 io_A_Valid_3_delay_1_3;
  reg                 io_A_Valid_3_delay_2_2;
  reg                 io_A_Valid_3_delay_3_1;
  reg                 io_A_Valid_3_delay_4;
  reg                 io_B_Valid_4_delay_1_2;
  reg                 io_B_Valid_4_delay_2_1;
  reg                 io_B_Valid_4_delay_3;
  reg                 io_A_Valid_3_delay_1_4;
  reg                 io_A_Valid_3_delay_2_3;
  reg                 io_A_Valid_3_delay_3_2;
  reg                 io_A_Valid_3_delay_4_1;
  reg                 io_A_Valid_3_delay_5;
  reg                 io_B_Valid_5_delay_1_2;
  reg                 io_B_Valid_5_delay_2_1;
  reg                 io_B_Valid_5_delay_3;
  reg                 io_A_Valid_3_delay_1_5;
  reg                 io_A_Valid_3_delay_2_4;
  reg                 io_A_Valid_3_delay_3_3;
  reg                 io_A_Valid_3_delay_4_2;
  reg                 io_A_Valid_3_delay_5_1;
  reg                 io_A_Valid_3_delay_6;
  reg                 io_B_Valid_6_delay_1_2;
  reg                 io_B_Valid_6_delay_2_1;
  reg                 io_B_Valid_6_delay_3;
  reg                 io_A_Valid_3_delay_1_6;
  reg                 io_A_Valid_3_delay_2_5;
  reg                 io_A_Valid_3_delay_3_4;
  reg                 io_A_Valid_3_delay_4_3;
  reg                 io_A_Valid_3_delay_5_2;
  reg                 io_A_Valid_3_delay_6_1;
  reg                 io_A_Valid_3_delay_7;
  reg                 io_B_Valid_7_delay_1_2;
  reg                 io_B_Valid_7_delay_2_1;
  reg                 io_B_Valid_7_delay_3;
  reg        [15:0]   io_signCount_regNextWhen_4;
  reg                 io_B_Valid_0_delay_1_3;
  reg                 io_B_Valid_0_delay_2_2;
  reg                 io_B_Valid_0_delay_3_1;
  reg                 io_B_Valid_0_delay_4;
  reg                 io_A_Valid_4_delay_1;
  reg                 io_B_Valid_1_delay_1_3;
  reg                 io_B_Valid_1_delay_2_2;
  reg                 io_B_Valid_1_delay_3_1;
  reg                 io_B_Valid_1_delay_4;
  reg                 io_A_Valid_4_delay_1_1;
  reg                 io_A_Valid_4_delay_2;
  reg                 io_B_Valid_2_delay_1_3;
  reg                 io_B_Valid_2_delay_2_2;
  reg                 io_B_Valid_2_delay_3_1;
  reg                 io_B_Valid_2_delay_4;
  reg                 io_A_Valid_4_delay_1_2;
  reg                 io_A_Valid_4_delay_2_1;
  reg                 io_A_Valid_4_delay_3;
  reg                 io_B_Valid_3_delay_1_3;
  reg                 io_B_Valid_3_delay_2_2;
  reg                 io_B_Valid_3_delay_3_1;
  reg                 io_B_Valid_3_delay_4;
  reg                 io_A_Valid_4_delay_1_3;
  reg                 io_A_Valid_4_delay_2_2;
  reg                 io_A_Valid_4_delay_3_1;
  reg                 io_A_Valid_4_delay_4;
  reg                 io_B_Valid_4_delay_1_3;
  reg                 io_B_Valid_4_delay_2_2;
  reg                 io_B_Valid_4_delay_3_1;
  reg                 io_B_Valid_4_delay_4;
  reg                 io_A_Valid_4_delay_1_4;
  reg                 io_A_Valid_4_delay_2_3;
  reg                 io_A_Valid_4_delay_3_2;
  reg                 io_A_Valid_4_delay_4_1;
  reg                 io_A_Valid_4_delay_5;
  reg                 io_B_Valid_5_delay_1_3;
  reg                 io_B_Valid_5_delay_2_2;
  reg                 io_B_Valid_5_delay_3_1;
  reg                 io_B_Valid_5_delay_4;
  reg                 io_A_Valid_4_delay_1_5;
  reg                 io_A_Valid_4_delay_2_4;
  reg                 io_A_Valid_4_delay_3_3;
  reg                 io_A_Valid_4_delay_4_2;
  reg                 io_A_Valid_4_delay_5_1;
  reg                 io_A_Valid_4_delay_6;
  reg                 io_B_Valid_6_delay_1_3;
  reg                 io_B_Valid_6_delay_2_2;
  reg                 io_B_Valid_6_delay_3_1;
  reg                 io_B_Valid_6_delay_4;
  reg                 io_A_Valid_4_delay_1_6;
  reg                 io_A_Valid_4_delay_2_5;
  reg                 io_A_Valid_4_delay_3_4;
  reg                 io_A_Valid_4_delay_4_3;
  reg                 io_A_Valid_4_delay_5_2;
  reg                 io_A_Valid_4_delay_6_1;
  reg                 io_A_Valid_4_delay_7;
  reg                 io_B_Valid_7_delay_1_3;
  reg                 io_B_Valid_7_delay_2_2;
  reg                 io_B_Valid_7_delay_3_1;
  reg                 io_B_Valid_7_delay_4;
  reg        [15:0]   io_signCount_regNextWhen_5;
  reg                 io_B_Valid_0_delay_1_4;
  reg                 io_B_Valid_0_delay_2_3;
  reg                 io_B_Valid_0_delay_3_2;
  reg                 io_B_Valid_0_delay_4_1;
  reg                 io_B_Valid_0_delay_5;
  reg                 io_A_Valid_5_delay_1;
  reg                 io_B_Valid_1_delay_1_4;
  reg                 io_B_Valid_1_delay_2_3;
  reg                 io_B_Valid_1_delay_3_2;
  reg                 io_B_Valid_1_delay_4_1;
  reg                 io_B_Valid_1_delay_5;
  reg                 io_A_Valid_5_delay_1_1;
  reg                 io_A_Valid_5_delay_2;
  reg                 io_B_Valid_2_delay_1_4;
  reg                 io_B_Valid_2_delay_2_3;
  reg                 io_B_Valid_2_delay_3_2;
  reg                 io_B_Valid_2_delay_4_1;
  reg                 io_B_Valid_2_delay_5;
  reg                 io_A_Valid_5_delay_1_2;
  reg                 io_A_Valid_5_delay_2_1;
  reg                 io_A_Valid_5_delay_3;
  reg                 io_B_Valid_3_delay_1_4;
  reg                 io_B_Valid_3_delay_2_3;
  reg                 io_B_Valid_3_delay_3_2;
  reg                 io_B_Valid_3_delay_4_1;
  reg                 io_B_Valid_3_delay_5;
  reg                 io_A_Valid_5_delay_1_3;
  reg                 io_A_Valid_5_delay_2_2;
  reg                 io_A_Valid_5_delay_3_1;
  reg                 io_A_Valid_5_delay_4;
  reg                 io_B_Valid_4_delay_1_4;
  reg                 io_B_Valid_4_delay_2_3;
  reg                 io_B_Valid_4_delay_3_2;
  reg                 io_B_Valid_4_delay_4_1;
  reg                 io_B_Valid_4_delay_5;
  reg                 io_A_Valid_5_delay_1_4;
  reg                 io_A_Valid_5_delay_2_3;
  reg                 io_A_Valid_5_delay_3_2;
  reg                 io_A_Valid_5_delay_4_1;
  reg                 io_A_Valid_5_delay_5;
  reg                 io_B_Valid_5_delay_1_4;
  reg                 io_B_Valid_5_delay_2_3;
  reg                 io_B_Valid_5_delay_3_2;
  reg                 io_B_Valid_5_delay_4_1;
  reg                 io_B_Valid_5_delay_5;
  reg                 io_A_Valid_5_delay_1_5;
  reg                 io_A_Valid_5_delay_2_4;
  reg                 io_A_Valid_5_delay_3_3;
  reg                 io_A_Valid_5_delay_4_2;
  reg                 io_A_Valid_5_delay_5_1;
  reg                 io_A_Valid_5_delay_6;
  reg                 io_B_Valid_6_delay_1_4;
  reg                 io_B_Valid_6_delay_2_3;
  reg                 io_B_Valid_6_delay_3_2;
  reg                 io_B_Valid_6_delay_4_1;
  reg                 io_B_Valid_6_delay_5;
  reg                 io_A_Valid_5_delay_1_6;
  reg                 io_A_Valid_5_delay_2_5;
  reg                 io_A_Valid_5_delay_3_4;
  reg                 io_A_Valid_5_delay_4_3;
  reg                 io_A_Valid_5_delay_5_2;
  reg                 io_A_Valid_5_delay_6_1;
  reg                 io_A_Valid_5_delay_7;
  reg                 io_B_Valid_7_delay_1_4;
  reg                 io_B_Valid_7_delay_2_3;
  reg                 io_B_Valid_7_delay_3_2;
  reg                 io_B_Valid_7_delay_4_1;
  reg                 io_B_Valid_7_delay_5;
  reg        [15:0]   io_signCount_regNextWhen_6;
  reg                 io_B_Valid_0_delay_1_5;
  reg                 io_B_Valid_0_delay_2_4;
  reg                 io_B_Valid_0_delay_3_3;
  reg                 io_B_Valid_0_delay_4_2;
  reg                 io_B_Valid_0_delay_5_1;
  reg                 io_B_Valid_0_delay_6;
  reg                 io_A_Valid_6_delay_1;
  reg                 io_B_Valid_1_delay_1_5;
  reg                 io_B_Valid_1_delay_2_4;
  reg                 io_B_Valid_1_delay_3_3;
  reg                 io_B_Valid_1_delay_4_2;
  reg                 io_B_Valid_1_delay_5_1;
  reg                 io_B_Valid_1_delay_6;
  reg                 io_A_Valid_6_delay_1_1;
  reg                 io_A_Valid_6_delay_2;
  reg                 io_B_Valid_2_delay_1_5;
  reg                 io_B_Valid_2_delay_2_4;
  reg                 io_B_Valid_2_delay_3_3;
  reg                 io_B_Valid_2_delay_4_2;
  reg                 io_B_Valid_2_delay_5_1;
  reg                 io_B_Valid_2_delay_6;
  reg                 io_A_Valid_6_delay_1_2;
  reg                 io_A_Valid_6_delay_2_1;
  reg                 io_A_Valid_6_delay_3;
  reg                 io_B_Valid_3_delay_1_5;
  reg                 io_B_Valid_3_delay_2_4;
  reg                 io_B_Valid_3_delay_3_3;
  reg                 io_B_Valid_3_delay_4_2;
  reg                 io_B_Valid_3_delay_5_1;
  reg                 io_B_Valid_3_delay_6;
  reg                 io_A_Valid_6_delay_1_3;
  reg                 io_A_Valid_6_delay_2_2;
  reg                 io_A_Valid_6_delay_3_1;
  reg                 io_A_Valid_6_delay_4;
  reg                 io_B_Valid_4_delay_1_5;
  reg                 io_B_Valid_4_delay_2_4;
  reg                 io_B_Valid_4_delay_3_3;
  reg                 io_B_Valid_4_delay_4_2;
  reg                 io_B_Valid_4_delay_5_1;
  reg                 io_B_Valid_4_delay_6;
  reg                 io_A_Valid_6_delay_1_4;
  reg                 io_A_Valid_6_delay_2_3;
  reg                 io_A_Valid_6_delay_3_2;
  reg                 io_A_Valid_6_delay_4_1;
  reg                 io_A_Valid_6_delay_5;
  reg                 io_B_Valid_5_delay_1_5;
  reg                 io_B_Valid_5_delay_2_4;
  reg                 io_B_Valid_5_delay_3_3;
  reg                 io_B_Valid_5_delay_4_2;
  reg                 io_B_Valid_5_delay_5_1;
  reg                 io_B_Valid_5_delay_6;
  reg                 io_A_Valid_6_delay_1_5;
  reg                 io_A_Valid_6_delay_2_4;
  reg                 io_A_Valid_6_delay_3_3;
  reg                 io_A_Valid_6_delay_4_2;
  reg                 io_A_Valid_6_delay_5_1;
  reg                 io_A_Valid_6_delay_6;
  reg                 io_B_Valid_6_delay_1_5;
  reg                 io_B_Valid_6_delay_2_4;
  reg                 io_B_Valid_6_delay_3_3;
  reg                 io_B_Valid_6_delay_4_2;
  reg                 io_B_Valid_6_delay_5_1;
  reg                 io_B_Valid_6_delay_6;
  reg                 io_A_Valid_6_delay_1_6;
  reg                 io_A_Valid_6_delay_2_5;
  reg                 io_A_Valid_6_delay_3_4;
  reg                 io_A_Valid_6_delay_4_3;
  reg                 io_A_Valid_6_delay_5_2;
  reg                 io_A_Valid_6_delay_6_1;
  reg                 io_A_Valid_6_delay_7;
  reg                 io_B_Valid_7_delay_1_5;
  reg                 io_B_Valid_7_delay_2_4;
  reg                 io_B_Valid_7_delay_3_3;
  reg                 io_B_Valid_7_delay_4_2;
  reg                 io_B_Valid_7_delay_5_1;
  reg                 io_B_Valid_7_delay_6;
  reg        [15:0]   io_signCount_regNextWhen_7;
  reg                 io_B_Valid_0_delay_1_6;
  reg                 io_B_Valid_0_delay_2_5;
  reg                 io_B_Valid_0_delay_3_4;
  reg                 io_B_Valid_0_delay_4_3;
  reg                 io_B_Valid_0_delay_5_2;
  reg                 io_B_Valid_0_delay_6_1;
  reg                 io_B_Valid_0_delay_7;
  reg                 io_A_Valid_7_delay_1;
  reg                 io_B_Valid_1_delay_1_6;
  reg                 io_B_Valid_1_delay_2_5;
  reg                 io_B_Valid_1_delay_3_4;
  reg                 io_B_Valid_1_delay_4_3;
  reg                 io_B_Valid_1_delay_5_2;
  reg                 io_B_Valid_1_delay_6_1;
  reg                 io_B_Valid_1_delay_7;
  reg                 io_A_Valid_7_delay_1_1;
  reg                 io_A_Valid_7_delay_2;
  reg                 io_B_Valid_2_delay_1_6;
  reg                 io_B_Valid_2_delay_2_5;
  reg                 io_B_Valid_2_delay_3_4;
  reg                 io_B_Valid_2_delay_4_3;
  reg                 io_B_Valid_2_delay_5_2;
  reg                 io_B_Valid_2_delay_6_1;
  reg                 io_B_Valid_2_delay_7;
  reg                 io_A_Valid_7_delay_1_2;
  reg                 io_A_Valid_7_delay_2_1;
  reg                 io_A_Valid_7_delay_3;
  reg                 io_B_Valid_3_delay_1_6;
  reg                 io_B_Valid_3_delay_2_5;
  reg                 io_B_Valid_3_delay_3_4;
  reg                 io_B_Valid_3_delay_4_3;
  reg                 io_B_Valid_3_delay_5_2;
  reg                 io_B_Valid_3_delay_6_1;
  reg                 io_B_Valid_3_delay_7;
  reg                 io_A_Valid_7_delay_1_3;
  reg                 io_A_Valid_7_delay_2_2;
  reg                 io_A_Valid_7_delay_3_1;
  reg                 io_A_Valid_7_delay_4;
  reg                 io_B_Valid_4_delay_1_6;
  reg                 io_B_Valid_4_delay_2_5;
  reg                 io_B_Valid_4_delay_3_4;
  reg                 io_B_Valid_4_delay_4_3;
  reg                 io_B_Valid_4_delay_5_2;
  reg                 io_B_Valid_4_delay_6_1;
  reg                 io_B_Valid_4_delay_7;
  reg                 io_A_Valid_7_delay_1_4;
  reg                 io_A_Valid_7_delay_2_3;
  reg                 io_A_Valid_7_delay_3_2;
  reg                 io_A_Valid_7_delay_4_1;
  reg                 io_A_Valid_7_delay_5;
  reg                 io_B_Valid_5_delay_1_6;
  reg                 io_B_Valid_5_delay_2_5;
  reg                 io_B_Valid_5_delay_3_4;
  reg                 io_B_Valid_5_delay_4_3;
  reg                 io_B_Valid_5_delay_5_2;
  reg                 io_B_Valid_5_delay_6_1;
  reg                 io_B_Valid_5_delay_7;
  reg                 io_A_Valid_7_delay_1_5;
  reg                 io_A_Valid_7_delay_2_4;
  reg                 io_A_Valid_7_delay_3_3;
  reg                 io_A_Valid_7_delay_4_2;
  reg                 io_A_Valid_7_delay_5_1;
  reg                 io_A_Valid_7_delay_6;
  reg                 io_B_Valid_6_delay_1_6;
  reg                 io_B_Valid_6_delay_2_5;
  reg                 io_B_Valid_6_delay_3_4;
  reg                 io_B_Valid_6_delay_4_3;
  reg                 io_B_Valid_6_delay_5_2;
  reg                 io_B_Valid_6_delay_6_1;
  reg                 io_B_Valid_6_delay_7;
  reg                 io_A_Valid_7_delay_1_6;
  reg                 io_A_Valid_7_delay_2_5;
  reg                 io_A_Valid_7_delay_3_4;
  reg                 io_A_Valid_7_delay_4_3;
  reg                 io_A_Valid_7_delay_5_2;
  reg                 io_A_Valid_7_delay_6_1;
  reg                 io_A_Valid_7_delay_7;
  reg                 io_B_Valid_7_delay_1_6;
  reg                 io_B_Valid_7_delay_2_5;
  reg                 io_B_Valid_7_delay_3_4;
  reg                 io_B_Valid_7_delay_4_3;
  reg                 io_B_Valid_7_delay_5_2;
  reg                 io_B_Valid_7_delay_6_1;
  reg                 io_B_Valid_7_delay_7;

  PE PE00 (
    .activate  (io_MatrixA_0[7:0]             ), //i
    .weight    (io_MatrixB_0[7:0]             ), //i
    .valid     (PE00_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE00_acount[7:0]              ), //o
    .bcount    (PE00_bcount[7:0]              ), //o
    .PE_OUT    (PE00_PE_OUT[31:0]             ), //o
    .finish    (PE00_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE01 (
    .activate  (PE00_acount[7:0]              ), //i
    .weight    (io_MatrixB_1[7:0]             ), //i
    .valid     (PE01_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE01_acount[7:0]              ), //o
    .bcount    (PE01_bcount[7:0]              ), //o
    .PE_OUT    (PE01_PE_OUT[31:0]             ), //o
    .finish    (PE01_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE02 (
    .activate  (PE01_acount[7:0]              ), //i
    .weight    (io_MatrixB_2[7:0]             ), //i
    .valid     (PE02_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE02_acount[7:0]              ), //o
    .bcount    (PE02_bcount[7:0]              ), //o
    .PE_OUT    (PE02_PE_OUT[31:0]             ), //o
    .finish    (PE02_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE03 (
    .activate  (PE02_acount[7:0]              ), //i
    .weight    (io_MatrixB_3[7:0]             ), //i
    .valid     (PE03_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE03_acount[7:0]              ), //o
    .bcount    (PE03_bcount[7:0]              ), //o
    .PE_OUT    (PE03_PE_OUT[31:0]             ), //o
    .finish    (PE03_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE04 (
    .activate  (PE03_acount[7:0]              ), //i
    .weight    (io_MatrixB_4[7:0]             ), //i
    .valid     (PE04_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE04_acount[7:0]              ), //o
    .bcount    (PE04_bcount[7:0]              ), //o
    .PE_OUT    (PE04_PE_OUT[31:0]             ), //o
    .finish    (PE04_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE05 (
    .activate  (PE04_acount[7:0]              ), //i
    .weight    (io_MatrixB_5[7:0]             ), //i
    .valid     (PE05_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE05_acount[7:0]              ), //o
    .bcount    (PE05_bcount[7:0]              ), //o
    .PE_OUT    (PE05_PE_OUT[31:0]             ), //o
    .finish    (PE05_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE06 (
    .activate  (PE05_acount[7:0]              ), //i
    .weight    (io_MatrixB_6[7:0]             ), //i
    .valid     (PE06_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE06_acount[7:0]              ), //o
    .bcount    (PE06_bcount[7:0]              ), //o
    .PE_OUT    (PE06_PE_OUT[31:0]             ), //o
    .finish    (PE06_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE07 (
    .activate  (PE06_acount[7:0]              ), //i
    .weight    (io_MatrixB_7[7:0]             ), //i
    .valid     (PE07_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE07_acount[7:0]              ), //o
    .bcount    (PE07_bcount[7:0]              ), //o
    .PE_OUT    (PE07_PE_OUT[31:0]             ), //o
    .finish    (PE07_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE10 (
    .activate  (io_MatrixA_1[7:0]               ), //i
    .weight    (PE00_bcount[7:0]                ), //i
    .valid     (PE10_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE10_acount[7:0]                ), //o
    .bcount    (PE10_bcount[7:0]                ), //o
    .PE_OUT    (PE10_PE_OUT[31:0]               ), //o
    .finish    (PE10_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE11 (
    .activate  (PE10_acount[7:0]                ), //i
    .weight    (PE01_bcount[7:0]                ), //i
    .valid     (PE11_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE11_acount[7:0]                ), //o
    .bcount    (PE11_bcount[7:0]                ), //o
    .PE_OUT    (PE11_PE_OUT[31:0]               ), //o
    .finish    (PE11_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE12 (
    .activate  (PE11_acount[7:0]                ), //i
    .weight    (PE02_bcount[7:0]                ), //i
    .valid     (PE12_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE12_acount[7:0]                ), //o
    .bcount    (PE12_bcount[7:0]                ), //o
    .PE_OUT    (PE12_PE_OUT[31:0]               ), //o
    .finish    (PE12_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE13 (
    .activate  (PE12_acount[7:0]                ), //i
    .weight    (PE03_bcount[7:0]                ), //i
    .valid     (PE13_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE13_acount[7:0]                ), //o
    .bcount    (PE13_bcount[7:0]                ), //o
    .PE_OUT    (PE13_PE_OUT[31:0]               ), //o
    .finish    (PE13_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE14 (
    .activate  (PE13_acount[7:0]                ), //i
    .weight    (PE04_bcount[7:0]                ), //i
    .valid     (PE14_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE14_acount[7:0]                ), //o
    .bcount    (PE14_bcount[7:0]                ), //o
    .PE_OUT    (PE14_PE_OUT[31:0]               ), //o
    .finish    (PE14_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE15 (
    .activate  (PE14_acount[7:0]                ), //i
    .weight    (PE05_bcount[7:0]                ), //i
    .valid     (PE15_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE15_acount[7:0]                ), //o
    .bcount    (PE15_bcount[7:0]                ), //o
    .PE_OUT    (PE15_PE_OUT[31:0]               ), //o
    .finish    (PE15_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE16 (
    .activate  (PE15_acount[7:0]                ), //i
    .weight    (PE06_bcount[7:0]                ), //i
    .valid     (PE16_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE16_acount[7:0]                ), //o
    .bcount    (PE16_bcount[7:0]                ), //o
    .PE_OUT    (PE16_PE_OUT[31:0]               ), //o
    .finish    (PE16_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE17 (
    .activate  (PE16_acount[7:0]                ), //i
    .weight    (PE07_bcount[7:0]                ), //i
    .valid     (PE17_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE17_acount[7:0]                ), //o
    .bcount    (PE17_bcount[7:0]                ), //o
    .PE_OUT    (PE17_PE_OUT[31:0]               ), //o
    .finish    (PE17_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE20 (
    .activate  (io_MatrixA_2[7:0]               ), //i
    .weight    (PE10_bcount[7:0]                ), //i
    .valid     (PE20_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE20_acount[7:0]                ), //o
    .bcount    (PE20_bcount[7:0]                ), //o
    .PE_OUT    (PE20_PE_OUT[31:0]               ), //o
    .finish    (PE20_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE21 (
    .activate  (PE20_acount[7:0]                ), //i
    .weight    (PE11_bcount[7:0]                ), //i
    .valid     (PE21_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE21_acount[7:0]                ), //o
    .bcount    (PE21_bcount[7:0]                ), //o
    .PE_OUT    (PE21_PE_OUT[31:0]               ), //o
    .finish    (PE21_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE22 (
    .activate  (PE21_acount[7:0]                ), //i
    .weight    (PE12_bcount[7:0]                ), //i
    .valid     (PE22_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE22_acount[7:0]                ), //o
    .bcount    (PE22_bcount[7:0]                ), //o
    .PE_OUT    (PE22_PE_OUT[31:0]               ), //o
    .finish    (PE22_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE23 (
    .activate  (PE22_acount[7:0]                ), //i
    .weight    (PE13_bcount[7:0]                ), //i
    .valid     (PE23_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE23_acount[7:0]                ), //o
    .bcount    (PE23_bcount[7:0]                ), //o
    .PE_OUT    (PE23_PE_OUT[31:0]               ), //o
    .finish    (PE23_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE24 (
    .activate  (PE23_acount[7:0]                ), //i
    .weight    (PE14_bcount[7:0]                ), //i
    .valid     (PE24_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE24_acount[7:0]                ), //o
    .bcount    (PE24_bcount[7:0]                ), //o
    .PE_OUT    (PE24_PE_OUT[31:0]               ), //o
    .finish    (PE24_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE25 (
    .activate  (PE24_acount[7:0]                ), //i
    .weight    (PE15_bcount[7:0]                ), //i
    .valid     (PE25_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE25_acount[7:0]                ), //o
    .bcount    (PE25_bcount[7:0]                ), //o
    .PE_OUT    (PE25_PE_OUT[31:0]               ), //o
    .finish    (PE25_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE26 (
    .activate  (PE25_acount[7:0]                ), //i
    .weight    (PE16_bcount[7:0]                ), //i
    .valid     (PE26_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE26_acount[7:0]                ), //o
    .bcount    (PE26_bcount[7:0]                ), //o
    .PE_OUT    (PE26_PE_OUT[31:0]               ), //o
    .finish    (PE26_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE27 (
    .activate  (PE26_acount[7:0]                ), //i
    .weight    (PE17_bcount[7:0]                ), //i
    .valid     (PE27_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE27_acount[7:0]                ), //o
    .bcount    (PE27_bcount[7:0]                ), //o
    .PE_OUT    (PE27_PE_OUT[31:0]               ), //o
    .finish    (PE27_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE30 (
    .activate  (io_MatrixA_3[7:0]               ), //i
    .weight    (PE20_bcount[7:0]                ), //i
    .valid     (PE30_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE30_acount[7:0]                ), //o
    .bcount    (PE30_bcount[7:0]                ), //o
    .PE_OUT    (PE30_PE_OUT[31:0]               ), //o
    .finish    (PE30_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE31 (
    .activate  (PE30_acount[7:0]                ), //i
    .weight    (PE21_bcount[7:0]                ), //i
    .valid     (PE31_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE31_acount[7:0]                ), //o
    .bcount    (PE31_bcount[7:0]                ), //o
    .PE_OUT    (PE31_PE_OUT[31:0]               ), //o
    .finish    (PE31_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE32 (
    .activate  (PE31_acount[7:0]                ), //i
    .weight    (PE22_bcount[7:0]                ), //i
    .valid     (PE32_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE32_acount[7:0]                ), //o
    .bcount    (PE32_bcount[7:0]                ), //o
    .PE_OUT    (PE32_PE_OUT[31:0]               ), //o
    .finish    (PE32_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE33 (
    .activate  (PE32_acount[7:0]                ), //i
    .weight    (PE23_bcount[7:0]                ), //i
    .valid     (PE33_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE33_acount[7:0]                ), //o
    .bcount    (PE33_bcount[7:0]                ), //o
    .PE_OUT    (PE33_PE_OUT[31:0]               ), //o
    .finish    (PE33_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE34 (
    .activate  (PE33_acount[7:0]                ), //i
    .weight    (PE24_bcount[7:0]                ), //i
    .valid     (PE34_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE34_acount[7:0]                ), //o
    .bcount    (PE34_bcount[7:0]                ), //o
    .PE_OUT    (PE34_PE_OUT[31:0]               ), //o
    .finish    (PE34_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE35 (
    .activate  (PE34_acount[7:0]                ), //i
    .weight    (PE25_bcount[7:0]                ), //i
    .valid     (PE35_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE35_acount[7:0]                ), //o
    .bcount    (PE35_bcount[7:0]                ), //o
    .PE_OUT    (PE35_PE_OUT[31:0]               ), //o
    .finish    (PE35_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE36 (
    .activate  (PE35_acount[7:0]                ), //i
    .weight    (PE26_bcount[7:0]                ), //i
    .valid     (PE36_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE36_acount[7:0]                ), //o
    .bcount    (PE36_bcount[7:0]                ), //o
    .PE_OUT    (PE36_PE_OUT[31:0]               ), //o
    .finish    (PE36_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE37 (
    .activate  (PE36_acount[7:0]                ), //i
    .weight    (PE27_bcount[7:0]                ), //i
    .valid     (PE37_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE37_acount[7:0]                ), //o
    .bcount    (PE37_bcount[7:0]                ), //o
    .PE_OUT    (PE37_PE_OUT[31:0]               ), //o
    .finish    (PE37_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE40 (
    .activate  (io_MatrixA_4[7:0]               ), //i
    .weight    (PE30_bcount[7:0]                ), //i
    .valid     (PE40_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE40_acount[7:0]                ), //o
    .bcount    (PE40_bcount[7:0]                ), //o
    .PE_OUT    (PE40_PE_OUT[31:0]               ), //o
    .finish    (PE40_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE41 (
    .activate  (PE40_acount[7:0]                ), //i
    .weight    (PE31_bcount[7:0]                ), //i
    .valid     (PE41_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE41_acount[7:0]                ), //o
    .bcount    (PE41_bcount[7:0]                ), //o
    .PE_OUT    (PE41_PE_OUT[31:0]               ), //o
    .finish    (PE41_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE42 (
    .activate  (PE41_acount[7:0]                ), //i
    .weight    (PE32_bcount[7:0]                ), //i
    .valid     (PE42_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE42_acount[7:0]                ), //o
    .bcount    (PE42_bcount[7:0]                ), //o
    .PE_OUT    (PE42_PE_OUT[31:0]               ), //o
    .finish    (PE42_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE43 (
    .activate  (PE42_acount[7:0]                ), //i
    .weight    (PE33_bcount[7:0]                ), //i
    .valid     (PE43_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE43_acount[7:0]                ), //o
    .bcount    (PE43_bcount[7:0]                ), //o
    .PE_OUT    (PE43_PE_OUT[31:0]               ), //o
    .finish    (PE43_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE44 (
    .activate  (PE43_acount[7:0]                ), //i
    .weight    (PE34_bcount[7:0]                ), //i
    .valid     (PE44_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE44_acount[7:0]                ), //o
    .bcount    (PE44_bcount[7:0]                ), //o
    .PE_OUT    (PE44_PE_OUT[31:0]               ), //o
    .finish    (PE44_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE45 (
    .activate  (PE44_acount[7:0]                ), //i
    .weight    (PE35_bcount[7:0]                ), //i
    .valid     (PE45_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE45_acount[7:0]                ), //o
    .bcount    (PE45_bcount[7:0]                ), //o
    .PE_OUT    (PE45_PE_OUT[31:0]               ), //o
    .finish    (PE45_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE46 (
    .activate  (PE45_acount[7:0]                ), //i
    .weight    (PE36_bcount[7:0]                ), //i
    .valid     (PE46_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE46_acount[7:0]                ), //o
    .bcount    (PE46_bcount[7:0]                ), //o
    .PE_OUT    (PE46_PE_OUT[31:0]               ), //o
    .finish    (PE46_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE47 (
    .activate  (PE46_acount[7:0]                ), //i
    .weight    (PE37_bcount[7:0]                ), //i
    .valid     (PE47_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE47_acount[7:0]                ), //o
    .bcount    (PE47_bcount[7:0]                ), //o
    .PE_OUT    (PE47_PE_OUT[31:0]               ), //o
    .finish    (PE47_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE50 (
    .activate  (io_MatrixA_5[7:0]               ), //i
    .weight    (PE40_bcount[7:0]                ), //i
    .valid     (PE50_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE50_acount[7:0]                ), //o
    .bcount    (PE50_bcount[7:0]                ), //o
    .PE_OUT    (PE50_PE_OUT[31:0]               ), //o
    .finish    (PE50_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE51 (
    .activate  (PE50_acount[7:0]                ), //i
    .weight    (PE41_bcount[7:0]                ), //i
    .valid     (PE51_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE51_acount[7:0]                ), //o
    .bcount    (PE51_bcount[7:0]                ), //o
    .PE_OUT    (PE51_PE_OUT[31:0]               ), //o
    .finish    (PE51_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE52 (
    .activate  (PE51_acount[7:0]                ), //i
    .weight    (PE42_bcount[7:0]                ), //i
    .valid     (PE52_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE52_acount[7:0]                ), //o
    .bcount    (PE52_bcount[7:0]                ), //o
    .PE_OUT    (PE52_PE_OUT[31:0]               ), //o
    .finish    (PE52_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE53 (
    .activate  (PE52_acount[7:0]                ), //i
    .weight    (PE43_bcount[7:0]                ), //i
    .valid     (PE53_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE53_acount[7:0]                ), //o
    .bcount    (PE53_bcount[7:0]                ), //o
    .PE_OUT    (PE53_PE_OUT[31:0]               ), //o
    .finish    (PE53_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE54 (
    .activate  (PE53_acount[7:0]                ), //i
    .weight    (PE44_bcount[7:0]                ), //i
    .valid     (PE54_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE54_acount[7:0]                ), //o
    .bcount    (PE54_bcount[7:0]                ), //o
    .PE_OUT    (PE54_PE_OUT[31:0]               ), //o
    .finish    (PE54_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE55 (
    .activate  (PE54_acount[7:0]                ), //i
    .weight    (PE45_bcount[7:0]                ), //i
    .valid     (PE55_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE55_acount[7:0]                ), //o
    .bcount    (PE55_bcount[7:0]                ), //o
    .PE_OUT    (PE55_PE_OUT[31:0]               ), //o
    .finish    (PE55_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE56 (
    .activate  (PE55_acount[7:0]                ), //i
    .weight    (PE46_bcount[7:0]                ), //i
    .valid     (PE56_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE56_acount[7:0]                ), //o
    .bcount    (PE56_bcount[7:0]                ), //o
    .PE_OUT    (PE56_PE_OUT[31:0]               ), //o
    .finish    (PE56_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE57 (
    .activate  (PE56_acount[7:0]                ), //i
    .weight    (PE47_bcount[7:0]                ), //i
    .valid     (PE57_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE57_acount[7:0]                ), //o
    .bcount    (PE57_bcount[7:0]                ), //o
    .PE_OUT    (PE57_PE_OUT[31:0]               ), //o
    .finish    (PE57_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE60 (
    .activate  (io_MatrixA_6[7:0]               ), //i
    .weight    (PE50_bcount[7:0]                ), //i
    .valid     (PE60_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE60_acount[7:0]                ), //o
    .bcount    (PE60_bcount[7:0]                ), //o
    .PE_OUT    (PE60_PE_OUT[31:0]               ), //o
    .finish    (PE60_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE61 (
    .activate  (PE60_acount[7:0]                ), //i
    .weight    (PE51_bcount[7:0]                ), //i
    .valid     (PE61_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE61_acount[7:0]                ), //o
    .bcount    (PE61_bcount[7:0]                ), //o
    .PE_OUT    (PE61_PE_OUT[31:0]               ), //o
    .finish    (PE61_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE62 (
    .activate  (PE61_acount[7:0]                ), //i
    .weight    (PE52_bcount[7:0]                ), //i
    .valid     (PE62_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE62_acount[7:0]                ), //o
    .bcount    (PE62_bcount[7:0]                ), //o
    .PE_OUT    (PE62_PE_OUT[31:0]               ), //o
    .finish    (PE62_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE63 (
    .activate  (PE62_acount[7:0]                ), //i
    .weight    (PE53_bcount[7:0]                ), //i
    .valid     (PE63_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE63_acount[7:0]                ), //o
    .bcount    (PE63_bcount[7:0]                ), //o
    .PE_OUT    (PE63_PE_OUT[31:0]               ), //o
    .finish    (PE63_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE64 (
    .activate  (PE63_acount[7:0]                ), //i
    .weight    (PE54_bcount[7:0]                ), //i
    .valid     (PE64_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE64_acount[7:0]                ), //o
    .bcount    (PE64_bcount[7:0]                ), //o
    .PE_OUT    (PE64_PE_OUT[31:0]               ), //o
    .finish    (PE64_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE65 (
    .activate  (PE64_acount[7:0]                ), //i
    .weight    (PE55_bcount[7:0]                ), //i
    .valid     (PE65_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE65_acount[7:0]                ), //o
    .bcount    (PE65_bcount[7:0]                ), //o
    .PE_OUT    (PE65_PE_OUT[31:0]               ), //o
    .finish    (PE65_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE66 (
    .activate  (PE65_acount[7:0]                ), //i
    .weight    (PE56_bcount[7:0]                ), //i
    .valid     (PE66_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE66_acount[7:0]                ), //o
    .bcount    (PE66_bcount[7:0]                ), //o
    .PE_OUT    (PE66_PE_OUT[31:0]               ), //o
    .finish    (PE66_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE67 (
    .activate  (PE66_acount[7:0]                ), //i
    .weight    (PE57_bcount[7:0]                ), //i
    .valid     (PE67_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE67_acount[7:0]                ), //o
    .bcount    (PE67_bcount[7:0]                ), //o
    .PE_OUT    (PE67_PE_OUT[31:0]               ), //o
    .finish    (PE67_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE70 (
    .activate  (io_MatrixA_7[7:0]               ), //i
    .weight    (PE60_bcount[7:0]                ), //i
    .valid     (PE70_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE70_acount[7:0]                ), //o
    .bcount    (PE70_bcount[7:0]                ), //o
    .PE_OUT    (PE70_PE_OUT[31:0]               ), //o
    .finish    (PE70_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE71 (
    .activate  (PE70_acount[7:0]                ), //i
    .weight    (PE61_bcount[7:0]                ), //i
    .valid     (PE71_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE71_acount[7:0]                ), //o
    .bcount    (PE71_bcount[7:0]                ), //o
    .PE_OUT    (PE71_PE_OUT[31:0]               ), //o
    .finish    (PE71_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE72 (
    .activate  (PE71_acount[7:0]                ), //i
    .weight    (PE62_bcount[7:0]                ), //i
    .valid     (PE72_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE72_acount[7:0]                ), //o
    .bcount    (PE72_bcount[7:0]                ), //o
    .PE_OUT    (PE72_PE_OUT[31:0]               ), //o
    .finish    (PE72_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE73 (
    .activate  (PE72_acount[7:0]                ), //i
    .weight    (PE63_bcount[7:0]                ), //i
    .valid     (PE73_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE73_acount[7:0]                ), //o
    .bcount    (PE73_bcount[7:0]                ), //o
    .PE_OUT    (PE73_PE_OUT[31:0]               ), //o
    .finish    (PE73_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE74 (
    .activate  (PE73_acount[7:0]                ), //i
    .weight    (PE64_bcount[7:0]                ), //i
    .valid     (PE74_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE74_acount[7:0]                ), //o
    .bcount    (PE74_bcount[7:0]                ), //o
    .PE_OUT    (PE74_PE_OUT[31:0]               ), //o
    .finish    (PE74_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE75 (
    .activate  (PE74_acount[7:0]                ), //i
    .weight    (PE65_bcount[7:0]                ), //i
    .valid     (PE75_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE75_acount[7:0]                ), //o
    .bcount    (PE75_bcount[7:0]                ), //o
    .PE_OUT    (PE75_PE_OUT[31:0]               ), //o
    .finish    (PE75_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE76 (
    .activate  (PE75_acount[7:0]                ), //i
    .weight    (PE66_bcount[7:0]                ), //i
    .valid     (PE76_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE76_acount[7:0]                ), //o
    .bcount    (PE76_bcount[7:0]                ), //o
    .PE_OUT    (PE76_PE_OUT[31:0]               ), //o
    .finish    (PE76_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE77 (
    .activate  (PE76_acount[7:0]                ), //i
    .weight    (PE67_bcount[7:0]                ), //i
    .valid     (PE77_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE77_acount[7:0]                ), //o
    .bcount    (PE77_bcount[7:0]                ), //o
    .PE_OUT    (PE77_PE_OUT[31:0]               ), //o
    .finish    (PE77_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  always @(*) begin
    MatrixC_0 = 32'h0;
    if(PE00_finish) begin
      MatrixC_0 = PE00_PE_OUT;
    end
    if(PE01_finish) begin
      MatrixC_0 = PE01_PE_OUT;
    end
    if(PE02_finish) begin
      MatrixC_0 = PE02_PE_OUT;
    end
    if(PE03_finish) begin
      MatrixC_0 = PE03_PE_OUT;
    end
    if(PE04_finish) begin
      MatrixC_0 = PE04_PE_OUT;
    end
    if(PE05_finish) begin
      MatrixC_0 = PE05_PE_OUT;
    end
    if(PE06_finish) begin
      MatrixC_0 = PE06_PE_OUT;
    end
    if(PE07_finish) begin
      MatrixC_0 = PE07_PE_OUT;
    end
  end

  always @(*) begin
    MatrixC_1 = 32'h0;
    if(PE10_finish) begin
      MatrixC_1 = PE10_PE_OUT;
    end
    if(PE11_finish) begin
      MatrixC_1 = PE11_PE_OUT;
    end
    if(PE12_finish) begin
      MatrixC_1 = PE12_PE_OUT;
    end
    if(PE13_finish) begin
      MatrixC_1 = PE13_PE_OUT;
    end
    if(PE14_finish) begin
      MatrixC_1 = PE14_PE_OUT;
    end
    if(PE15_finish) begin
      MatrixC_1 = PE15_PE_OUT;
    end
    if(PE16_finish) begin
      MatrixC_1 = PE16_PE_OUT;
    end
    if(PE17_finish) begin
      MatrixC_1 = PE17_PE_OUT;
    end
  end

  always @(*) begin
    MatrixC_2 = 32'h0;
    if(PE20_finish) begin
      MatrixC_2 = PE20_PE_OUT;
    end
    if(PE21_finish) begin
      MatrixC_2 = PE21_PE_OUT;
    end
    if(PE22_finish) begin
      MatrixC_2 = PE22_PE_OUT;
    end
    if(PE23_finish) begin
      MatrixC_2 = PE23_PE_OUT;
    end
    if(PE24_finish) begin
      MatrixC_2 = PE24_PE_OUT;
    end
    if(PE25_finish) begin
      MatrixC_2 = PE25_PE_OUT;
    end
    if(PE26_finish) begin
      MatrixC_2 = PE26_PE_OUT;
    end
    if(PE27_finish) begin
      MatrixC_2 = PE27_PE_OUT;
    end
  end

  always @(*) begin
    MatrixC_3 = 32'h0;
    if(PE30_finish) begin
      MatrixC_3 = PE30_PE_OUT;
    end
    if(PE31_finish) begin
      MatrixC_3 = PE31_PE_OUT;
    end
    if(PE32_finish) begin
      MatrixC_3 = PE32_PE_OUT;
    end
    if(PE33_finish) begin
      MatrixC_3 = PE33_PE_OUT;
    end
    if(PE34_finish) begin
      MatrixC_3 = PE34_PE_OUT;
    end
    if(PE35_finish) begin
      MatrixC_3 = PE35_PE_OUT;
    end
    if(PE36_finish) begin
      MatrixC_3 = PE36_PE_OUT;
    end
    if(PE37_finish) begin
      MatrixC_3 = PE37_PE_OUT;
    end
  end

  always @(*) begin
    MatrixC_4 = 32'h0;
    if(PE40_finish) begin
      MatrixC_4 = PE40_PE_OUT;
    end
    if(PE41_finish) begin
      MatrixC_4 = PE41_PE_OUT;
    end
    if(PE42_finish) begin
      MatrixC_4 = PE42_PE_OUT;
    end
    if(PE43_finish) begin
      MatrixC_4 = PE43_PE_OUT;
    end
    if(PE44_finish) begin
      MatrixC_4 = PE44_PE_OUT;
    end
    if(PE45_finish) begin
      MatrixC_4 = PE45_PE_OUT;
    end
    if(PE46_finish) begin
      MatrixC_4 = PE46_PE_OUT;
    end
    if(PE47_finish) begin
      MatrixC_4 = PE47_PE_OUT;
    end
  end

  always @(*) begin
    MatrixC_5 = 32'h0;
    if(PE50_finish) begin
      MatrixC_5 = PE50_PE_OUT;
    end
    if(PE51_finish) begin
      MatrixC_5 = PE51_PE_OUT;
    end
    if(PE52_finish) begin
      MatrixC_5 = PE52_PE_OUT;
    end
    if(PE53_finish) begin
      MatrixC_5 = PE53_PE_OUT;
    end
    if(PE54_finish) begin
      MatrixC_5 = PE54_PE_OUT;
    end
    if(PE55_finish) begin
      MatrixC_5 = PE55_PE_OUT;
    end
    if(PE56_finish) begin
      MatrixC_5 = PE56_PE_OUT;
    end
    if(PE57_finish) begin
      MatrixC_5 = PE57_PE_OUT;
    end
  end

  always @(*) begin
    MatrixC_6 = 32'h0;
    if(PE60_finish) begin
      MatrixC_6 = PE60_PE_OUT;
    end
    if(PE61_finish) begin
      MatrixC_6 = PE61_PE_OUT;
    end
    if(PE62_finish) begin
      MatrixC_6 = PE62_PE_OUT;
    end
    if(PE63_finish) begin
      MatrixC_6 = PE63_PE_OUT;
    end
    if(PE64_finish) begin
      MatrixC_6 = PE64_PE_OUT;
    end
    if(PE65_finish) begin
      MatrixC_6 = PE65_PE_OUT;
    end
    if(PE66_finish) begin
      MatrixC_6 = PE66_PE_OUT;
    end
    if(PE67_finish) begin
      MatrixC_6 = PE67_PE_OUT;
    end
  end

  always @(*) begin
    MatrixC_7 = 32'h0;
    if(PE70_finish) begin
      MatrixC_7 = PE70_PE_OUT;
    end
    if(PE71_finish) begin
      MatrixC_7 = PE71_PE_OUT;
    end
    if(PE72_finish) begin
      MatrixC_7 = PE72_PE_OUT;
    end
    if(PE73_finish) begin
      MatrixC_7 = PE73_PE_OUT;
    end
    if(PE74_finish) begin
      MatrixC_7 = PE74_PE_OUT;
    end
    if(PE75_finish) begin
      MatrixC_7 = PE75_PE_OUT;
    end
    if(PE76_finish) begin
      MatrixC_7 = PE76_PE_OUT;
    end
    if(PE77_finish) begin
      MatrixC_7 = PE77_PE_OUT;
    end
  end

  assign PE00_valid = (io_A_Valid_0 && io_B_Valid_0);
  assign PE01_valid = (io_A_Valid_0_delay_1 && io_B_Valid_1);
  assign PE02_valid = (io_A_Valid_0_delay_2 && io_B_Valid_2);
  assign PE03_valid = (io_A_Valid_0_delay_3 && io_B_Valid_3);
  assign PE04_valid = (io_A_Valid_0_delay_4 && io_B_Valid_4);
  assign PE05_valid = (io_A_Valid_0_delay_5 && io_B_Valid_5);
  assign PE06_valid = (io_A_Valid_0_delay_6 && io_B_Valid_6);
  assign PE07_valid = (io_A_Valid_0_delay_7 && io_B_Valid_7);
  assign PE10_valid = (io_A_Valid_1 && io_B_Valid_0_delay_1);
  assign PE11_valid = (io_A_Valid_1_delay_1 && io_B_Valid_1_delay_1);
  assign PE12_valid = (io_A_Valid_1_delay_2 && io_B_Valid_2_delay_1);
  assign PE13_valid = (io_A_Valid_1_delay_3 && io_B_Valid_3_delay_1);
  assign PE14_valid = (io_A_Valid_1_delay_4 && io_B_Valid_4_delay_1);
  assign PE15_valid = (io_A_Valid_1_delay_5 && io_B_Valid_5_delay_1);
  assign PE16_valid = (io_A_Valid_1_delay_6 && io_B_Valid_6_delay_1);
  assign PE17_valid = (io_A_Valid_1_delay_7 && io_B_Valid_7_delay_1);
  assign PE20_valid = (io_A_Valid_2 && io_B_Valid_0_delay_2);
  assign PE21_valid = (io_A_Valid_2_delay_1 && io_B_Valid_1_delay_2);
  assign PE22_valid = (io_A_Valid_2_delay_2 && io_B_Valid_2_delay_2);
  assign PE23_valid = (io_A_Valid_2_delay_3 && io_B_Valid_3_delay_2);
  assign PE24_valid = (io_A_Valid_2_delay_4 && io_B_Valid_4_delay_2);
  assign PE25_valid = (io_A_Valid_2_delay_5 && io_B_Valid_5_delay_2);
  assign PE26_valid = (io_A_Valid_2_delay_6 && io_B_Valid_6_delay_2);
  assign PE27_valid = (io_A_Valid_2_delay_7 && io_B_Valid_7_delay_2);
  assign PE30_valid = (io_A_Valid_3 && io_B_Valid_0_delay_3);
  assign PE31_valid = (io_A_Valid_3_delay_1 && io_B_Valid_1_delay_3);
  assign PE32_valid = (io_A_Valid_3_delay_2 && io_B_Valid_2_delay_3);
  assign PE33_valid = (io_A_Valid_3_delay_3 && io_B_Valid_3_delay_3);
  assign PE34_valid = (io_A_Valid_3_delay_4 && io_B_Valid_4_delay_3);
  assign PE35_valid = (io_A_Valid_3_delay_5 && io_B_Valid_5_delay_3);
  assign PE36_valid = (io_A_Valid_3_delay_6 && io_B_Valid_6_delay_3);
  assign PE37_valid = (io_A_Valid_3_delay_7 && io_B_Valid_7_delay_3);
  assign PE40_valid = (io_A_Valid_4 && io_B_Valid_0_delay_4);
  assign PE41_valid = (io_A_Valid_4_delay_1 && io_B_Valid_1_delay_4);
  assign PE42_valid = (io_A_Valid_4_delay_2 && io_B_Valid_2_delay_4);
  assign PE43_valid = (io_A_Valid_4_delay_3 && io_B_Valid_3_delay_4);
  assign PE44_valid = (io_A_Valid_4_delay_4 && io_B_Valid_4_delay_4);
  assign PE45_valid = (io_A_Valid_4_delay_5 && io_B_Valid_5_delay_4);
  assign PE46_valid = (io_A_Valid_4_delay_6 && io_B_Valid_6_delay_4);
  assign PE47_valid = (io_A_Valid_4_delay_7 && io_B_Valid_7_delay_4);
  assign PE50_valid = (io_A_Valid_5 && io_B_Valid_0_delay_5);
  assign PE51_valid = (io_A_Valid_5_delay_1 && io_B_Valid_1_delay_5);
  assign PE52_valid = (io_A_Valid_5_delay_2 && io_B_Valid_2_delay_5);
  assign PE53_valid = (io_A_Valid_5_delay_3 && io_B_Valid_3_delay_5);
  assign PE54_valid = (io_A_Valid_5_delay_4 && io_B_Valid_4_delay_5);
  assign PE55_valid = (io_A_Valid_5_delay_5 && io_B_Valid_5_delay_5);
  assign PE56_valid = (io_A_Valid_5_delay_6 && io_B_Valid_6_delay_5);
  assign PE57_valid = (io_A_Valid_5_delay_7 && io_B_Valid_7_delay_5);
  assign PE60_valid = (io_A_Valid_6 && io_B_Valid_0_delay_6);
  assign PE61_valid = (io_A_Valid_6_delay_1 && io_B_Valid_1_delay_6);
  assign PE62_valid = (io_A_Valid_6_delay_2 && io_B_Valid_2_delay_6);
  assign PE63_valid = (io_A_Valid_6_delay_3 && io_B_Valid_3_delay_6);
  assign PE64_valid = (io_A_Valid_6_delay_4 && io_B_Valid_4_delay_6);
  assign PE65_valid = (io_A_Valid_6_delay_5 && io_B_Valid_5_delay_6);
  assign PE66_valid = (io_A_Valid_6_delay_6 && io_B_Valid_6_delay_6);
  assign PE67_valid = (io_A_Valid_6_delay_7 && io_B_Valid_7_delay_6);
  assign PE70_valid = (io_A_Valid_7 && io_B_Valid_0_delay_7);
  assign PE71_valid = (io_A_Valid_7_delay_1 && io_B_Valid_1_delay_7);
  assign PE72_valid = (io_A_Valid_7_delay_2 && io_B_Valid_2_delay_7);
  assign PE73_valid = (io_A_Valid_7_delay_3 && io_B_Valid_3_delay_7);
  assign PE74_valid = (io_A_Valid_7_delay_4 && io_B_Valid_4_delay_7);
  assign PE75_valid = (io_A_Valid_7_delay_5 && io_B_Valid_5_delay_7);
  assign PE76_valid = (io_A_Valid_7_delay_6 && io_B_Valid_6_delay_7);
  assign PE77_valid = (io_A_Valid_7_delay_7 && io_B_Valid_7_delay_7);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      io_signCount_regNextWhen <= 16'h0;
      io_signCount_regNextWhen_1 <= 16'h0;
      io_signCount_regNextWhen_2 <= 16'h0;
      io_signCount_regNextWhen_3 <= 16'h0;
      io_signCount_regNextWhen_4 <= 16'h0;
      io_signCount_regNextWhen_5 <= 16'h0;
      io_signCount_regNextWhen_6 <= 16'h0;
      io_signCount_regNextWhen_7 <= 16'h0;
    end else begin
      if(start) begin
        io_signCount_regNextWhen <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_1 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_2 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_3 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_4 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_5 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_6 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_7 <= io_signCount;
      end
    end
  end

  always @(posedge clk) begin
    io_A_Valid_0_delay_1 <= io_A_Valid_0;
    io_A_Valid_0_delay_1_1 <= io_A_Valid_0;
    io_A_Valid_0_delay_2 <= io_A_Valid_0_delay_1_1;
    io_A_Valid_0_delay_1_2 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_1 <= io_A_Valid_0_delay_1_2;
    io_A_Valid_0_delay_3 <= io_A_Valid_0_delay_2_1;
    io_A_Valid_0_delay_1_3 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_2 <= io_A_Valid_0_delay_1_3;
    io_A_Valid_0_delay_3_1 <= io_A_Valid_0_delay_2_2;
    io_A_Valid_0_delay_4 <= io_A_Valid_0_delay_3_1;
    io_A_Valid_0_delay_1_4 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_3 <= io_A_Valid_0_delay_1_4;
    io_A_Valid_0_delay_3_2 <= io_A_Valid_0_delay_2_3;
    io_A_Valid_0_delay_4_1 <= io_A_Valid_0_delay_3_2;
    io_A_Valid_0_delay_5 <= io_A_Valid_0_delay_4_1;
    io_A_Valid_0_delay_1_5 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_4 <= io_A_Valid_0_delay_1_5;
    io_A_Valid_0_delay_3_3 <= io_A_Valid_0_delay_2_4;
    io_A_Valid_0_delay_4_2 <= io_A_Valid_0_delay_3_3;
    io_A_Valid_0_delay_5_1 <= io_A_Valid_0_delay_4_2;
    io_A_Valid_0_delay_6 <= io_A_Valid_0_delay_5_1;
    io_A_Valid_0_delay_1_6 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_5 <= io_A_Valid_0_delay_1_6;
    io_A_Valid_0_delay_3_4 <= io_A_Valid_0_delay_2_5;
    io_A_Valid_0_delay_4_3 <= io_A_Valid_0_delay_3_4;
    io_A_Valid_0_delay_5_2 <= io_A_Valid_0_delay_4_3;
    io_A_Valid_0_delay_6_1 <= io_A_Valid_0_delay_5_2;
    io_A_Valid_0_delay_7 <= io_A_Valid_0_delay_6_1;
    io_B_Valid_0_delay_1 <= io_B_Valid_0;
    io_A_Valid_1_delay_1 <= io_A_Valid_1;
    io_B_Valid_1_delay_1 <= io_B_Valid_1;
    io_A_Valid_1_delay_1_1 <= io_A_Valid_1;
    io_A_Valid_1_delay_2 <= io_A_Valid_1_delay_1_1;
    io_B_Valid_2_delay_1 <= io_B_Valid_2;
    io_A_Valid_1_delay_1_2 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_1 <= io_A_Valid_1_delay_1_2;
    io_A_Valid_1_delay_3 <= io_A_Valid_1_delay_2_1;
    io_B_Valid_3_delay_1 <= io_B_Valid_3;
    io_A_Valid_1_delay_1_3 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_2 <= io_A_Valid_1_delay_1_3;
    io_A_Valid_1_delay_3_1 <= io_A_Valid_1_delay_2_2;
    io_A_Valid_1_delay_4 <= io_A_Valid_1_delay_3_1;
    io_B_Valid_4_delay_1 <= io_B_Valid_4;
    io_A_Valid_1_delay_1_4 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_3 <= io_A_Valid_1_delay_1_4;
    io_A_Valid_1_delay_3_2 <= io_A_Valid_1_delay_2_3;
    io_A_Valid_1_delay_4_1 <= io_A_Valid_1_delay_3_2;
    io_A_Valid_1_delay_5 <= io_A_Valid_1_delay_4_1;
    io_B_Valid_5_delay_1 <= io_B_Valid_5;
    io_A_Valid_1_delay_1_5 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_4 <= io_A_Valid_1_delay_1_5;
    io_A_Valid_1_delay_3_3 <= io_A_Valid_1_delay_2_4;
    io_A_Valid_1_delay_4_2 <= io_A_Valid_1_delay_3_3;
    io_A_Valid_1_delay_5_1 <= io_A_Valid_1_delay_4_2;
    io_A_Valid_1_delay_6 <= io_A_Valid_1_delay_5_1;
    io_B_Valid_6_delay_1 <= io_B_Valid_6;
    io_A_Valid_1_delay_1_6 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_5 <= io_A_Valid_1_delay_1_6;
    io_A_Valid_1_delay_3_4 <= io_A_Valid_1_delay_2_5;
    io_A_Valid_1_delay_4_3 <= io_A_Valid_1_delay_3_4;
    io_A_Valid_1_delay_5_2 <= io_A_Valid_1_delay_4_3;
    io_A_Valid_1_delay_6_1 <= io_A_Valid_1_delay_5_2;
    io_A_Valid_1_delay_7 <= io_A_Valid_1_delay_6_1;
    io_B_Valid_7_delay_1 <= io_B_Valid_7;
    io_B_Valid_0_delay_1_1 <= io_B_Valid_0;
    io_B_Valid_0_delay_2 <= io_B_Valid_0_delay_1_1;
    io_A_Valid_2_delay_1 <= io_A_Valid_2;
    io_B_Valid_1_delay_1_1 <= io_B_Valid_1;
    io_B_Valid_1_delay_2 <= io_B_Valid_1_delay_1_1;
    io_A_Valid_2_delay_1_1 <= io_A_Valid_2;
    io_A_Valid_2_delay_2 <= io_A_Valid_2_delay_1_1;
    io_B_Valid_2_delay_1_1 <= io_B_Valid_2;
    io_B_Valid_2_delay_2 <= io_B_Valid_2_delay_1_1;
    io_A_Valid_2_delay_1_2 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_1 <= io_A_Valid_2_delay_1_2;
    io_A_Valid_2_delay_3 <= io_A_Valid_2_delay_2_1;
    io_B_Valid_3_delay_1_1 <= io_B_Valid_3;
    io_B_Valid_3_delay_2 <= io_B_Valid_3_delay_1_1;
    io_A_Valid_2_delay_1_3 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_2 <= io_A_Valid_2_delay_1_3;
    io_A_Valid_2_delay_3_1 <= io_A_Valid_2_delay_2_2;
    io_A_Valid_2_delay_4 <= io_A_Valid_2_delay_3_1;
    io_B_Valid_4_delay_1_1 <= io_B_Valid_4;
    io_B_Valid_4_delay_2 <= io_B_Valid_4_delay_1_1;
    io_A_Valid_2_delay_1_4 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_3 <= io_A_Valid_2_delay_1_4;
    io_A_Valid_2_delay_3_2 <= io_A_Valid_2_delay_2_3;
    io_A_Valid_2_delay_4_1 <= io_A_Valid_2_delay_3_2;
    io_A_Valid_2_delay_5 <= io_A_Valid_2_delay_4_1;
    io_B_Valid_5_delay_1_1 <= io_B_Valid_5;
    io_B_Valid_5_delay_2 <= io_B_Valid_5_delay_1_1;
    io_A_Valid_2_delay_1_5 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_4 <= io_A_Valid_2_delay_1_5;
    io_A_Valid_2_delay_3_3 <= io_A_Valid_2_delay_2_4;
    io_A_Valid_2_delay_4_2 <= io_A_Valid_2_delay_3_3;
    io_A_Valid_2_delay_5_1 <= io_A_Valid_2_delay_4_2;
    io_A_Valid_2_delay_6 <= io_A_Valid_2_delay_5_1;
    io_B_Valid_6_delay_1_1 <= io_B_Valid_6;
    io_B_Valid_6_delay_2 <= io_B_Valid_6_delay_1_1;
    io_A_Valid_2_delay_1_6 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_5 <= io_A_Valid_2_delay_1_6;
    io_A_Valid_2_delay_3_4 <= io_A_Valid_2_delay_2_5;
    io_A_Valid_2_delay_4_3 <= io_A_Valid_2_delay_3_4;
    io_A_Valid_2_delay_5_2 <= io_A_Valid_2_delay_4_3;
    io_A_Valid_2_delay_6_1 <= io_A_Valid_2_delay_5_2;
    io_A_Valid_2_delay_7 <= io_A_Valid_2_delay_6_1;
    io_B_Valid_7_delay_1_1 <= io_B_Valid_7;
    io_B_Valid_7_delay_2 <= io_B_Valid_7_delay_1_1;
    io_B_Valid_0_delay_1_2 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_1 <= io_B_Valid_0_delay_1_2;
    io_B_Valid_0_delay_3 <= io_B_Valid_0_delay_2_1;
    io_A_Valid_3_delay_1 <= io_A_Valid_3;
    io_B_Valid_1_delay_1_2 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_1 <= io_B_Valid_1_delay_1_2;
    io_B_Valid_1_delay_3 <= io_B_Valid_1_delay_2_1;
    io_A_Valid_3_delay_1_1 <= io_A_Valid_3;
    io_A_Valid_3_delay_2 <= io_A_Valid_3_delay_1_1;
    io_B_Valid_2_delay_1_2 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_1 <= io_B_Valid_2_delay_1_2;
    io_B_Valid_2_delay_3 <= io_B_Valid_2_delay_2_1;
    io_A_Valid_3_delay_1_2 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_1 <= io_A_Valid_3_delay_1_2;
    io_A_Valid_3_delay_3 <= io_A_Valid_3_delay_2_1;
    io_B_Valid_3_delay_1_2 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_1 <= io_B_Valid_3_delay_1_2;
    io_B_Valid_3_delay_3 <= io_B_Valid_3_delay_2_1;
    io_A_Valid_3_delay_1_3 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_2 <= io_A_Valid_3_delay_1_3;
    io_A_Valid_3_delay_3_1 <= io_A_Valid_3_delay_2_2;
    io_A_Valid_3_delay_4 <= io_A_Valid_3_delay_3_1;
    io_B_Valid_4_delay_1_2 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_1 <= io_B_Valid_4_delay_1_2;
    io_B_Valid_4_delay_3 <= io_B_Valid_4_delay_2_1;
    io_A_Valid_3_delay_1_4 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_3 <= io_A_Valid_3_delay_1_4;
    io_A_Valid_3_delay_3_2 <= io_A_Valid_3_delay_2_3;
    io_A_Valid_3_delay_4_1 <= io_A_Valid_3_delay_3_2;
    io_A_Valid_3_delay_5 <= io_A_Valid_3_delay_4_1;
    io_B_Valid_5_delay_1_2 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_1 <= io_B_Valid_5_delay_1_2;
    io_B_Valid_5_delay_3 <= io_B_Valid_5_delay_2_1;
    io_A_Valid_3_delay_1_5 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_4 <= io_A_Valid_3_delay_1_5;
    io_A_Valid_3_delay_3_3 <= io_A_Valid_3_delay_2_4;
    io_A_Valid_3_delay_4_2 <= io_A_Valid_3_delay_3_3;
    io_A_Valid_3_delay_5_1 <= io_A_Valid_3_delay_4_2;
    io_A_Valid_3_delay_6 <= io_A_Valid_3_delay_5_1;
    io_B_Valid_6_delay_1_2 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_1 <= io_B_Valid_6_delay_1_2;
    io_B_Valid_6_delay_3 <= io_B_Valid_6_delay_2_1;
    io_A_Valid_3_delay_1_6 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_5 <= io_A_Valid_3_delay_1_6;
    io_A_Valid_3_delay_3_4 <= io_A_Valid_3_delay_2_5;
    io_A_Valid_3_delay_4_3 <= io_A_Valid_3_delay_3_4;
    io_A_Valid_3_delay_5_2 <= io_A_Valid_3_delay_4_3;
    io_A_Valid_3_delay_6_1 <= io_A_Valid_3_delay_5_2;
    io_A_Valid_3_delay_7 <= io_A_Valid_3_delay_6_1;
    io_B_Valid_7_delay_1_2 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_1 <= io_B_Valid_7_delay_1_2;
    io_B_Valid_7_delay_3 <= io_B_Valid_7_delay_2_1;
    io_B_Valid_0_delay_1_3 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_2 <= io_B_Valid_0_delay_1_3;
    io_B_Valid_0_delay_3_1 <= io_B_Valid_0_delay_2_2;
    io_B_Valid_0_delay_4 <= io_B_Valid_0_delay_3_1;
    io_A_Valid_4_delay_1 <= io_A_Valid_4;
    io_B_Valid_1_delay_1_3 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_2 <= io_B_Valid_1_delay_1_3;
    io_B_Valid_1_delay_3_1 <= io_B_Valid_1_delay_2_2;
    io_B_Valid_1_delay_4 <= io_B_Valid_1_delay_3_1;
    io_A_Valid_4_delay_1_1 <= io_A_Valid_4;
    io_A_Valid_4_delay_2 <= io_A_Valid_4_delay_1_1;
    io_B_Valid_2_delay_1_3 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_2 <= io_B_Valid_2_delay_1_3;
    io_B_Valid_2_delay_3_1 <= io_B_Valid_2_delay_2_2;
    io_B_Valid_2_delay_4 <= io_B_Valid_2_delay_3_1;
    io_A_Valid_4_delay_1_2 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_1 <= io_A_Valid_4_delay_1_2;
    io_A_Valid_4_delay_3 <= io_A_Valid_4_delay_2_1;
    io_B_Valid_3_delay_1_3 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_2 <= io_B_Valid_3_delay_1_3;
    io_B_Valid_3_delay_3_1 <= io_B_Valid_3_delay_2_2;
    io_B_Valid_3_delay_4 <= io_B_Valid_3_delay_3_1;
    io_A_Valid_4_delay_1_3 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_2 <= io_A_Valid_4_delay_1_3;
    io_A_Valid_4_delay_3_1 <= io_A_Valid_4_delay_2_2;
    io_A_Valid_4_delay_4 <= io_A_Valid_4_delay_3_1;
    io_B_Valid_4_delay_1_3 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_2 <= io_B_Valid_4_delay_1_3;
    io_B_Valid_4_delay_3_1 <= io_B_Valid_4_delay_2_2;
    io_B_Valid_4_delay_4 <= io_B_Valid_4_delay_3_1;
    io_A_Valid_4_delay_1_4 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_3 <= io_A_Valid_4_delay_1_4;
    io_A_Valid_4_delay_3_2 <= io_A_Valid_4_delay_2_3;
    io_A_Valid_4_delay_4_1 <= io_A_Valid_4_delay_3_2;
    io_A_Valid_4_delay_5 <= io_A_Valid_4_delay_4_1;
    io_B_Valid_5_delay_1_3 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_2 <= io_B_Valid_5_delay_1_3;
    io_B_Valid_5_delay_3_1 <= io_B_Valid_5_delay_2_2;
    io_B_Valid_5_delay_4 <= io_B_Valid_5_delay_3_1;
    io_A_Valid_4_delay_1_5 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_4 <= io_A_Valid_4_delay_1_5;
    io_A_Valid_4_delay_3_3 <= io_A_Valid_4_delay_2_4;
    io_A_Valid_4_delay_4_2 <= io_A_Valid_4_delay_3_3;
    io_A_Valid_4_delay_5_1 <= io_A_Valid_4_delay_4_2;
    io_A_Valid_4_delay_6 <= io_A_Valid_4_delay_5_1;
    io_B_Valid_6_delay_1_3 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_2 <= io_B_Valid_6_delay_1_3;
    io_B_Valid_6_delay_3_1 <= io_B_Valid_6_delay_2_2;
    io_B_Valid_6_delay_4 <= io_B_Valid_6_delay_3_1;
    io_A_Valid_4_delay_1_6 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_5 <= io_A_Valid_4_delay_1_6;
    io_A_Valid_4_delay_3_4 <= io_A_Valid_4_delay_2_5;
    io_A_Valid_4_delay_4_3 <= io_A_Valid_4_delay_3_4;
    io_A_Valid_4_delay_5_2 <= io_A_Valid_4_delay_4_3;
    io_A_Valid_4_delay_6_1 <= io_A_Valid_4_delay_5_2;
    io_A_Valid_4_delay_7 <= io_A_Valid_4_delay_6_1;
    io_B_Valid_7_delay_1_3 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_2 <= io_B_Valid_7_delay_1_3;
    io_B_Valid_7_delay_3_1 <= io_B_Valid_7_delay_2_2;
    io_B_Valid_7_delay_4 <= io_B_Valid_7_delay_3_1;
    io_B_Valid_0_delay_1_4 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_3 <= io_B_Valid_0_delay_1_4;
    io_B_Valid_0_delay_3_2 <= io_B_Valid_0_delay_2_3;
    io_B_Valid_0_delay_4_1 <= io_B_Valid_0_delay_3_2;
    io_B_Valid_0_delay_5 <= io_B_Valid_0_delay_4_1;
    io_A_Valid_5_delay_1 <= io_A_Valid_5;
    io_B_Valid_1_delay_1_4 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_3 <= io_B_Valid_1_delay_1_4;
    io_B_Valid_1_delay_3_2 <= io_B_Valid_1_delay_2_3;
    io_B_Valid_1_delay_4_1 <= io_B_Valid_1_delay_3_2;
    io_B_Valid_1_delay_5 <= io_B_Valid_1_delay_4_1;
    io_A_Valid_5_delay_1_1 <= io_A_Valid_5;
    io_A_Valid_5_delay_2 <= io_A_Valid_5_delay_1_1;
    io_B_Valid_2_delay_1_4 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_3 <= io_B_Valid_2_delay_1_4;
    io_B_Valid_2_delay_3_2 <= io_B_Valid_2_delay_2_3;
    io_B_Valid_2_delay_4_1 <= io_B_Valid_2_delay_3_2;
    io_B_Valid_2_delay_5 <= io_B_Valid_2_delay_4_1;
    io_A_Valid_5_delay_1_2 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_1 <= io_A_Valid_5_delay_1_2;
    io_A_Valid_5_delay_3 <= io_A_Valid_5_delay_2_1;
    io_B_Valid_3_delay_1_4 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_3 <= io_B_Valid_3_delay_1_4;
    io_B_Valid_3_delay_3_2 <= io_B_Valid_3_delay_2_3;
    io_B_Valid_3_delay_4_1 <= io_B_Valid_3_delay_3_2;
    io_B_Valid_3_delay_5 <= io_B_Valid_3_delay_4_1;
    io_A_Valid_5_delay_1_3 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_2 <= io_A_Valid_5_delay_1_3;
    io_A_Valid_5_delay_3_1 <= io_A_Valid_5_delay_2_2;
    io_A_Valid_5_delay_4 <= io_A_Valid_5_delay_3_1;
    io_B_Valid_4_delay_1_4 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_3 <= io_B_Valid_4_delay_1_4;
    io_B_Valid_4_delay_3_2 <= io_B_Valid_4_delay_2_3;
    io_B_Valid_4_delay_4_1 <= io_B_Valid_4_delay_3_2;
    io_B_Valid_4_delay_5 <= io_B_Valid_4_delay_4_1;
    io_A_Valid_5_delay_1_4 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_3 <= io_A_Valid_5_delay_1_4;
    io_A_Valid_5_delay_3_2 <= io_A_Valid_5_delay_2_3;
    io_A_Valid_5_delay_4_1 <= io_A_Valid_5_delay_3_2;
    io_A_Valid_5_delay_5 <= io_A_Valid_5_delay_4_1;
    io_B_Valid_5_delay_1_4 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_3 <= io_B_Valid_5_delay_1_4;
    io_B_Valid_5_delay_3_2 <= io_B_Valid_5_delay_2_3;
    io_B_Valid_5_delay_4_1 <= io_B_Valid_5_delay_3_2;
    io_B_Valid_5_delay_5 <= io_B_Valid_5_delay_4_1;
    io_A_Valid_5_delay_1_5 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_4 <= io_A_Valid_5_delay_1_5;
    io_A_Valid_5_delay_3_3 <= io_A_Valid_5_delay_2_4;
    io_A_Valid_5_delay_4_2 <= io_A_Valid_5_delay_3_3;
    io_A_Valid_5_delay_5_1 <= io_A_Valid_5_delay_4_2;
    io_A_Valid_5_delay_6 <= io_A_Valid_5_delay_5_1;
    io_B_Valid_6_delay_1_4 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_3 <= io_B_Valid_6_delay_1_4;
    io_B_Valid_6_delay_3_2 <= io_B_Valid_6_delay_2_3;
    io_B_Valid_6_delay_4_1 <= io_B_Valid_6_delay_3_2;
    io_B_Valid_6_delay_5 <= io_B_Valid_6_delay_4_1;
    io_A_Valid_5_delay_1_6 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_5 <= io_A_Valid_5_delay_1_6;
    io_A_Valid_5_delay_3_4 <= io_A_Valid_5_delay_2_5;
    io_A_Valid_5_delay_4_3 <= io_A_Valid_5_delay_3_4;
    io_A_Valid_5_delay_5_2 <= io_A_Valid_5_delay_4_3;
    io_A_Valid_5_delay_6_1 <= io_A_Valid_5_delay_5_2;
    io_A_Valid_5_delay_7 <= io_A_Valid_5_delay_6_1;
    io_B_Valid_7_delay_1_4 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_3 <= io_B_Valid_7_delay_1_4;
    io_B_Valid_7_delay_3_2 <= io_B_Valid_7_delay_2_3;
    io_B_Valid_7_delay_4_1 <= io_B_Valid_7_delay_3_2;
    io_B_Valid_7_delay_5 <= io_B_Valid_7_delay_4_1;
    io_B_Valid_0_delay_1_5 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_4 <= io_B_Valid_0_delay_1_5;
    io_B_Valid_0_delay_3_3 <= io_B_Valid_0_delay_2_4;
    io_B_Valid_0_delay_4_2 <= io_B_Valid_0_delay_3_3;
    io_B_Valid_0_delay_5_1 <= io_B_Valid_0_delay_4_2;
    io_B_Valid_0_delay_6 <= io_B_Valid_0_delay_5_1;
    io_A_Valid_6_delay_1 <= io_A_Valid_6;
    io_B_Valid_1_delay_1_5 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_4 <= io_B_Valid_1_delay_1_5;
    io_B_Valid_1_delay_3_3 <= io_B_Valid_1_delay_2_4;
    io_B_Valid_1_delay_4_2 <= io_B_Valid_1_delay_3_3;
    io_B_Valid_1_delay_5_1 <= io_B_Valid_1_delay_4_2;
    io_B_Valid_1_delay_6 <= io_B_Valid_1_delay_5_1;
    io_A_Valid_6_delay_1_1 <= io_A_Valid_6;
    io_A_Valid_6_delay_2 <= io_A_Valid_6_delay_1_1;
    io_B_Valid_2_delay_1_5 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_4 <= io_B_Valid_2_delay_1_5;
    io_B_Valid_2_delay_3_3 <= io_B_Valid_2_delay_2_4;
    io_B_Valid_2_delay_4_2 <= io_B_Valid_2_delay_3_3;
    io_B_Valid_2_delay_5_1 <= io_B_Valid_2_delay_4_2;
    io_B_Valid_2_delay_6 <= io_B_Valid_2_delay_5_1;
    io_A_Valid_6_delay_1_2 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_1 <= io_A_Valid_6_delay_1_2;
    io_A_Valid_6_delay_3 <= io_A_Valid_6_delay_2_1;
    io_B_Valid_3_delay_1_5 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_4 <= io_B_Valid_3_delay_1_5;
    io_B_Valid_3_delay_3_3 <= io_B_Valid_3_delay_2_4;
    io_B_Valid_3_delay_4_2 <= io_B_Valid_3_delay_3_3;
    io_B_Valid_3_delay_5_1 <= io_B_Valid_3_delay_4_2;
    io_B_Valid_3_delay_6 <= io_B_Valid_3_delay_5_1;
    io_A_Valid_6_delay_1_3 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_2 <= io_A_Valid_6_delay_1_3;
    io_A_Valid_6_delay_3_1 <= io_A_Valid_6_delay_2_2;
    io_A_Valid_6_delay_4 <= io_A_Valid_6_delay_3_1;
    io_B_Valid_4_delay_1_5 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_4 <= io_B_Valid_4_delay_1_5;
    io_B_Valid_4_delay_3_3 <= io_B_Valid_4_delay_2_4;
    io_B_Valid_4_delay_4_2 <= io_B_Valid_4_delay_3_3;
    io_B_Valid_4_delay_5_1 <= io_B_Valid_4_delay_4_2;
    io_B_Valid_4_delay_6 <= io_B_Valid_4_delay_5_1;
    io_A_Valid_6_delay_1_4 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_3 <= io_A_Valid_6_delay_1_4;
    io_A_Valid_6_delay_3_2 <= io_A_Valid_6_delay_2_3;
    io_A_Valid_6_delay_4_1 <= io_A_Valid_6_delay_3_2;
    io_A_Valid_6_delay_5 <= io_A_Valid_6_delay_4_1;
    io_B_Valid_5_delay_1_5 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_4 <= io_B_Valid_5_delay_1_5;
    io_B_Valid_5_delay_3_3 <= io_B_Valid_5_delay_2_4;
    io_B_Valid_5_delay_4_2 <= io_B_Valid_5_delay_3_3;
    io_B_Valid_5_delay_5_1 <= io_B_Valid_5_delay_4_2;
    io_B_Valid_5_delay_6 <= io_B_Valid_5_delay_5_1;
    io_A_Valid_6_delay_1_5 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_4 <= io_A_Valid_6_delay_1_5;
    io_A_Valid_6_delay_3_3 <= io_A_Valid_6_delay_2_4;
    io_A_Valid_6_delay_4_2 <= io_A_Valid_6_delay_3_3;
    io_A_Valid_6_delay_5_1 <= io_A_Valid_6_delay_4_2;
    io_A_Valid_6_delay_6 <= io_A_Valid_6_delay_5_1;
    io_B_Valid_6_delay_1_5 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_4 <= io_B_Valid_6_delay_1_5;
    io_B_Valid_6_delay_3_3 <= io_B_Valid_6_delay_2_4;
    io_B_Valid_6_delay_4_2 <= io_B_Valid_6_delay_3_3;
    io_B_Valid_6_delay_5_1 <= io_B_Valid_6_delay_4_2;
    io_B_Valid_6_delay_6 <= io_B_Valid_6_delay_5_1;
    io_A_Valid_6_delay_1_6 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_5 <= io_A_Valid_6_delay_1_6;
    io_A_Valid_6_delay_3_4 <= io_A_Valid_6_delay_2_5;
    io_A_Valid_6_delay_4_3 <= io_A_Valid_6_delay_3_4;
    io_A_Valid_6_delay_5_2 <= io_A_Valid_6_delay_4_3;
    io_A_Valid_6_delay_6_1 <= io_A_Valid_6_delay_5_2;
    io_A_Valid_6_delay_7 <= io_A_Valid_6_delay_6_1;
    io_B_Valid_7_delay_1_5 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_4 <= io_B_Valid_7_delay_1_5;
    io_B_Valid_7_delay_3_3 <= io_B_Valid_7_delay_2_4;
    io_B_Valid_7_delay_4_2 <= io_B_Valid_7_delay_3_3;
    io_B_Valid_7_delay_5_1 <= io_B_Valid_7_delay_4_2;
    io_B_Valid_7_delay_6 <= io_B_Valid_7_delay_5_1;
    io_B_Valid_0_delay_1_6 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_5 <= io_B_Valid_0_delay_1_6;
    io_B_Valid_0_delay_3_4 <= io_B_Valid_0_delay_2_5;
    io_B_Valid_0_delay_4_3 <= io_B_Valid_0_delay_3_4;
    io_B_Valid_0_delay_5_2 <= io_B_Valid_0_delay_4_3;
    io_B_Valid_0_delay_6_1 <= io_B_Valid_0_delay_5_2;
    io_B_Valid_0_delay_7 <= io_B_Valid_0_delay_6_1;
    io_A_Valid_7_delay_1 <= io_A_Valid_7;
    io_B_Valid_1_delay_1_6 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_5 <= io_B_Valid_1_delay_1_6;
    io_B_Valid_1_delay_3_4 <= io_B_Valid_1_delay_2_5;
    io_B_Valid_1_delay_4_3 <= io_B_Valid_1_delay_3_4;
    io_B_Valid_1_delay_5_2 <= io_B_Valid_1_delay_4_3;
    io_B_Valid_1_delay_6_1 <= io_B_Valid_1_delay_5_2;
    io_B_Valid_1_delay_7 <= io_B_Valid_1_delay_6_1;
    io_A_Valid_7_delay_1_1 <= io_A_Valid_7;
    io_A_Valid_7_delay_2 <= io_A_Valid_7_delay_1_1;
    io_B_Valid_2_delay_1_6 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_5 <= io_B_Valid_2_delay_1_6;
    io_B_Valid_2_delay_3_4 <= io_B_Valid_2_delay_2_5;
    io_B_Valid_2_delay_4_3 <= io_B_Valid_2_delay_3_4;
    io_B_Valid_2_delay_5_2 <= io_B_Valid_2_delay_4_3;
    io_B_Valid_2_delay_6_1 <= io_B_Valid_2_delay_5_2;
    io_B_Valid_2_delay_7 <= io_B_Valid_2_delay_6_1;
    io_A_Valid_7_delay_1_2 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_1 <= io_A_Valid_7_delay_1_2;
    io_A_Valid_7_delay_3 <= io_A_Valid_7_delay_2_1;
    io_B_Valid_3_delay_1_6 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_5 <= io_B_Valid_3_delay_1_6;
    io_B_Valid_3_delay_3_4 <= io_B_Valid_3_delay_2_5;
    io_B_Valid_3_delay_4_3 <= io_B_Valid_3_delay_3_4;
    io_B_Valid_3_delay_5_2 <= io_B_Valid_3_delay_4_3;
    io_B_Valid_3_delay_6_1 <= io_B_Valid_3_delay_5_2;
    io_B_Valid_3_delay_7 <= io_B_Valid_3_delay_6_1;
    io_A_Valid_7_delay_1_3 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_2 <= io_A_Valid_7_delay_1_3;
    io_A_Valid_7_delay_3_1 <= io_A_Valid_7_delay_2_2;
    io_A_Valid_7_delay_4 <= io_A_Valid_7_delay_3_1;
    io_B_Valid_4_delay_1_6 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_5 <= io_B_Valid_4_delay_1_6;
    io_B_Valid_4_delay_3_4 <= io_B_Valid_4_delay_2_5;
    io_B_Valid_4_delay_4_3 <= io_B_Valid_4_delay_3_4;
    io_B_Valid_4_delay_5_2 <= io_B_Valid_4_delay_4_3;
    io_B_Valid_4_delay_6_1 <= io_B_Valid_4_delay_5_2;
    io_B_Valid_4_delay_7 <= io_B_Valid_4_delay_6_1;
    io_A_Valid_7_delay_1_4 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_3 <= io_A_Valid_7_delay_1_4;
    io_A_Valid_7_delay_3_2 <= io_A_Valid_7_delay_2_3;
    io_A_Valid_7_delay_4_1 <= io_A_Valid_7_delay_3_2;
    io_A_Valid_7_delay_5 <= io_A_Valid_7_delay_4_1;
    io_B_Valid_5_delay_1_6 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_5 <= io_B_Valid_5_delay_1_6;
    io_B_Valid_5_delay_3_4 <= io_B_Valid_5_delay_2_5;
    io_B_Valid_5_delay_4_3 <= io_B_Valid_5_delay_3_4;
    io_B_Valid_5_delay_5_2 <= io_B_Valid_5_delay_4_3;
    io_B_Valid_5_delay_6_1 <= io_B_Valid_5_delay_5_2;
    io_B_Valid_5_delay_7 <= io_B_Valid_5_delay_6_1;
    io_A_Valid_7_delay_1_5 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_4 <= io_A_Valid_7_delay_1_5;
    io_A_Valid_7_delay_3_3 <= io_A_Valid_7_delay_2_4;
    io_A_Valid_7_delay_4_2 <= io_A_Valid_7_delay_3_3;
    io_A_Valid_7_delay_5_1 <= io_A_Valid_7_delay_4_2;
    io_A_Valid_7_delay_6 <= io_A_Valid_7_delay_5_1;
    io_B_Valid_6_delay_1_6 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_5 <= io_B_Valid_6_delay_1_6;
    io_B_Valid_6_delay_3_4 <= io_B_Valid_6_delay_2_5;
    io_B_Valid_6_delay_4_3 <= io_B_Valid_6_delay_3_4;
    io_B_Valid_6_delay_5_2 <= io_B_Valid_6_delay_4_3;
    io_B_Valid_6_delay_6_1 <= io_B_Valid_6_delay_5_2;
    io_B_Valid_6_delay_7 <= io_B_Valid_6_delay_6_1;
    io_A_Valid_7_delay_1_6 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_5 <= io_A_Valid_7_delay_1_6;
    io_A_Valid_7_delay_3_4 <= io_A_Valid_7_delay_2_5;
    io_A_Valid_7_delay_4_3 <= io_A_Valid_7_delay_3_4;
    io_A_Valid_7_delay_5_2 <= io_A_Valid_7_delay_4_3;
    io_A_Valid_7_delay_6_1 <= io_A_Valid_7_delay_5_2;
    io_A_Valid_7_delay_7 <= io_A_Valid_7_delay_6_1;
    io_B_Valid_7_delay_1_6 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_5 <= io_B_Valid_7_delay_1_6;
    io_B_Valid_7_delay_3_4 <= io_B_Valid_7_delay_2_5;
    io_B_Valid_7_delay_4_3 <= io_B_Valid_7_delay_3_4;
    io_B_Valid_7_delay_5_2 <= io_B_Valid_7_delay_4_3;
    io_B_Valid_7_delay_6_1 <= io_B_Valid_7_delay_5_2;
    io_B_Valid_7_delay_7 <= io_B_Valid_7_delay_6_1;
  end


endmodule

//PE_63 replaced by PE

//PE_62 replaced by PE

//PE_61 replaced by PE

//PE_60 replaced by PE

//PE_59 replaced by PE

//PE_58 replaced by PE

//PE_57 replaced by PE

//PE_56 replaced by PE

//PE_55 replaced by PE

//PE_54 replaced by PE

//PE_53 replaced by PE

//PE_52 replaced by PE

//PE_51 replaced by PE

//PE_50 replaced by PE

//PE_49 replaced by PE

//PE_48 replaced by PE

//PE_47 replaced by PE

//PE_46 replaced by PE

//PE_45 replaced by PE

//PE_44 replaced by PE

//PE_43 replaced by PE

//PE_42 replaced by PE

//PE_41 replaced by PE

//PE_40 replaced by PE

//PE_39 replaced by PE

//PE_38 replaced by PE

//PE_37 replaced by PE

//PE_36 replaced by PE

//PE_35 replaced by PE

//PE_34 replaced by PE

//PE_33 replaced by PE

//PE_32 replaced by PE

//PE_31 replaced by PE

//PE_30 replaced by PE

//PE_29 replaced by PE

//PE_28 replaced by PE

//PE_27 replaced by PE

//PE_26 replaced by PE

//PE_25 replaced by PE

//PE_24 replaced by PE

//PE_23 replaced by PE

//PE_22 replaced by PE

//PE_21 replaced by PE

//PE_20 replaced by PE

//PE_19 replaced by PE

//PE_18 replaced by PE

//PE_17 replaced by PE

//PE_16 replaced by PE

//PE_15 replaced by PE

//PE_14 replaced by PE

//PE_13 replaced by PE

//PE_12 replaced by PE

//PE_11 replaced by PE

//PE_10 replaced by PE

//PE_9 replaced by PE

//PE_8 replaced by PE

//PE_7 replaced by PE

//PE_6 replaced by PE

//PE_5 replaced by PE

//PE_4 replaced by PE

//PE_3 replaced by PE

//PE_2 replaced by PE

//PE_1 replaced by PE

module PE (
  input      [7:0]    activate,
  input      [7:0]    weight,
  input               valid,
  input      [15:0]   signCount,
  output     [7:0]    acount,
  output     [7:0]    bcount,
  output reg [31:0]   PE_OUT,
  output              finish,
  input               clk,
  input               reset
);

  wire       [15:0]   dsp_P;
  wire       [31:0]   _zz_reg1;
  wire       [31:0]   _zz_reg1_1;
  wire       [31:0]   _zz_reg1_2;
  reg        [31:0]   reg1;
  reg                 valid_regNext;
  reg                 valid_regNext_regNext;
  reg        [15:0]   finishCnt_count;
  wire                finishCnt_valid;
  reg                 valid_regNext_1;
  reg        [7:0]    activate_regNext;
  reg        [7:0]    weight_regNext;

  assign _zz_reg1 = {{16{dsp_P[15]}}, dsp_P};
  assign _zz_reg1_1 = 32'h0;
  assign _zz_reg1_2 = {{16{dsp_P[15]}}, dsp_P};
  dsp_marco dsp (
    .CLK (clk          ), //i
    .A   (activate[7:0]), //i
    .B   (weight[7:0]  ), //i
    .P   (dsp_P[15:0]  )  //o
  );
  assign finishCnt_valid = ((finishCnt_count == signCount) && valid_regNext_regNext);
  assign finish = finishCnt_valid;
  always @(*) begin
    PE_OUT = 32'h0;
    if(finishCnt_valid) begin
      PE_OUT = reg1;
    end
  end

  assign acount = activate_regNext;
  assign bcount = weight_regNext;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      reg1 <= 32'h0;
      finishCnt_count <= 16'h0;
    end else begin
      if(valid_regNext_regNext) begin
        if(finishCnt_valid) begin
          finishCnt_count <= 16'h0;
        end else begin
          finishCnt_count <= (finishCnt_count + 16'h0001);
        end
      end
      if(finishCnt_valid) begin
        reg1 <= (valid ? _zz_reg1 : _zz_reg1_1);
      end else begin
        if(valid_regNext_1) begin
          reg1 <= ($signed(_zz_reg1_2) + $signed(reg1));
        end
      end
    end
  end

  always @(posedge clk) begin
    valid_regNext <= valid;
    valid_regNext_regNext <= valid_regNext;
    valid_regNext_1 <= valid;
    activate_regNext <= activate;
    weight_regNext <= weight;
  end


endmodule
