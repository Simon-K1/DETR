// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : SA3D_Top
// Git hash  : 72a3ba00bf8112f87f4c70cf56c4d31a0db88aa8

`timescale 1ns/1ps

module SA3D_Top (
  input               Control_start,
  input               Control_Switch_Conv,
  input      [63:0]   s_axis_s2mm_tdata,
  input      [7:0]    s_axis_s2mm_tkeep,
  input               s_axis_s2mm_tlast,
  output              s_axis_s2mm_tready,
  input               s_axis_s2mm_tvalid,
  input      [4:0]    Img2Col_Stride,
  input      [4:0]    Img2Col_Kernel_Size,
  input      [15:0]   Img2Col_Window_Size,
  input      [15:0]   Img2Col_InFeature_Size,
  input      [15:0]   Img2Col_InFeature_Channel,
  input      [15:0]   Img2Col_OutFeature_Channel,
  input      [15:0]   Img2Col_OutFeature_Size,
  input      [12:0]   Img2Col_Sliding_Size,
  input      [15:0]   Img2Col_OutCol_Count_Times,
  input      [15:0]   Img2Col_InCol_Count_Times,
  input      [15:0]   Img2Col_OutRow_Count_Times,
  input      [15:0]   Img2Col_OutFeature_Channel_Count_Times,
  input      [15:0]   Img2Col_WeightMatrix_Row,
  input      [11:0]   Img2Col_OutMatrix_Col,
  input      [19:0]   Img2Col_OutMatrix_Row,
  input               clk,
  output     [63:0]   m_axis_mm2s_tdata,
  output     [7:0]    m_axis_mm2s_tkeep,
  output              m_axis_mm2s_tlast,
  input               m_axis_mm2s_tready,
  output              m_axis_mm2s_tvalid,
  input               reset
);
  localparam TopCtrl_Enum_IDLE = 6'd1;
  localparam TopCtrl_Enum_INIT = 6'd2;
  localparam TopCtrl_Enum_WEIGHT_CACHE = 6'd4;
  localparam TopCtrl_Enum_RECEIVE_PICTURE = 6'd8;
  localparam TopCtrl_Enum_RECEIVE_MATRIX = 6'd16;
  localparam TopCtrl_Enum_WAIT_COMPUTE_END = 6'd32;

  reg        [1:0]    InputSwitch_Switch;
  reg                 InputSwitch_m_0_axis_mm2s_tready;
  wire                SubModule_Img2Col_start;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_0;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_1;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_2;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_3;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_4;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_5;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_6;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixA_7;
  wire       [7:0]    SubModule_SA_3D__zz_io_MatrixB_0;
  wire                SubModule_SA_3D__zz_io_A_Valid_0;
  wire                SubModule_SA_3D__zz_io_A_Valid_1;
  wire                SubModule_SA_3D__zz_io_A_Valid_2;
  wire                SubModule_SA_3D__zz_io_A_Valid_3;
  wire                SubModule_SA_3D__zz_io_A_Valid_4;
  wire                SubModule_SA_3D__zz_io_A_Valid_5;
  wire                SubModule_SA_3D__zz_io_A_Valid_6;
  wire                SubModule_SA_3D__zz_io_A_Valid_7;
  wire                SubModule_SA_3D__zz_io_B_Valid_0;
  wire       [15:0]   SubModule_SA_3D__zz_io_signCount;
  wire       [7:0]    SubModule_DataArrange_sData_0;
  wire       [7:0]    SubModule_DataArrange_sData_1;
  wire       [7:0]    SubModule_DataArrange_sData_2;
  wire       [7:0]    SubModule_DataArrange_sData_3;
  wire       [7:0]    SubModule_DataArrange_sData_4;
  wire       [7:0]    SubModule_DataArrange_sData_5;
  wire       [7:0]    SubModule_DataArrange_sData_6;
  wire       [7:0]    SubModule_DataArrange_sData_7;
  reg        [7:0]    SubModule_DataArrange_sValid;
  wire       [9:0]    SubModule_DataArrange_OutChannel;
  wire                InputSwitch_s0_axis_s2mm_tready;
  wire       [63:0]   InputSwitch_m_0_axis_mm2s_tdata;
  wire       [7:0]    InputSwitch_m_0_axis_mm2s_tkeep;
  wire                InputSwitch_m_0_axis_mm2s_tlast;
  wire                InputSwitch_m_0_axis_mm2s_tvalid;
  wire       [63:0]   InputSwitch_m_1_axis_mm2s_tdata;
  wire       [7:0]    InputSwitch_m_1_axis_mm2s_tkeep;
  wire                InputSwitch_m_1_axis_mm2s_tlast;
  wire                InputSwitch_m_1_axis_mm2s_tvalid;
  wire       [63:0]   SubModule_Img2Col_mData;
  wire       [7:0]    SubModule_Img2Col_mValid;
  wire                SubModule_Img2Col_s_axis_s2mm_tready;
  wire                SubModule_Img2Col_Raddr_Valid;
  wire                SubModule_Img2Col_LayerEnd;
  wire                SubModule_SA_3D_Matrix_C_valid_0;
  wire                SubModule_SA_3D_Matrix_C_valid_1;
  wire                SubModule_SA_3D_Matrix_C_valid_2;
  wire                SubModule_SA_3D_Matrix_C_valid_3;
  wire                SubModule_SA_3D_Matrix_C_valid_4;
  wire                SubModule_SA_3D_Matrix_C_valid_5;
  wire                SubModule_SA_3D_Matrix_C_valid_6;
  wire                SubModule_SA_3D_Matrix_C_valid_7;
  wire       [31:0]   SubModule_SA_3D_Matrix_C_payload_0;
  wire       [31:0]   SubModule_SA_3D_Matrix_C_payload_1;
  wire       [31:0]   SubModule_SA_3D_Matrix_C_payload_2;
  wire       [31:0]   SubModule_SA_3D_Matrix_C_payload_3;
  wire       [31:0]   SubModule_SA_3D_Matrix_C_payload_4;
  wire       [31:0]   SubModule_SA_3D_Matrix_C_payload_5;
  wire       [31:0]   SubModule_SA_3D_Matrix_C_payload_6;
  wire       [31:0]   SubModule_SA_3D_Matrix_C_payload_7;
  wire                SubModule_WeightCache_s_axis_s2mm_tready;
  wire       [7:0]    SubModule_WeightCache_mData_0;
  wire       [7:0]    SubModule_WeightCache_mData_1;
  wire       [7:0]    SubModule_WeightCache_mData_2;
  wire       [7:0]    SubModule_WeightCache_mData_3;
  wire       [7:0]    SubModule_WeightCache_mData_4;
  wire       [7:0]    SubModule_WeightCache_mData_5;
  wire       [7:0]    SubModule_WeightCache_mData_6;
  wire       [7:0]    SubModule_WeightCache_mData_7;
  wire       [7:0]    SubModule_WeightCache_mData_8;
  wire       [7:0]    SubModule_WeightCache_mData_9;
  wire       [7:0]    SubModule_WeightCache_mData_10;
  wire       [7:0]    SubModule_WeightCache_mData_11;
  wire       [7:0]    SubModule_WeightCache_mData_12;
  wire       [7:0]    SubModule_WeightCache_mData_13;
  wire       [7:0]    SubModule_WeightCache_mData_14;
  wire       [7:0]    SubModule_WeightCache_mData_15;
  wire       [7:0]    SubModule_WeightCache_mData_16;
  wire       [7:0]    SubModule_WeightCache_mData_17;
  wire       [7:0]    SubModule_WeightCache_mData_18;
  wire       [7:0]    SubModule_WeightCache_mData_19;
  wire       [7:0]    SubModule_WeightCache_mData_20;
  wire       [7:0]    SubModule_WeightCache_mData_21;
  wire       [7:0]    SubModule_WeightCache_mData_22;
  wire       [7:0]    SubModule_WeightCache_mData_23;
  wire       [7:0]    SubModule_WeightCache_mData_24;
  wire       [7:0]    SubModule_WeightCache_mData_25;
  wire       [7:0]    SubModule_WeightCache_mData_26;
  wire       [7:0]    SubModule_WeightCache_mData_27;
  wire       [7:0]    SubModule_WeightCache_mData_28;
  wire       [7:0]    SubModule_WeightCache_mData_29;
  wire       [7:0]    SubModule_WeightCache_mData_30;
  wire       [7:0]    SubModule_WeightCache_mData_31;
  wire       [7:0]    SubModule_WeightCache_mData_32;
  wire       [7:0]    SubModule_WeightCache_mData_33;
  wire       [7:0]    SubModule_WeightCache_mData_34;
  wire       [7:0]    SubModule_WeightCache_mData_35;
  wire       [7:0]    SubModule_WeightCache_mData_36;
  wire       [7:0]    SubModule_WeightCache_mData_37;
  wire       [7:0]    SubModule_WeightCache_mData_38;
  wire       [7:0]    SubModule_WeightCache_mData_39;
  wire       [7:0]    SubModule_WeightCache_mData_40;
  wire       [7:0]    SubModule_WeightCache_mData_41;
  wire       [7:0]    SubModule_WeightCache_mData_42;
  wire       [7:0]    SubModule_WeightCache_mData_43;
  wire       [7:0]    SubModule_WeightCache_mData_44;
  wire       [7:0]    SubModule_WeightCache_mData_45;
  wire       [7:0]    SubModule_WeightCache_mData_46;
  wire       [7:0]    SubModule_WeightCache_mData_47;
  wire       [7:0]    SubModule_WeightCache_mData_48;
  wire       [7:0]    SubModule_WeightCache_mData_49;
  wire       [7:0]    SubModule_WeightCache_mData_50;
  wire       [7:0]    SubModule_WeightCache_mData_51;
  wire       [7:0]    SubModule_WeightCache_mData_52;
  wire       [7:0]    SubModule_WeightCache_mData_53;
  wire       [7:0]    SubModule_WeightCache_mData_54;
  wire       [7:0]    SubModule_WeightCache_mData_55;
  wire       [7:0]    SubModule_WeightCache_mData_56;
  wire       [7:0]    SubModule_WeightCache_mData_57;
  wire       [7:0]    SubModule_WeightCache_mData_58;
  wire       [7:0]    SubModule_WeightCache_mData_59;
  wire       [7:0]    SubModule_WeightCache_mData_60;
  wire       [7:0]    SubModule_WeightCache_mData_61;
  wire       [7:0]    SubModule_WeightCache_mData_62;
  wire       [7:0]    SubModule_WeightCache_mData_63;
  wire                SubModule_WeightCache_Weight_Cached;
  wire       [63:0]   SubModule_WeightCache_MatrixCol_Switch;
  wire                SubModule_DataArrange_sReady;
  wire                SubModule_DataArrange_mData_valid;
  wire       [63:0]   SubModule_DataArrange_mData_payload;
  wire                SubModule_DataArrange_mLast;
  wire                SubModule_DataArrange_LayerEnd;
  reg        [5:0]    Fsm_currentState;
  reg        [5:0]    Fsm_nextState;
  wire                Fsm_Inited;
  wire                Fsm_WeightCached;
  wire                Fsm_Picture_Received;
  wire                Fsm_Matrix_Received;
  wire                Fsm_Compute_End;
  wire                Fsm_Switch_Conv;
  wire                when_SA3D_Top_l46;
  wire                when_SA3D_Top_l48;
  wire                LayerEnd;
  wire                when_WaCounter_l19;
  reg        [2:0]    InitCnt_count;
  reg                 InitCnt_valid;
  wire                when_WaCounter_l14;
  wire                when_SA3D_Top_l131;
  reg        [7:0]    _zz_io_MatrixB_1;
  reg                 _zz_io_B_Valid_1;
  reg        [7:0]    _zz_io_MatrixB_2;
  reg        [7:0]    _zz_io_MatrixB_2_1;
  reg                 _zz_io_B_Valid_2;
  reg                 _zz_io_B_Valid_2_1;
  reg        [7:0]    _zz_io_MatrixB_3;
  reg        [7:0]    _zz_io_MatrixB_3_1;
  reg        [7:0]    _zz_io_MatrixB_3_2;
  reg                 _zz_io_B_Valid_3;
  reg                 _zz_io_B_Valid_3_1;
  reg                 _zz_io_B_Valid_3_2;
  reg        [7:0]    _zz_io_MatrixB_4;
  reg        [7:0]    _zz_io_MatrixB_4_1;
  reg        [7:0]    _zz_io_MatrixB_4_2;
  reg        [7:0]    _zz_io_MatrixB_4_3;
  reg                 _zz_io_B_Valid_4;
  reg                 _zz_io_B_Valid_4_1;
  reg                 _zz_io_B_Valid_4_2;
  reg                 _zz_io_B_Valid_4_3;
  reg        [7:0]    _zz_io_MatrixB_5;
  reg        [7:0]    _zz_io_MatrixB_5_1;
  reg        [7:0]    _zz_io_MatrixB_5_2;
  reg        [7:0]    _zz_io_MatrixB_5_3;
  reg        [7:0]    _zz_io_MatrixB_5_4;
  reg                 _zz_io_B_Valid_5;
  reg                 _zz_io_B_Valid_5_1;
  reg                 _zz_io_B_Valid_5_2;
  reg                 _zz_io_B_Valid_5_3;
  reg                 _zz_io_B_Valid_5_4;
  reg        [7:0]    _zz_io_MatrixB_6;
  reg        [7:0]    _zz_io_MatrixB_6_1;
  reg        [7:0]    _zz_io_MatrixB_6_2;
  reg        [7:0]    _zz_io_MatrixB_6_3;
  reg        [7:0]    _zz_io_MatrixB_6_4;
  reg        [7:0]    _zz_io_MatrixB_6_5;
  reg                 _zz_io_B_Valid_6;
  reg                 _zz_io_B_Valid_6_1;
  reg                 _zz_io_B_Valid_6_2;
  reg                 _zz_io_B_Valid_6_3;
  reg                 _zz_io_B_Valid_6_4;
  reg                 _zz_io_B_Valid_6_5;
  reg        [7:0]    _zz_io_MatrixB_7;
  reg        [7:0]    _zz_io_MatrixB_7_1;
  reg        [7:0]    _zz_io_MatrixB_7_2;
  reg        [7:0]    _zz_io_MatrixB_7_3;
  reg        [7:0]    _zz_io_MatrixB_7_4;
  reg        [7:0]    _zz_io_MatrixB_7_5;
  reg        [7:0]    _zz_io_MatrixB_7_6;
  reg                 _zz_io_B_Valid_7;
  reg                 _zz_io_B_Valid_7_1;
  reg                 _zz_io_B_Valid_7_2;
  reg                 _zz_io_B_Valid_7_3;
  reg                 _zz_io_B_Valid_7_4;
  reg                 _zz_io_B_Valid_7_5;
  reg                 _zz_io_B_Valid_7_6;
  reg        [7:0]    _zz_io_MatrixB_8;
  reg        [7:0]    _zz_io_MatrixB_8_1;
  reg        [7:0]    _zz_io_MatrixB_8_2;
  reg        [7:0]    _zz_io_MatrixB_8_3;
  reg        [7:0]    _zz_io_MatrixB_8_4;
  reg        [7:0]    _zz_io_MatrixB_8_5;
  reg        [7:0]    _zz_io_MatrixB_8_6;
  reg        [7:0]    _zz_io_MatrixB_8_7;
  reg                 _zz_io_B_Valid_8;
  reg                 _zz_io_B_Valid_8_1;
  reg                 _zz_io_B_Valid_8_2;
  reg                 _zz_io_B_Valid_8_3;
  reg                 _zz_io_B_Valid_8_4;
  reg                 _zz_io_B_Valid_8_5;
  reg                 _zz_io_B_Valid_8_6;
  reg                 _zz_io_B_Valid_8_7;
  reg        [7:0]    _zz_io_MatrixB_9;
  reg        [7:0]    _zz_io_MatrixB_9_1;
  reg        [7:0]    _zz_io_MatrixB_9_2;
  reg        [7:0]    _zz_io_MatrixB_9_3;
  reg        [7:0]    _zz_io_MatrixB_9_4;
  reg        [7:0]    _zz_io_MatrixB_9_5;
  reg        [7:0]    _zz_io_MatrixB_9_6;
  reg        [7:0]    _zz_io_MatrixB_9_7;
  reg        [7:0]    _zz_io_MatrixB_9_8;
  reg                 _zz_io_B_Valid_9;
  reg                 _zz_io_B_Valid_9_1;
  reg                 _zz_io_B_Valid_9_2;
  reg                 _zz_io_B_Valid_9_3;
  reg                 _zz_io_B_Valid_9_4;
  reg                 _zz_io_B_Valid_9_5;
  reg                 _zz_io_B_Valid_9_6;
  reg                 _zz_io_B_Valid_9_7;
  reg                 _zz_io_B_Valid_9_8;
  reg        [7:0]    _zz_io_MatrixB_10;
  reg        [7:0]    _zz_io_MatrixB_10_1;
  reg        [7:0]    _zz_io_MatrixB_10_2;
  reg        [7:0]    _zz_io_MatrixB_10_3;
  reg        [7:0]    _zz_io_MatrixB_10_4;
  reg        [7:0]    _zz_io_MatrixB_10_5;
  reg        [7:0]    _zz_io_MatrixB_10_6;
  reg        [7:0]    _zz_io_MatrixB_10_7;
  reg        [7:0]    _zz_io_MatrixB_10_8;
  reg        [7:0]    _zz_io_MatrixB_10_9;
  reg                 _zz_io_B_Valid_10;
  reg                 _zz_io_B_Valid_10_1;
  reg                 _zz_io_B_Valid_10_2;
  reg                 _zz_io_B_Valid_10_3;
  reg                 _zz_io_B_Valid_10_4;
  reg                 _zz_io_B_Valid_10_5;
  reg                 _zz_io_B_Valid_10_6;
  reg                 _zz_io_B_Valid_10_7;
  reg                 _zz_io_B_Valid_10_8;
  reg                 _zz_io_B_Valid_10_9;
  reg        [7:0]    _zz_io_MatrixB_11;
  reg        [7:0]    _zz_io_MatrixB_11_1;
  reg        [7:0]    _zz_io_MatrixB_11_2;
  reg        [7:0]    _zz_io_MatrixB_11_3;
  reg        [7:0]    _zz_io_MatrixB_11_4;
  reg        [7:0]    _zz_io_MatrixB_11_5;
  reg        [7:0]    _zz_io_MatrixB_11_6;
  reg        [7:0]    _zz_io_MatrixB_11_7;
  reg        [7:0]    _zz_io_MatrixB_11_8;
  reg        [7:0]    _zz_io_MatrixB_11_9;
  reg        [7:0]    _zz_io_MatrixB_11_10;
  reg                 _zz_io_B_Valid_11;
  reg                 _zz_io_B_Valid_11_1;
  reg                 _zz_io_B_Valid_11_2;
  reg                 _zz_io_B_Valid_11_3;
  reg                 _zz_io_B_Valid_11_4;
  reg                 _zz_io_B_Valid_11_5;
  reg                 _zz_io_B_Valid_11_6;
  reg                 _zz_io_B_Valid_11_7;
  reg                 _zz_io_B_Valid_11_8;
  reg                 _zz_io_B_Valid_11_9;
  reg                 _zz_io_B_Valid_11_10;
  reg        [7:0]    _zz_io_MatrixB_12;
  reg        [7:0]    _zz_io_MatrixB_12_1;
  reg        [7:0]    _zz_io_MatrixB_12_2;
  reg        [7:0]    _zz_io_MatrixB_12_3;
  reg        [7:0]    _zz_io_MatrixB_12_4;
  reg        [7:0]    _zz_io_MatrixB_12_5;
  reg        [7:0]    _zz_io_MatrixB_12_6;
  reg        [7:0]    _zz_io_MatrixB_12_7;
  reg        [7:0]    _zz_io_MatrixB_12_8;
  reg        [7:0]    _zz_io_MatrixB_12_9;
  reg        [7:0]    _zz_io_MatrixB_12_10;
  reg        [7:0]    _zz_io_MatrixB_12_11;
  reg                 _zz_io_B_Valid_12;
  reg                 _zz_io_B_Valid_12_1;
  reg                 _zz_io_B_Valid_12_2;
  reg                 _zz_io_B_Valid_12_3;
  reg                 _zz_io_B_Valid_12_4;
  reg                 _zz_io_B_Valid_12_5;
  reg                 _zz_io_B_Valid_12_6;
  reg                 _zz_io_B_Valid_12_7;
  reg                 _zz_io_B_Valid_12_8;
  reg                 _zz_io_B_Valid_12_9;
  reg                 _zz_io_B_Valid_12_10;
  reg                 _zz_io_B_Valid_12_11;
  reg        [7:0]    _zz_io_MatrixB_13;
  reg        [7:0]    _zz_io_MatrixB_13_1;
  reg        [7:0]    _zz_io_MatrixB_13_2;
  reg        [7:0]    _zz_io_MatrixB_13_3;
  reg        [7:0]    _zz_io_MatrixB_13_4;
  reg        [7:0]    _zz_io_MatrixB_13_5;
  reg        [7:0]    _zz_io_MatrixB_13_6;
  reg        [7:0]    _zz_io_MatrixB_13_7;
  reg        [7:0]    _zz_io_MatrixB_13_8;
  reg        [7:0]    _zz_io_MatrixB_13_9;
  reg        [7:0]    _zz_io_MatrixB_13_10;
  reg        [7:0]    _zz_io_MatrixB_13_11;
  reg        [7:0]    _zz_io_MatrixB_13_12;
  reg                 _zz_io_B_Valid_13;
  reg                 _zz_io_B_Valid_13_1;
  reg                 _zz_io_B_Valid_13_2;
  reg                 _zz_io_B_Valid_13_3;
  reg                 _zz_io_B_Valid_13_4;
  reg                 _zz_io_B_Valid_13_5;
  reg                 _zz_io_B_Valid_13_6;
  reg                 _zz_io_B_Valid_13_7;
  reg                 _zz_io_B_Valid_13_8;
  reg                 _zz_io_B_Valid_13_9;
  reg                 _zz_io_B_Valid_13_10;
  reg                 _zz_io_B_Valid_13_11;
  reg                 _zz_io_B_Valid_13_12;
  reg        [7:0]    _zz_io_MatrixB_14;
  reg        [7:0]    _zz_io_MatrixB_14_1;
  reg        [7:0]    _zz_io_MatrixB_14_2;
  reg        [7:0]    _zz_io_MatrixB_14_3;
  reg        [7:0]    _zz_io_MatrixB_14_4;
  reg        [7:0]    _zz_io_MatrixB_14_5;
  reg        [7:0]    _zz_io_MatrixB_14_6;
  reg        [7:0]    _zz_io_MatrixB_14_7;
  reg        [7:0]    _zz_io_MatrixB_14_8;
  reg        [7:0]    _zz_io_MatrixB_14_9;
  reg        [7:0]    _zz_io_MatrixB_14_10;
  reg        [7:0]    _zz_io_MatrixB_14_11;
  reg        [7:0]    _zz_io_MatrixB_14_12;
  reg        [7:0]    _zz_io_MatrixB_14_13;
  reg                 _zz_io_B_Valid_14;
  reg                 _zz_io_B_Valid_14_1;
  reg                 _zz_io_B_Valid_14_2;
  reg                 _zz_io_B_Valid_14_3;
  reg                 _zz_io_B_Valid_14_4;
  reg                 _zz_io_B_Valid_14_5;
  reg                 _zz_io_B_Valid_14_6;
  reg                 _zz_io_B_Valid_14_7;
  reg                 _zz_io_B_Valid_14_8;
  reg                 _zz_io_B_Valid_14_9;
  reg                 _zz_io_B_Valid_14_10;
  reg                 _zz_io_B_Valid_14_11;
  reg                 _zz_io_B_Valid_14_12;
  reg                 _zz_io_B_Valid_14_13;
  reg        [7:0]    _zz_io_MatrixB_15;
  reg        [7:0]    _zz_io_MatrixB_15_1;
  reg        [7:0]    _zz_io_MatrixB_15_2;
  reg        [7:0]    _zz_io_MatrixB_15_3;
  reg        [7:0]    _zz_io_MatrixB_15_4;
  reg        [7:0]    _zz_io_MatrixB_15_5;
  reg        [7:0]    _zz_io_MatrixB_15_6;
  reg        [7:0]    _zz_io_MatrixB_15_7;
  reg        [7:0]    _zz_io_MatrixB_15_8;
  reg        [7:0]    _zz_io_MatrixB_15_9;
  reg        [7:0]    _zz_io_MatrixB_15_10;
  reg        [7:0]    _zz_io_MatrixB_15_11;
  reg        [7:0]    _zz_io_MatrixB_15_12;
  reg        [7:0]    _zz_io_MatrixB_15_13;
  reg        [7:0]    _zz_io_MatrixB_15_14;
  reg                 _zz_io_B_Valid_15;
  reg                 _zz_io_B_Valid_15_1;
  reg                 _zz_io_B_Valid_15_2;
  reg                 _zz_io_B_Valid_15_3;
  reg                 _zz_io_B_Valid_15_4;
  reg                 _zz_io_B_Valid_15_5;
  reg                 _zz_io_B_Valid_15_6;
  reg                 _zz_io_B_Valid_15_7;
  reg                 _zz_io_B_Valid_15_8;
  reg                 _zz_io_B_Valid_15_9;
  reg                 _zz_io_B_Valid_15_10;
  reg                 _zz_io_B_Valid_15_11;
  reg                 _zz_io_B_Valid_15_12;
  reg                 _zz_io_B_Valid_15_13;
  reg                 _zz_io_B_Valid_15_14;
  reg        [7:0]    _zz_io_MatrixB_16;
  reg        [7:0]    _zz_io_MatrixB_16_1;
  reg        [7:0]    _zz_io_MatrixB_16_2;
  reg        [7:0]    _zz_io_MatrixB_16_3;
  reg        [7:0]    _zz_io_MatrixB_16_4;
  reg        [7:0]    _zz_io_MatrixB_16_5;
  reg        [7:0]    _zz_io_MatrixB_16_6;
  reg        [7:0]    _zz_io_MatrixB_16_7;
  reg        [7:0]    _zz_io_MatrixB_16_8;
  reg        [7:0]    _zz_io_MatrixB_16_9;
  reg        [7:0]    _zz_io_MatrixB_16_10;
  reg        [7:0]    _zz_io_MatrixB_16_11;
  reg        [7:0]    _zz_io_MatrixB_16_12;
  reg        [7:0]    _zz_io_MatrixB_16_13;
  reg        [7:0]    _zz_io_MatrixB_16_14;
  reg        [7:0]    _zz_io_MatrixB_16_15;
  reg                 _zz_io_B_Valid_16;
  reg                 _zz_io_B_Valid_16_1;
  reg                 _zz_io_B_Valid_16_2;
  reg                 _zz_io_B_Valid_16_3;
  reg                 _zz_io_B_Valid_16_4;
  reg                 _zz_io_B_Valid_16_5;
  reg                 _zz_io_B_Valid_16_6;
  reg                 _zz_io_B_Valid_16_7;
  reg                 _zz_io_B_Valid_16_8;
  reg                 _zz_io_B_Valid_16_9;
  reg                 _zz_io_B_Valid_16_10;
  reg                 _zz_io_B_Valid_16_11;
  reg                 _zz_io_B_Valid_16_12;
  reg                 _zz_io_B_Valid_16_13;
  reg                 _zz_io_B_Valid_16_14;
  reg                 _zz_io_B_Valid_16_15;
  reg        [7:0]    _zz_io_MatrixB_17;
  reg        [7:0]    _zz_io_MatrixB_17_1;
  reg        [7:0]    _zz_io_MatrixB_17_2;
  reg        [7:0]    _zz_io_MatrixB_17_3;
  reg        [7:0]    _zz_io_MatrixB_17_4;
  reg        [7:0]    _zz_io_MatrixB_17_5;
  reg        [7:0]    _zz_io_MatrixB_17_6;
  reg        [7:0]    _zz_io_MatrixB_17_7;
  reg        [7:0]    _zz_io_MatrixB_17_8;
  reg        [7:0]    _zz_io_MatrixB_17_9;
  reg        [7:0]    _zz_io_MatrixB_17_10;
  reg        [7:0]    _zz_io_MatrixB_17_11;
  reg        [7:0]    _zz_io_MatrixB_17_12;
  reg        [7:0]    _zz_io_MatrixB_17_13;
  reg        [7:0]    _zz_io_MatrixB_17_14;
  reg        [7:0]    _zz_io_MatrixB_17_15;
  reg        [7:0]    _zz_io_MatrixB_17_16;
  reg                 _zz_io_B_Valid_17;
  reg                 _zz_io_B_Valid_17_1;
  reg                 _zz_io_B_Valid_17_2;
  reg                 _zz_io_B_Valid_17_3;
  reg                 _zz_io_B_Valid_17_4;
  reg                 _zz_io_B_Valid_17_5;
  reg                 _zz_io_B_Valid_17_6;
  reg                 _zz_io_B_Valid_17_7;
  reg                 _zz_io_B_Valid_17_8;
  reg                 _zz_io_B_Valid_17_9;
  reg                 _zz_io_B_Valid_17_10;
  reg                 _zz_io_B_Valid_17_11;
  reg                 _zz_io_B_Valid_17_12;
  reg                 _zz_io_B_Valid_17_13;
  reg                 _zz_io_B_Valid_17_14;
  reg                 _zz_io_B_Valid_17_15;
  reg                 _zz_io_B_Valid_17_16;
  reg        [7:0]    _zz_io_MatrixB_18;
  reg        [7:0]    _zz_io_MatrixB_18_1;
  reg        [7:0]    _zz_io_MatrixB_18_2;
  reg        [7:0]    _zz_io_MatrixB_18_3;
  reg        [7:0]    _zz_io_MatrixB_18_4;
  reg        [7:0]    _zz_io_MatrixB_18_5;
  reg        [7:0]    _zz_io_MatrixB_18_6;
  reg        [7:0]    _zz_io_MatrixB_18_7;
  reg        [7:0]    _zz_io_MatrixB_18_8;
  reg        [7:0]    _zz_io_MatrixB_18_9;
  reg        [7:0]    _zz_io_MatrixB_18_10;
  reg        [7:0]    _zz_io_MatrixB_18_11;
  reg        [7:0]    _zz_io_MatrixB_18_12;
  reg        [7:0]    _zz_io_MatrixB_18_13;
  reg        [7:0]    _zz_io_MatrixB_18_14;
  reg        [7:0]    _zz_io_MatrixB_18_15;
  reg        [7:0]    _zz_io_MatrixB_18_16;
  reg        [7:0]    _zz_io_MatrixB_18_17;
  reg                 _zz_io_B_Valid_18;
  reg                 _zz_io_B_Valid_18_1;
  reg                 _zz_io_B_Valid_18_2;
  reg                 _zz_io_B_Valid_18_3;
  reg                 _zz_io_B_Valid_18_4;
  reg                 _zz_io_B_Valid_18_5;
  reg                 _zz_io_B_Valid_18_6;
  reg                 _zz_io_B_Valid_18_7;
  reg                 _zz_io_B_Valid_18_8;
  reg                 _zz_io_B_Valid_18_9;
  reg                 _zz_io_B_Valid_18_10;
  reg                 _zz_io_B_Valid_18_11;
  reg                 _zz_io_B_Valid_18_12;
  reg                 _zz_io_B_Valid_18_13;
  reg                 _zz_io_B_Valid_18_14;
  reg                 _zz_io_B_Valid_18_15;
  reg                 _zz_io_B_Valid_18_16;
  reg                 _zz_io_B_Valid_18_17;
  reg        [7:0]    _zz_io_MatrixB_19;
  reg        [7:0]    _zz_io_MatrixB_19_1;
  reg        [7:0]    _zz_io_MatrixB_19_2;
  reg        [7:0]    _zz_io_MatrixB_19_3;
  reg        [7:0]    _zz_io_MatrixB_19_4;
  reg        [7:0]    _zz_io_MatrixB_19_5;
  reg        [7:0]    _zz_io_MatrixB_19_6;
  reg        [7:0]    _zz_io_MatrixB_19_7;
  reg        [7:0]    _zz_io_MatrixB_19_8;
  reg        [7:0]    _zz_io_MatrixB_19_9;
  reg        [7:0]    _zz_io_MatrixB_19_10;
  reg        [7:0]    _zz_io_MatrixB_19_11;
  reg        [7:0]    _zz_io_MatrixB_19_12;
  reg        [7:0]    _zz_io_MatrixB_19_13;
  reg        [7:0]    _zz_io_MatrixB_19_14;
  reg        [7:0]    _zz_io_MatrixB_19_15;
  reg        [7:0]    _zz_io_MatrixB_19_16;
  reg        [7:0]    _zz_io_MatrixB_19_17;
  reg        [7:0]    _zz_io_MatrixB_19_18;
  reg                 _zz_io_B_Valid_19;
  reg                 _zz_io_B_Valid_19_1;
  reg                 _zz_io_B_Valid_19_2;
  reg                 _zz_io_B_Valid_19_3;
  reg                 _zz_io_B_Valid_19_4;
  reg                 _zz_io_B_Valid_19_5;
  reg                 _zz_io_B_Valid_19_6;
  reg                 _zz_io_B_Valid_19_7;
  reg                 _zz_io_B_Valid_19_8;
  reg                 _zz_io_B_Valid_19_9;
  reg                 _zz_io_B_Valid_19_10;
  reg                 _zz_io_B_Valid_19_11;
  reg                 _zz_io_B_Valid_19_12;
  reg                 _zz_io_B_Valid_19_13;
  reg                 _zz_io_B_Valid_19_14;
  reg                 _zz_io_B_Valid_19_15;
  reg                 _zz_io_B_Valid_19_16;
  reg                 _zz_io_B_Valid_19_17;
  reg                 _zz_io_B_Valid_19_18;
  reg        [7:0]    _zz_io_MatrixB_20;
  reg        [7:0]    _zz_io_MatrixB_20_1;
  reg        [7:0]    _zz_io_MatrixB_20_2;
  reg        [7:0]    _zz_io_MatrixB_20_3;
  reg        [7:0]    _zz_io_MatrixB_20_4;
  reg        [7:0]    _zz_io_MatrixB_20_5;
  reg        [7:0]    _zz_io_MatrixB_20_6;
  reg        [7:0]    _zz_io_MatrixB_20_7;
  reg        [7:0]    _zz_io_MatrixB_20_8;
  reg        [7:0]    _zz_io_MatrixB_20_9;
  reg        [7:0]    _zz_io_MatrixB_20_10;
  reg        [7:0]    _zz_io_MatrixB_20_11;
  reg        [7:0]    _zz_io_MatrixB_20_12;
  reg        [7:0]    _zz_io_MatrixB_20_13;
  reg        [7:0]    _zz_io_MatrixB_20_14;
  reg        [7:0]    _zz_io_MatrixB_20_15;
  reg        [7:0]    _zz_io_MatrixB_20_16;
  reg        [7:0]    _zz_io_MatrixB_20_17;
  reg        [7:0]    _zz_io_MatrixB_20_18;
  reg        [7:0]    _zz_io_MatrixB_20_19;
  reg                 _zz_io_B_Valid_20;
  reg                 _zz_io_B_Valid_20_1;
  reg                 _zz_io_B_Valid_20_2;
  reg                 _zz_io_B_Valid_20_3;
  reg                 _zz_io_B_Valid_20_4;
  reg                 _zz_io_B_Valid_20_5;
  reg                 _zz_io_B_Valid_20_6;
  reg                 _zz_io_B_Valid_20_7;
  reg                 _zz_io_B_Valid_20_8;
  reg                 _zz_io_B_Valid_20_9;
  reg                 _zz_io_B_Valid_20_10;
  reg                 _zz_io_B_Valid_20_11;
  reg                 _zz_io_B_Valid_20_12;
  reg                 _zz_io_B_Valid_20_13;
  reg                 _zz_io_B_Valid_20_14;
  reg                 _zz_io_B_Valid_20_15;
  reg                 _zz_io_B_Valid_20_16;
  reg                 _zz_io_B_Valid_20_17;
  reg                 _zz_io_B_Valid_20_18;
  reg                 _zz_io_B_Valid_20_19;
  reg        [7:0]    _zz_io_MatrixB_21;
  reg        [7:0]    _zz_io_MatrixB_21_1;
  reg        [7:0]    _zz_io_MatrixB_21_2;
  reg        [7:0]    _zz_io_MatrixB_21_3;
  reg        [7:0]    _zz_io_MatrixB_21_4;
  reg        [7:0]    _zz_io_MatrixB_21_5;
  reg        [7:0]    _zz_io_MatrixB_21_6;
  reg        [7:0]    _zz_io_MatrixB_21_7;
  reg        [7:0]    _zz_io_MatrixB_21_8;
  reg        [7:0]    _zz_io_MatrixB_21_9;
  reg        [7:0]    _zz_io_MatrixB_21_10;
  reg        [7:0]    _zz_io_MatrixB_21_11;
  reg        [7:0]    _zz_io_MatrixB_21_12;
  reg        [7:0]    _zz_io_MatrixB_21_13;
  reg        [7:0]    _zz_io_MatrixB_21_14;
  reg        [7:0]    _zz_io_MatrixB_21_15;
  reg        [7:0]    _zz_io_MatrixB_21_16;
  reg        [7:0]    _zz_io_MatrixB_21_17;
  reg        [7:0]    _zz_io_MatrixB_21_18;
  reg        [7:0]    _zz_io_MatrixB_21_19;
  reg        [7:0]    _zz_io_MatrixB_21_20;
  reg                 _zz_io_B_Valid_21;
  reg                 _zz_io_B_Valid_21_1;
  reg                 _zz_io_B_Valid_21_2;
  reg                 _zz_io_B_Valid_21_3;
  reg                 _zz_io_B_Valid_21_4;
  reg                 _zz_io_B_Valid_21_5;
  reg                 _zz_io_B_Valid_21_6;
  reg                 _zz_io_B_Valid_21_7;
  reg                 _zz_io_B_Valid_21_8;
  reg                 _zz_io_B_Valid_21_9;
  reg                 _zz_io_B_Valid_21_10;
  reg                 _zz_io_B_Valid_21_11;
  reg                 _zz_io_B_Valid_21_12;
  reg                 _zz_io_B_Valid_21_13;
  reg                 _zz_io_B_Valid_21_14;
  reg                 _zz_io_B_Valid_21_15;
  reg                 _zz_io_B_Valid_21_16;
  reg                 _zz_io_B_Valid_21_17;
  reg                 _zz_io_B_Valid_21_18;
  reg                 _zz_io_B_Valid_21_19;
  reg                 _zz_io_B_Valid_21_20;
  reg        [7:0]    _zz_io_MatrixB_22;
  reg        [7:0]    _zz_io_MatrixB_22_1;
  reg        [7:0]    _zz_io_MatrixB_22_2;
  reg        [7:0]    _zz_io_MatrixB_22_3;
  reg        [7:0]    _zz_io_MatrixB_22_4;
  reg        [7:0]    _zz_io_MatrixB_22_5;
  reg        [7:0]    _zz_io_MatrixB_22_6;
  reg        [7:0]    _zz_io_MatrixB_22_7;
  reg        [7:0]    _zz_io_MatrixB_22_8;
  reg        [7:0]    _zz_io_MatrixB_22_9;
  reg        [7:0]    _zz_io_MatrixB_22_10;
  reg        [7:0]    _zz_io_MatrixB_22_11;
  reg        [7:0]    _zz_io_MatrixB_22_12;
  reg        [7:0]    _zz_io_MatrixB_22_13;
  reg        [7:0]    _zz_io_MatrixB_22_14;
  reg        [7:0]    _zz_io_MatrixB_22_15;
  reg        [7:0]    _zz_io_MatrixB_22_16;
  reg        [7:0]    _zz_io_MatrixB_22_17;
  reg        [7:0]    _zz_io_MatrixB_22_18;
  reg        [7:0]    _zz_io_MatrixB_22_19;
  reg        [7:0]    _zz_io_MatrixB_22_20;
  reg        [7:0]    _zz_io_MatrixB_22_21;
  reg                 _zz_io_B_Valid_22;
  reg                 _zz_io_B_Valid_22_1;
  reg                 _zz_io_B_Valid_22_2;
  reg                 _zz_io_B_Valid_22_3;
  reg                 _zz_io_B_Valid_22_4;
  reg                 _zz_io_B_Valid_22_5;
  reg                 _zz_io_B_Valid_22_6;
  reg                 _zz_io_B_Valid_22_7;
  reg                 _zz_io_B_Valid_22_8;
  reg                 _zz_io_B_Valid_22_9;
  reg                 _zz_io_B_Valid_22_10;
  reg                 _zz_io_B_Valid_22_11;
  reg                 _zz_io_B_Valid_22_12;
  reg                 _zz_io_B_Valid_22_13;
  reg                 _zz_io_B_Valid_22_14;
  reg                 _zz_io_B_Valid_22_15;
  reg                 _zz_io_B_Valid_22_16;
  reg                 _zz_io_B_Valid_22_17;
  reg                 _zz_io_B_Valid_22_18;
  reg                 _zz_io_B_Valid_22_19;
  reg                 _zz_io_B_Valid_22_20;
  reg                 _zz_io_B_Valid_22_21;
  reg        [7:0]    _zz_io_MatrixB_23;
  reg        [7:0]    _zz_io_MatrixB_23_1;
  reg        [7:0]    _zz_io_MatrixB_23_2;
  reg        [7:0]    _zz_io_MatrixB_23_3;
  reg        [7:0]    _zz_io_MatrixB_23_4;
  reg        [7:0]    _zz_io_MatrixB_23_5;
  reg        [7:0]    _zz_io_MatrixB_23_6;
  reg        [7:0]    _zz_io_MatrixB_23_7;
  reg        [7:0]    _zz_io_MatrixB_23_8;
  reg        [7:0]    _zz_io_MatrixB_23_9;
  reg        [7:0]    _zz_io_MatrixB_23_10;
  reg        [7:0]    _zz_io_MatrixB_23_11;
  reg        [7:0]    _zz_io_MatrixB_23_12;
  reg        [7:0]    _zz_io_MatrixB_23_13;
  reg        [7:0]    _zz_io_MatrixB_23_14;
  reg        [7:0]    _zz_io_MatrixB_23_15;
  reg        [7:0]    _zz_io_MatrixB_23_16;
  reg        [7:0]    _zz_io_MatrixB_23_17;
  reg        [7:0]    _zz_io_MatrixB_23_18;
  reg        [7:0]    _zz_io_MatrixB_23_19;
  reg        [7:0]    _zz_io_MatrixB_23_20;
  reg        [7:0]    _zz_io_MatrixB_23_21;
  reg        [7:0]    _zz_io_MatrixB_23_22;
  reg                 _zz_io_B_Valid_23;
  reg                 _zz_io_B_Valid_23_1;
  reg                 _zz_io_B_Valid_23_2;
  reg                 _zz_io_B_Valid_23_3;
  reg                 _zz_io_B_Valid_23_4;
  reg                 _zz_io_B_Valid_23_5;
  reg                 _zz_io_B_Valid_23_6;
  reg                 _zz_io_B_Valid_23_7;
  reg                 _zz_io_B_Valid_23_8;
  reg                 _zz_io_B_Valid_23_9;
  reg                 _zz_io_B_Valid_23_10;
  reg                 _zz_io_B_Valid_23_11;
  reg                 _zz_io_B_Valid_23_12;
  reg                 _zz_io_B_Valid_23_13;
  reg                 _zz_io_B_Valid_23_14;
  reg                 _zz_io_B_Valid_23_15;
  reg                 _zz_io_B_Valid_23_16;
  reg                 _zz_io_B_Valid_23_17;
  reg                 _zz_io_B_Valid_23_18;
  reg                 _zz_io_B_Valid_23_19;
  reg                 _zz_io_B_Valid_23_20;
  reg                 _zz_io_B_Valid_23_21;
  reg                 _zz_io_B_Valid_23_22;
  reg        [7:0]    _zz_io_MatrixB_24;
  reg        [7:0]    _zz_io_MatrixB_24_1;
  reg        [7:0]    _zz_io_MatrixB_24_2;
  reg        [7:0]    _zz_io_MatrixB_24_3;
  reg        [7:0]    _zz_io_MatrixB_24_4;
  reg        [7:0]    _zz_io_MatrixB_24_5;
  reg        [7:0]    _zz_io_MatrixB_24_6;
  reg        [7:0]    _zz_io_MatrixB_24_7;
  reg        [7:0]    _zz_io_MatrixB_24_8;
  reg        [7:0]    _zz_io_MatrixB_24_9;
  reg        [7:0]    _zz_io_MatrixB_24_10;
  reg        [7:0]    _zz_io_MatrixB_24_11;
  reg        [7:0]    _zz_io_MatrixB_24_12;
  reg        [7:0]    _zz_io_MatrixB_24_13;
  reg        [7:0]    _zz_io_MatrixB_24_14;
  reg        [7:0]    _zz_io_MatrixB_24_15;
  reg        [7:0]    _zz_io_MatrixB_24_16;
  reg        [7:0]    _zz_io_MatrixB_24_17;
  reg        [7:0]    _zz_io_MatrixB_24_18;
  reg        [7:0]    _zz_io_MatrixB_24_19;
  reg        [7:0]    _zz_io_MatrixB_24_20;
  reg        [7:0]    _zz_io_MatrixB_24_21;
  reg        [7:0]    _zz_io_MatrixB_24_22;
  reg        [7:0]    _zz_io_MatrixB_24_23;
  reg                 _zz_io_B_Valid_24;
  reg                 _zz_io_B_Valid_24_1;
  reg                 _zz_io_B_Valid_24_2;
  reg                 _zz_io_B_Valid_24_3;
  reg                 _zz_io_B_Valid_24_4;
  reg                 _zz_io_B_Valid_24_5;
  reg                 _zz_io_B_Valid_24_6;
  reg                 _zz_io_B_Valid_24_7;
  reg                 _zz_io_B_Valid_24_8;
  reg                 _zz_io_B_Valid_24_9;
  reg                 _zz_io_B_Valid_24_10;
  reg                 _zz_io_B_Valid_24_11;
  reg                 _zz_io_B_Valid_24_12;
  reg                 _zz_io_B_Valid_24_13;
  reg                 _zz_io_B_Valid_24_14;
  reg                 _zz_io_B_Valid_24_15;
  reg                 _zz_io_B_Valid_24_16;
  reg                 _zz_io_B_Valid_24_17;
  reg                 _zz_io_B_Valid_24_18;
  reg                 _zz_io_B_Valid_24_19;
  reg                 _zz_io_B_Valid_24_20;
  reg                 _zz_io_B_Valid_24_21;
  reg                 _zz_io_B_Valid_24_22;
  reg                 _zz_io_B_Valid_24_23;
  reg        [7:0]    _zz_io_MatrixB_25;
  reg        [7:0]    _zz_io_MatrixB_25_1;
  reg        [7:0]    _zz_io_MatrixB_25_2;
  reg        [7:0]    _zz_io_MatrixB_25_3;
  reg        [7:0]    _zz_io_MatrixB_25_4;
  reg        [7:0]    _zz_io_MatrixB_25_5;
  reg        [7:0]    _zz_io_MatrixB_25_6;
  reg        [7:0]    _zz_io_MatrixB_25_7;
  reg        [7:0]    _zz_io_MatrixB_25_8;
  reg        [7:0]    _zz_io_MatrixB_25_9;
  reg        [7:0]    _zz_io_MatrixB_25_10;
  reg        [7:0]    _zz_io_MatrixB_25_11;
  reg        [7:0]    _zz_io_MatrixB_25_12;
  reg        [7:0]    _zz_io_MatrixB_25_13;
  reg        [7:0]    _zz_io_MatrixB_25_14;
  reg        [7:0]    _zz_io_MatrixB_25_15;
  reg        [7:0]    _zz_io_MatrixB_25_16;
  reg        [7:0]    _zz_io_MatrixB_25_17;
  reg        [7:0]    _zz_io_MatrixB_25_18;
  reg        [7:0]    _zz_io_MatrixB_25_19;
  reg        [7:0]    _zz_io_MatrixB_25_20;
  reg        [7:0]    _zz_io_MatrixB_25_21;
  reg        [7:0]    _zz_io_MatrixB_25_22;
  reg        [7:0]    _zz_io_MatrixB_25_23;
  reg        [7:0]    _zz_io_MatrixB_25_24;
  reg                 _zz_io_B_Valid_25;
  reg                 _zz_io_B_Valid_25_1;
  reg                 _zz_io_B_Valid_25_2;
  reg                 _zz_io_B_Valid_25_3;
  reg                 _zz_io_B_Valid_25_4;
  reg                 _zz_io_B_Valid_25_5;
  reg                 _zz_io_B_Valid_25_6;
  reg                 _zz_io_B_Valid_25_7;
  reg                 _zz_io_B_Valid_25_8;
  reg                 _zz_io_B_Valid_25_9;
  reg                 _zz_io_B_Valid_25_10;
  reg                 _zz_io_B_Valid_25_11;
  reg                 _zz_io_B_Valid_25_12;
  reg                 _zz_io_B_Valid_25_13;
  reg                 _zz_io_B_Valid_25_14;
  reg                 _zz_io_B_Valid_25_15;
  reg                 _zz_io_B_Valid_25_16;
  reg                 _zz_io_B_Valid_25_17;
  reg                 _zz_io_B_Valid_25_18;
  reg                 _zz_io_B_Valid_25_19;
  reg                 _zz_io_B_Valid_25_20;
  reg                 _zz_io_B_Valid_25_21;
  reg                 _zz_io_B_Valid_25_22;
  reg                 _zz_io_B_Valid_25_23;
  reg                 _zz_io_B_Valid_25_24;
  reg        [7:0]    _zz_io_MatrixB_26;
  reg        [7:0]    _zz_io_MatrixB_26_1;
  reg        [7:0]    _zz_io_MatrixB_26_2;
  reg        [7:0]    _zz_io_MatrixB_26_3;
  reg        [7:0]    _zz_io_MatrixB_26_4;
  reg        [7:0]    _zz_io_MatrixB_26_5;
  reg        [7:0]    _zz_io_MatrixB_26_6;
  reg        [7:0]    _zz_io_MatrixB_26_7;
  reg        [7:0]    _zz_io_MatrixB_26_8;
  reg        [7:0]    _zz_io_MatrixB_26_9;
  reg        [7:0]    _zz_io_MatrixB_26_10;
  reg        [7:0]    _zz_io_MatrixB_26_11;
  reg        [7:0]    _zz_io_MatrixB_26_12;
  reg        [7:0]    _zz_io_MatrixB_26_13;
  reg        [7:0]    _zz_io_MatrixB_26_14;
  reg        [7:0]    _zz_io_MatrixB_26_15;
  reg        [7:0]    _zz_io_MatrixB_26_16;
  reg        [7:0]    _zz_io_MatrixB_26_17;
  reg        [7:0]    _zz_io_MatrixB_26_18;
  reg        [7:0]    _zz_io_MatrixB_26_19;
  reg        [7:0]    _zz_io_MatrixB_26_20;
  reg        [7:0]    _zz_io_MatrixB_26_21;
  reg        [7:0]    _zz_io_MatrixB_26_22;
  reg        [7:0]    _zz_io_MatrixB_26_23;
  reg        [7:0]    _zz_io_MatrixB_26_24;
  reg        [7:0]    _zz_io_MatrixB_26_25;
  reg                 _zz_io_B_Valid_26;
  reg                 _zz_io_B_Valid_26_1;
  reg                 _zz_io_B_Valid_26_2;
  reg                 _zz_io_B_Valid_26_3;
  reg                 _zz_io_B_Valid_26_4;
  reg                 _zz_io_B_Valid_26_5;
  reg                 _zz_io_B_Valid_26_6;
  reg                 _zz_io_B_Valid_26_7;
  reg                 _zz_io_B_Valid_26_8;
  reg                 _zz_io_B_Valid_26_9;
  reg                 _zz_io_B_Valid_26_10;
  reg                 _zz_io_B_Valid_26_11;
  reg                 _zz_io_B_Valid_26_12;
  reg                 _zz_io_B_Valid_26_13;
  reg                 _zz_io_B_Valid_26_14;
  reg                 _zz_io_B_Valid_26_15;
  reg                 _zz_io_B_Valid_26_16;
  reg                 _zz_io_B_Valid_26_17;
  reg                 _zz_io_B_Valid_26_18;
  reg                 _zz_io_B_Valid_26_19;
  reg                 _zz_io_B_Valid_26_20;
  reg                 _zz_io_B_Valid_26_21;
  reg                 _zz_io_B_Valid_26_22;
  reg                 _zz_io_B_Valid_26_23;
  reg                 _zz_io_B_Valid_26_24;
  reg                 _zz_io_B_Valid_26_25;
  reg        [7:0]    _zz_io_MatrixB_27;
  reg        [7:0]    _zz_io_MatrixB_27_1;
  reg        [7:0]    _zz_io_MatrixB_27_2;
  reg        [7:0]    _zz_io_MatrixB_27_3;
  reg        [7:0]    _zz_io_MatrixB_27_4;
  reg        [7:0]    _zz_io_MatrixB_27_5;
  reg        [7:0]    _zz_io_MatrixB_27_6;
  reg        [7:0]    _zz_io_MatrixB_27_7;
  reg        [7:0]    _zz_io_MatrixB_27_8;
  reg        [7:0]    _zz_io_MatrixB_27_9;
  reg        [7:0]    _zz_io_MatrixB_27_10;
  reg        [7:0]    _zz_io_MatrixB_27_11;
  reg        [7:0]    _zz_io_MatrixB_27_12;
  reg        [7:0]    _zz_io_MatrixB_27_13;
  reg        [7:0]    _zz_io_MatrixB_27_14;
  reg        [7:0]    _zz_io_MatrixB_27_15;
  reg        [7:0]    _zz_io_MatrixB_27_16;
  reg        [7:0]    _zz_io_MatrixB_27_17;
  reg        [7:0]    _zz_io_MatrixB_27_18;
  reg        [7:0]    _zz_io_MatrixB_27_19;
  reg        [7:0]    _zz_io_MatrixB_27_20;
  reg        [7:0]    _zz_io_MatrixB_27_21;
  reg        [7:0]    _zz_io_MatrixB_27_22;
  reg        [7:0]    _zz_io_MatrixB_27_23;
  reg        [7:0]    _zz_io_MatrixB_27_24;
  reg        [7:0]    _zz_io_MatrixB_27_25;
  reg        [7:0]    _zz_io_MatrixB_27_26;
  reg                 _zz_io_B_Valid_27;
  reg                 _zz_io_B_Valid_27_1;
  reg                 _zz_io_B_Valid_27_2;
  reg                 _zz_io_B_Valid_27_3;
  reg                 _zz_io_B_Valid_27_4;
  reg                 _zz_io_B_Valid_27_5;
  reg                 _zz_io_B_Valid_27_6;
  reg                 _zz_io_B_Valid_27_7;
  reg                 _zz_io_B_Valid_27_8;
  reg                 _zz_io_B_Valid_27_9;
  reg                 _zz_io_B_Valid_27_10;
  reg                 _zz_io_B_Valid_27_11;
  reg                 _zz_io_B_Valid_27_12;
  reg                 _zz_io_B_Valid_27_13;
  reg                 _zz_io_B_Valid_27_14;
  reg                 _zz_io_B_Valid_27_15;
  reg                 _zz_io_B_Valid_27_16;
  reg                 _zz_io_B_Valid_27_17;
  reg                 _zz_io_B_Valid_27_18;
  reg                 _zz_io_B_Valid_27_19;
  reg                 _zz_io_B_Valid_27_20;
  reg                 _zz_io_B_Valid_27_21;
  reg                 _zz_io_B_Valid_27_22;
  reg                 _zz_io_B_Valid_27_23;
  reg                 _zz_io_B_Valid_27_24;
  reg                 _zz_io_B_Valid_27_25;
  reg                 _zz_io_B_Valid_27_26;
  reg        [7:0]    _zz_io_MatrixB_28;
  reg        [7:0]    _zz_io_MatrixB_28_1;
  reg        [7:0]    _zz_io_MatrixB_28_2;
  reg        [7:0]    _zz_io_MatrixB_28_3;
  reg        [7:0]    _zz_io_MatrixB_28_4;
  reg        [7:0]    _zz_io_MatrixB_28_5;
  reg        [7:0]    _zz_io_MatrixB_28_6;
  reg        [7:0]    _zz_io_MatrixB_28_7;
  reg        [7:0]    _zz_io_MatrixB_28_8;
  reg        [7:0]    _zz_io_MatrixB_28_9;
  reg        [7:0]    _zz_io_MatrixB_28_10;
  reg        [7:0]    _zz_io_MatrixB_28_11;
  reg        [7:0]    _zz_io_MatrixB_28_12;
  reg        [7:0]    _zz_io_MatrixB_28_13;
  reg        [7:0]    _zz_io_MatrixB_28_14;
  reg        [7:0]    _zz_io_MatrixB_28_15;
  reg        [7:0]    _zz_io_MatrixB_28_16;
  reg        [7:0]    _zz_io_MatrixB_28_17;
  reg        [7:0]    _zz_io_MatrixB_28_18;
  reg        [7:0]    _zz_io_MatrixB_28_19;
  reg        [7:0]    _zz_io_MatrixB_28_20;
  reg        [7:0]    _zz_io_MatrixB_28_21;
  reg        [7:0]    _zz_io_MatrixB_28_22;
  reg        [7:0]    _zz_io_MatrixB_28_23;
  reg        [7:0]    _zz_io_MatrixB_28_24;
  reg        [7:0]    _zz_io_MatrixB_28_25;
  reg        [7:0]    _zz_io_MatrixB_28_26;
  reg        [7:0]    _zz_io_MatrixB_28_27;
  reg                 _zz_io_B_Valid_28;
  reg                 _zz_io_B_Valid_28_1;
  reg                 _zz_io_B_Valid_28_2;
  reg                 _zz_io_B_Valid_28_3;
  reg                 _zz_io_B_Valid_28_4;
  reg                 _zz_io_B_Valid_28_5;
  reg                 _zz_io_B_Valid_28_6;
  reg                 _zz_io_B_Valid_28_7;
  reg                 _zz_io_B_Valid_28_8;
  reg                 _zz_io_B_Valid_28_9;
  reg                 _zz_io_B_Valid_28_10;
  reg                 _zz_io_B_Valid_28_11;
  reg                 _zz_io_B_Valid_28_12;
  reg                 _zz_io_B_Valid_28_13;
  reg                 _zz_io_B_Valid_28_14;
  reg                 _zz_io_B_Valid_28_15;
  reg                 _zz_io_B_Valid_28_16;
  reg                 _zz_io_B_Valid_28_17;
  reg                 _zz_io_B_Valid_28_18;
  reg                 _zz_io_B_Valid_28_19;
  reg                 _zz_io_B_Valid_28_20;
  reg                 _zz_io_B_Valid_28_21;
  reg                 _zz_io_B_Valid_28_22;
  reg                 _zz_io_B_Valid_28_23;
  reg                 _zz_io_B_Valid_28_24;
  reg                 _zz_io_B_Valid_28_25;
  reg                 _zz_io_B_Valid_28_26;
  reg                 _zz_io_B_Valid_28_27;
  reg        [7:0]    _zz_io_MatrixB_29;
  reg        [7:0]    _zz_io_MatrixB_29_1;
  reg        [7:0]    _zz_io_MatrixB_29_2;
  reg        [7:0]    _zz_io_MatrixB_29_3;
  reg        [7:0]    _zz_io_MatrixB_29_4;
  reg        [7:0]    _zz_io_MatrixB_29_5;
  reg        [7:0]    _zz_io_MatrixB_29_6;
  reg        [7:0]    _zz_io_MatrixB_29_7;
  reg        [7:0]    _zz_io_MatrixB_29_8;
  reg        [7:0]    _zz_io_MatrixB_29_9;
  reg        [7:0]    _zz_io_MatrixB_29_10;
  reg        [7:0]    _zz_io_MatrixB_29_11;
  reg        [7:0]    _zz_io_MatrixB_29_12;
  reg        [7:0]    _zz_io_MatrixB_29_13;
  reg        [7:0]    _zz_io_MatrixB_29_14;
  reg        [7:0]    _zz_io_MatrixB_29_15;
  reg        [7:0]    _zz_io_MatrixB_29_16;
  reg        [7:0]    _zz_io_MatrixB_29_17;
  reg        [7:0]    _zz_io_MatrixB_29_18;
  reg        [7:0]    _zz_io_MatrixB_29_19;
  reg        [7:0]    _zz_io_MatrixB_29_20;
  reg        [7:0]    _zz_io_MatrixB_29_21;
  reg        [7:0]    _zz_io_MatrixB_29_22;
  reg        [7:0]    _zz_io_MatrixB_29_23;
  reg        [7:0]    _zz_io_MatrixB_29_24;
  reg        [7:0]    _zz_io_MatrixB_29_25;
  reg        [7:0]    _zz_io_MatrixB_29_26;
  reg        [7:0]    _zz_io_MatrixB_29_27;
  reg        [7:0]    _zz_io_MatrixB_29_28;
  reg                 _zz_io_B_Valid_29;
  reg                 _zz_io_B_Valid_29_1;
  reg                 _zz_io_B_Valid_29_2;
  reg                 _zz_io_B_Valid_29_3;
  reg                 _zz_io_B_Valid_29_4;
  reg                 _zz_io_B_Valid_29_5;
  reg                 _zz_io_B_Valid_29_6;
  reg                 _zz_io_B_Valid_29_7;
  reg                 _zz_io_B_Valid_29_8;
  reg                 _zz_io_B_Valid_29_9;
  reg                 _zz_io_B_Valid_29_10;
  reg                 _zz_io_B_Valid_29_11;
  reg                 _zz_io_B_Valid_29_12;
  reg                 _zz_io_B_Valid_29_13;
  reg                 _zz_io_B_Valid_29_14;
  reg                 _zz_io_B_Valid_29_15;
  reg                 _zz_io_B_Valid_29_16;
  reg                 _zz_io_B_Valid_29_17;
  reg                 _zz_io_B_Valid_29_18;
  reg                 _zz_io_B_Valid_29_19;
  reg                 _zz_io_B_Valid_29_20;
  reg                 _zz_io_B_Valid_29_21;
  reg                 _zz_io_B_Valid_29_22;
  reg                 _zz_io_B_Valid_29_23;
  reg                 _zz_io_B_Valid_29_24;
  reg                 _zz_io_B_Valid_29_25;
  reg                 _zz_io_B_Valid_29_26;
  reg                 _zz_io_B_Valid_29_27;
  reg                 _zz_io_B_Valid_29_28;
  reg        [7:0]    _zz_io_MatrixB_30;
  reg        [7:0]    _zz_io_MatrixB_30_1;
  reg        [7:0]    _zz_io_MatrixB_30_2;
  reg        [7:0]    _zz_io_MatrixB_30_3;
  reg        [7:0]    _zz_io_MatrixB_30_4;
  reg        [7:0]    _zz_io_MatrixB_30_5;
  reg        [7:0]    _zz_io_MatrixB_30_6;
  reg        [7:0]    _zz_io_MatrixB_30_7;
  reg        [7:0]    _zz_io_MatrixB_30_8;
  reg        [7:0]    _zz_io_MatrixB_30_9;
  reg        [7:0]    _zz_io_MatrixB_30_10;
  reg        [7:0]    _zz_io_MatrixB_30_11;
  reg        [7:0]    _zz_io_MatrixB_30_12;
  reg        [7:0]    _zz_io_MatrixB_30_13;
  reg        [7:0]    _zz_io_MatrixB_30_14;
  reg        [7:0]    _zz_io_MatrixB_30_15;
  reg        [7:0]    _zz_io_MatrixB_30_16;
  reg        [7:0]    _zz_io_MatrixB_30_17;
  reg        [7:0]    _zz_io_MatrixB_30_18;
  reg        [7:0]    _zz_io_MatrixB_30_19;
  reg        [7:0]    _zz_io_MatrixB_30_20;
  reg        [7:0]    _zz_io_MatrixB_30_21;
  reg        [7:0]    _zz_io_MatrixB_30_22;
  reg        [7:0]    _zz_io_MatrixB_30_23;
  reg        [7:0]    _zz_io_MatrixB_30_24;
  reg        [7:0]    _zz_io_MatrixB_30_25;
  reg        [7:0]    _zz_io_MatrixB_30_26;
  reg        [7:0]    _zz_io_MatrixB_30_27;
  reg        [7:0]    _zz_io_MatrixB_30_28;
  reg        [7:0]    _zz_io_MatrixB_30_29;
  reg                 _zz_io_B_Valid_30;
  reg                 _zz_io_B_Valid_30_1;
  reg                 _zz_io_B_Valid_30_2;
  reg                 _zz_io_B_Valid_30_3;
  reg                 _zz_io_B_Valid_30_4;
  reg                 _zz_io_B_Valid_30_5;
  reg                 _zz_io_B_Valid_30_6;
  reg                 _zz_io_B_Valid_30_7;
  reg                 _zz_io_B_Valid_30_8;
  reg                 _zz_io_B_Valid_30_9;
  reg                 _zz_io_B_Valid_30_10;
  reg                 _zz_io_B_Valid_30_11;
  reg                 _zz_io_B_Valid_30_12;
  reg                 _zz_io_B_Valid_30_13;
  reg                 _zz_io_B_Valid_30_14;
  reg                 _zz_io_B_Valid_30_15;
  reg                 _zz_io_B_Valid_30_16;
  reg                 _zz_io_B_Valid_30_17;
  reg                 _zz_io_B_Valid_30_18;
  reg                 _zz_io_B_Valid_30_19;
  reg                 _zz_io_B_Valid_30_20;
  reg                 _zz_io_B_Valid_30_21;
  reg                 _zz_io_B_Valid_30_22;
  reg                 _zz_io_B_Valid_30_23;
  reg                 _zz_io_B_Valid_30_24;
  reg                 _zz_io_B_Valid_30_25;
  reg                 _zz_io_B_Valid_30_26;
  reg                 _zz_io_B_Valid_30_27;
  reg                 _zz_io_B_Valid_30_28;
  reg                 _zz_io_B_Valid_30_29;
  reg        [7:0]    _zz_io_MatrixB_31;
  reg        [7:0]    _zz_io_MatrixB_31_1;
  reg        [7:0]    _zz_io_MatrixB_31_2;
  reg        [7:0]    _zz_io_MatrixB_31_3;
  reg        [7:0]    _zz_io_MatrixB_31_4;
  reg        [7:0]    _zz_io_MatrixB_31_5;
  reg        [7:0]    _zz_io_MatrixB_31_6;
  reg        [7:0]    _zz_io_MatrixB_31_7;
  reg        [7:0]    _zz_io_MatrixB_31_8;
  reg        [7:0]    _zz_io_MatrixB_31_9;
  reg        [7:0]    _zz_io_MatrixB_31_10;
  reg        [7:0]    _zz_io_MatrixB_31_11;
  reg        [7:0]    _zz_io_MatrixB_31_12;
  reg        [7:0]    _zz_io_MatrixB_31_13;
  reg        [7:0]    _zz_io_MatrixB_31_14;
  reg        [7:0]    _zz_io_MatrixB_31_15;
  reg        [7:0]    _zz_io_MatrixB_31_16;
  reg        [7:0]    _zz_io_MatrixB_31_17;
  reg        [7:0]    _zz_io_MatrixB_31_18;
  reg        [7:0]    _zz_io_MatrixB_31_19;
  reg        [7:0]    _zz_io_MatrixB_31_20;
  reg        [7:0]    _zz_io_MatrixB_31_21;
  reg        [7:0]    _zz_io_MatrixB_31_22;
  reg        [7:0]    _zz_io_MatrixB_31_23;
  reg        [7:0]    _zz_io_MatrixB_31_24;
  reg        [7:0]    _zz_io_MatrixB_31_25;
  reg        [7:0]    _zz_io_MatrixB_31_26;
  reg        [7:0]    _zz_io_MatrixB_31_27;
  reg        [7:0]    _zz_io_MatrixB_31_28;
  reg        [7:0]    _zz_io_MatrixB_31_29;
  reg        [7:0]    _zz_io_MatrixB_31_30;
  reg                 _zz_io_B_Valid_31;
  reg                 _zz_io_B_Valid_31_1;
  reg                 _zz_io_B_Valid_31_2;
  reg                 _zz_io_B_Valid_31_3;
  reg                 _zz_io_B_Valid_31_4;
  reg                 _zz_io_B_Valid_31_5;
  reg                 _zz_io_B_Valid_31_6;
  reg                 _zz_io_B_Valid_31_7;
  reg                 _zz_io_B_Valid_31_8;
  reg                 _zz_io_B_Valid_31_9;
  reg                 _zz_io_B_Valid_31_10;
  reg                 _zz_io_B_Valid_31_11;
  reg                 _zz_io_B_Valid_31_12;
  reg                 _zz_io_B_Valid_31_13;
  reg                 _zz_io_B_Valid_31_14;
  reg                 _zz_io_B_Valid_31_15;
  reg                 _zz_io_B_Valid_31_16;
  reg                 _zz_io_B_Valid_31_17;
  reg                 _zz_io_B_Valid_31_18;
  reg                 _zz_io_B_Valid_31_19;
  reg                 _zz_io_B_Valid_31_20;
  reg                 _zz_io_B_Valid_31_21;
  reg                 _zz_io_B_Valid_31_22;
  reg                 _zz_io_B_Valid_31_23;
  reg                 _zz_io_B_Valid_31_24;
  reg                 _zz_io_B_Valid_31_25;
  reg                 _zz_io_B_Valid_31_26;
  reg                 _zz_io_B_Valid_31_27;
  reg                 _zz_io_B_Valid_31_28;
  reg                 _zz_io_B_Valid_31_29;
  reg                 _zz_io_B_Valid_31_30;
  reg        [7:0]    _zz_io_MatrixB_32;
  reg        [7:0]    _zz_io_MatrixB_32_1;
  reg        [7:0]    _zz_io_MatrixB_32_2;
  reg        [7:0]    _zz_io_MatrixB_32_3;
  reg        [7:0]    _zz_io_MatrixB_32_4;
  reg        [7:0]    _zz_io_MatrixB_32_5;
  reg        [7:0]    _zz_io_MatrixB_32_6;
  reg        [7:0]    _zz_io_MatrixB_32_7;
  reg        [7:0]    _zz_io_MatrixB_32_8;
  reg        [7:0]    _zz_io_MatrixB_32_9;
  reg        [7:0]    _zz_io_MatrixB_32_10;
  reg        [7:0]    _zz_io_MatrixB_32_11;
  reg        [7:0]    _zz_io_MatrixB_32_12;
  reg        [7:0]    _zz_io_MatrixB_32_13;
  reg        [7:0]    _zz_io_MatrixB_32_14;
  reg        [7:0]    _zz_io_MatrixB_32_15;
  reg        [7:0]    _zz_io_MatrixB_32_16;
  reg        [7:0]    _zz_io_MatrixB_32_17;
  reg        [7:0]    _zz_io_MatrixB_32_18;
  reg        [7:0]    _zz_io_MatrixB_32_19;
  reg        [7:0]    _zz_io_MatrixB_32_20;
  reg        [7:0]    _zz_io_MatrixB_32_21;
  reg        [7:0]    _zz_io_MatrixB_32_22;
  reg        [7:0]    _zz_io_MatrixB_32_23;
  reg        [7:0]    _zz_io_MatrixB_32_24;
  reg        [7:0]    _zz_io_MatrixB_32_25;
  reg        [7:0]    _zz_io_MatrixB_32_26;
  reg        [7:0]    _zz_io_MatrixB_32_27;
  reg        [7:0]    _zz_io_MatrixB_32_28;
  reg        [7:0]    _zz_io_MatrixB_32_29;
  reg        [7:0]    _zz_io_MatrixB_32_30;
  reg        [7:0]    _zz_io_MatrixB_32_31;
  reg                 _zz_io_B_Valid_32;
  reg                 _zz_io_B_Valid_32_1;
  reg                 _zz_io_B_Valid_32_2;
  reg                 _zz_io_B_Valid_32_3;
  reg                 _zz_io_B_Valid_32_4;
  reg                 _zz_io_B_Valid_32_5;
  reg                 _zz_io_B_Valid_32_6;
  reg                 _zz_io_B_Valid_32_7;
  reg                 _zz_io_B_Valid_32_8;
  reg                 _zz_io_B_Valid_32_9;
  reg                 _zz_io_B_Valid_32_10;
  reg                 _zz_io_B_Valid_32_11;
  reg                 _zz_io_B_Valid_32_12;
  reg                 _zz_io_B_Valid_32_13;
  reg                 _zz_io_B_Valid_32_14;
  reg                 _zz_io_B_Valid_32_15;
  reg                 _zz_io_B_Valid_32_16;
  reg                 _zz_io_B_Valid_32_17;
  reg                 _zz_io_B_Valid_32_18;
  reg                 _zz_io_B_Valid_32_19;
  reg                 _zz_io_B_Valid_32_20;
  reg                 _zz_io_B_Valid_32_21;
  reg                 _zz_io_B_Valid_32_22;
  reg                 _zz_io_B_Valid_32_23;
  reg                 _zz_io_B_Valid_32_24;
  reg                 _zz_io_B_Valid_32_25;
  reg                 _zz_io_B_Valid_32_26;
  reg                 _zz_io_B_Valid_32_27;
  reg                 _zz_io_B_Valid_32_28;
  reg                 _zz_io_B_Valid_32_29;
  reg                 _zz_io_B_Valid_32_30;
  reg                 _zz_io_B_Valid_32_31;
  reg        [7:0]    _zz_io_MatrixB_33;
  reg        [7:0]    _zz_io_MatrixB_33_1;
  reg        [7:0]    _zz_io_MatrixB_33_2;
  reg        [7:0]    _zz_io_MatrixB_33_3;
  reg        [7:0]    _zz_io_MatrixB_33_4;
  reg        [7:0]    _zz_io_MatrixB_33_5;
  reg        [7:0]    _zz_io_MatrixB_33_6;
  reg        [7:0]    _zz_io_MatrixB_33_7;
  reg        [7:0]    _zz_io_MatrixB_33_8;
  reg        [7:0]    _zz_io_MatrixB_33_9;
  reg        [7:0]    _zz_io_MatrixB_33_10;
  reg        [7:0]    _zz_io_MatrixB_33_11;
  reg        [7:0]    _zz_io_MatrixB_33_12;
  reg        [7:0]    _zz_io_MatrixB_33_13;
  reg        [7:0]    _zz_io_MatrixB_33_14;
  reg        [7:0]    _zz_io_MatrixB_33_15;
  reg        [7:0]    _zz_io_MatrixB_33_16;
  reg        [7:0]    _zz_io_MatrixB_33_17;
  reg        [7:0]    _zz_io_MatrixB_33_18;
  reg        [7:0]    _zz_io_MatrixB_33_19;
  reg        [7:0]    _zz_io_MatrixB_33_20;
  reg        [7:0]    _zz_io_MatrixB_33_21;
  reg        [7:0]    _zz_io_MatrixB_33_22;
  reg        [7:0]    _zz_io_MatrixB_33_23;
  reg        [7:0]    _zz_io_MatrixB_33_24;
  reg        [7:0]    _zz_io_MatrixB_33_25;
  reg        [7:0]    _zz_io_MatrixB_33_26;
  reg        [7:0]    _zz_io_MatrixB_33_27;
  reg        [7:0]    _zz_io_MatrixB_33_28;
  reg        [7:0]    _zz_io_MatrixB_33_29;
  reg        [7:0]    _zz_io_MatrixB_33_30;
  reg        [7:0]    _zz_io_MatrixB_33_31;
  reg        [7:0]    _zz_io_MatrixB_33_32;
  reg                 _zz_io_B_Valid_33;
  reg                 _zz_io_B_Valid_33_1;
  reg                 _zz_io_B_Valid_33_2;
  reg                 _zz_io_B_Valid_33_3;
  reg                 _zz_io_B_Valid_33_4;
  reg                 _zz_io_B_Valid_33_5;
  reg                 _zz_io_B_Valid_33_6;
  reg                 _zz_io_B_Valid_33_7;
  reg                 _zz_io_B_Valid_33_8;
  reg                 _zz_io_B_Valid_33_9;
  reg                 _zz_io_B_Valid_33_10;
  reg                 _zz_io_B_Valid_33_11;
  reg                 _zz_io_B_Valid_33_12;
  reg                 _zz_io_B_Valid_33_13;
  reg                 _zz_io_B_Valid_33_14;
  reg                 _zz_io_B_Valid_33_15;
  reg                 _zz_io_B_Valid_33_16;
  reg                 _zz_io_B_Valid_33_17;
  reg                 _zz_io_B_Valid_33_18;
  reg                 _zz_io_B_Valid_33_19;
  reg                 _zz_io_B_Valid_33_20;
  reg                 _zz_io_B_Valid_33_21;
  reg                 _zz_io_B_Valid_33_22;
  reg                 _zz_io_B_Valid_33_23;
  reg                 _zz_io_B_Valid_33_24;
  reg                 _zz_io_B_Valid_33_25;
  reg                 _zz_io_B_Valid_33_26;
  reg                 _zz_io_B_Valid_33_27;
  reg                 _zz_io_B_Valid_33_28;
  reg                 _zz_io_B_Valid_33_29;
  reg                 _zz_io_B_Valid_33_30;
  reg                 _zz_io_B_Valid_33_31;
  reg                 _zz_io_B_Valid_33_32;
  reg        [7:0]    _zz_io_MatrixB_34;
  reg        [7:0]    _zz_io_MatrixB_34_1;
  reg        [7:0]    _zz_io_MatrixB_34_2;
  reg        [7:0]    _zz_io_MatrixB_34_3;
  reg        [7:0]    _zz_io_MatrixB_34_4;
  reg        [7:0]    _zz_io_MatrixB_34_5;
  reg        [7:0]    _zz_io_MatrixB_34_6;
  reg        [7:0]    _zz_io_MatrixB_34_7;
  reg        [7:0]    _zz_io_MatrixB_34_8;
  reg        [7:0]    _zz_io_MatrixB_34_9;
  reg        [7:0]    _zz_io_MatrixB_34_10;
  reg        [7:0]    _zz_io_MatrixB_34_11;
  reg        [7:0]    _zz_io_MatrixB_34_12;
  reg        [7:0]    _zz_io_MatrixB_34_13;
  reg        [7:0]    _zz_io_MatrixB_34_14;
  reg        [7:0]    _zz_io_MatrixB_34_15;
  reg        [7:0]    _zz_io_MatrixB_34_16;
  reg        [7:0]    _zz_io_MatrixB_34_17;
  reg        [7:0]    _zz_io_MatrixB_34_18;
  reg        [7:0]    _zz_io_MatrixB_34_19;
  reg        [7:0]    _zz_io_MatrixB_34_20;
  reg        [7:0]    _zz_io_MatrixB_34_21;
  reg        [7:0]    _zz_io_MatrixB_34_22;
  reg        [7:0]    _zz_io_MatrixB_34_23;
  reg        [7:0]    _zz_io_MatrixB_34_24;
  reg        [7:0]    _zz_io_MatrixB_34_25;
  reg        [7:0]    _zz_io_MatrixB_34_26;
  reg        [7:0]    _zz_io_MatrixB_34_27;
  reg        [7:0]    _zz_io_MatrixB_34_28;
  reg        [7:0]    _zz_io_MatrixB_34_29;
  reg        [7:0]    _zz_io_MatrixB_34_30;
  reg        [7:0]    _zz_io_MatrixB_34_31;
  reg        [7:0]    _zz_io_MatrixB_34_32;
  reg        [7:0]    _zz_io_MatrixB_34_33;
  reg                 _zz_io_B_Valid_34;
  reg                 _zz_io_B_Valid_34_1;
  reg                 _zz_io_B_Valid_34_2;
  reg                 _zz_io_B_Valid_34_3;
  reg                 _zz_io_B_Valid_34_4;
  reg                 _zz_io_B_Valid_34_5;
  reg                 _zz_io_B_Valid_34_6;
  reg                 _zz_io_B_Valid_34_7;
  reg                 _zz_io_B_Valid_34_8;
  reg                 _zz_io_B_Valid_34_9;
  reg                 _zz_io_B_Valid_34_10;
  reg                 _zz_io_B_Valid_34_11;
  reg                 _zz_io_B_Valid_34_12;
  reg                 _zz_io_B_Valid_34_13;
  reg                 _zz_io_B_Valid_34_14;
  reg                 _zz_io_B_Valid_34_15;
  reg                 _zz_io_B_Valid_34_16;
  reg                 _zz_io_B_Valid_34_17;
  reg                 _zz_io_B_Valid_34_18;
  reg                 _zz_io_B_Valid_34_19;
  reg                 _zz_io_B_Valid_34_20;
  reg                 _zz_io_B_Valid_34_21;
  reg                 _zz_io_B_Valid_34_22;
  reg                 _zz_io_B_Valid_34_23;
  reg                 _zz_io_B_Valid_34_24;
  reg                 _zz_io_B_Valid_34_25;
  reg                 _zz_io_B_Valid_34_26;
  reg                 _zz_io_B_Valid_34_27;
  reg                 _zz_io_B_Valid_34_28;
  reg                 _zz_io_B_Valid_34_29;
  reg                 _zz_io_B_Valid_34_30;
  reg                 _zz_io_B_Valid_34_31;
  reg                 _zz_io_B_Valid_34_32;
  reg                 _zz_io_B_Valid_34_33;
  reg        [7:0]    _zz_io_MatrixB_35;
  reg        [7:0]    _zz_io_MatrixB_35_1;
  reg        [7:0]    _zz_io_MatrixB_35_2;
  reg        [7:0]    _zz_io_MatrixB_35_3;
  reg        [7:0]    _zz_io_MatrixB_35_4;
  reg        [7:0]    _zz_io_MatrixB_35_5;
  reg        [7:0]    _zz_io_MatrixB_35_6;
  reg        [7:0]    _zz_io_MatrixB_35_7;
  reg        [7:0]    _zz_io_MatrixB_35_8;
  reg        [7:0]    _zz_io_MatrixB_35_9;
  reg        [7:0]    _zz_io_MatrixB_35_10;
  reg        [7:0]    _zz_io_MatrixB_35_11;
  reg        [7:0]    _zz_io_MatrixB_35_12;
  reg        [7:0]    _zz_io_MatrixB_35_13;
  reg        [7:0]    _zz_io_MatrixB_35_14;
  reg        [7:0]    _zz_io_MatrixB_35_15;
  reg        [7:0]    _zz_io_MatrixB_35_16;
  reg        [7:0]    _zz_io_MatrixB_35_17;
  reg        [7:0]    _zz_io_MatrixB_35_18;
  reg        [7:0]    _zz_io_MatrixB_35_19;
  reg        [7:0]    _zz_io_MatrixB_35_20;
  reg        [7:0]    _zz_io_MatrixB_35_21;
  reg        [7:0]    _zz_io_MatrixB_35_22;
  reg        [7:0]    _zz_io_MatrixB_35_23;
  reg        [7:0]    _zz_io_MatrixB_35_24;
  reg        [7:0]    _zz_io_MatrixB_35_25;
  reg        [7:0]    _zz_io_MatrixB_35_26;
  reg        [7:0]    _zz_io_MatrixB_35_27;
  reg        [7:0]    _zz_io_MatrixB_35_28;
  reg        [7:0]    _zz_io_MatrixB_35_29;
  reg        [7:0]    _zz_io_MatrixB_35_30;
  reg        [7:0]    _zz_io_MatrixB_35_31;
  reg        [7:0]    _zz_io_MatrixB_35_32;
  reg        [7:0]    _zz_io_MatrixB_35_33;
  reg        [7:0]    _zz_io_MatrixB_35_34;
  reg                 _zz_io_B_Valid_35;
  reg                 _zz_io_B_Valid_35_1;
  reg                 _zz_io_B_Valid_35_2;
  reg                 _zz_io_B_Valid_35_3;
  reg                 _zz_io_B_Valid_35_4;
  reg                 _zz_io_B_Valid_35_5;
  reg                 _zz_io_B_Valid_35_6;
  reg                 _zz_io_B_Valid_35_7;
  reg                 _zz_io_B_Valid_35_8;
  reg                 _zz_io_B_Valid_35_9;
  reg                 _zz_io_B_Valid_35_10;
  reg                 _zz_io_B_Valid_35_11;
  reg                 _zz_io_B_Valid_35_12;
  reg                 _zz_io_B_Valid_35_13;
  reg                 _zz_io_B_Valid_35_14;
  reg                 _zz_io_B_Valid_35_15;
  reg                 _zz_io_B_Valid_35_16;
  reg                 _zz_io_B_Valid_35_17;
  reg                 _zz_io_B_Valid_35_18;
  reg                 _zz_io_B_Valid_35_19;
  reg                 _zz_io_B_Valid_35_20;
  reg                 _zz_io_B_Valid_35_21;
  reg                 _zz_io_B_Valid_35_22;
  reg                 _zz_io_B_Valid_35_23;
  reg                 _zz_io_B_Valid_35_24;
  reg                 _zz_io_B_Valid_35_25;
  reg                 _zz_io_B_Valid_35_26;
  reg                 _zz_io_B_Valid_35_27;
  reg                 _zz_io_B_Valid_35_28;
  reg                 _zz_io_B_Valid_35_29;
  reg                 _zz_io_B_Valid_35_30;
  reg                 _zz_io_B_Valid_35_31;
  reg                 _zz_io_B_Valid_35_32;
  reg                 _zz_io_B_Valid_35_33;
  reg                 _zz_io_B_Valid_35_34;
  reg        [7:0]    _zz_io_MatrixB_36;
  reg        [7:0]    _zz_io_MatrixB_36_1;
  reg        [7:0]    _zz_io_MatrixB_36_2;
  reg        [7:0]    _zz_io_MatrixB_36_3;
  reg        [7:0]    _zz_io_MatrixB_36_4;
  reg        [7:0]    _zz_io_MatrixB_36_5;
  reg        [7:0]    _zz_io_MatrixB_36_6;
  reg        [7:0]    _zz_io_MatrixB_36_7;
  reg        [7:0]    _zz_io_MatrixB_36_8;
  reg        [7:0]    _zz_io_MatrixB_36_9;
  reg        [7:0]    _zz_io_MatrixB_36_10;
  reg        [7:0]    _zz_io_MatrixB_36_11;
  reg        [7:0]    _zz_io_MatrixB_36_12;
  reg        [7:0]    _zz_io_MatrixB_36_13;
  reg        [7:0]    _zz_io_MatrixB_36_14;
  reg        [7:0]    _zz_io_MatrixB_36_15;
  reg        [7:0]    _zz_io_MatrixB_36_16;
  reg        [7:0]    _zz_io_MatrixB_36_17;
  reg        [7:0]    _zz_io_MatrixB_36_18;
  reg        [7:0]    _zz_io_MatrixB_36_19;
  reg        [7:0]    _zz_io_MatrixB_36_20;
  reg        [7:0]    _zz_io_MatrixB_36_21;
  reg        [7:0]    _zz_io_MatrixB_36_22;
  reg        [7:0]    _zz_io_MatrixB_36_23;
  reg        [7:0]    _zz_io_MatrixB_36_24;
  reg        [7:0]    _zz_io_MatrixB_36_25;
  reg        [7:0]    _zz_io_MatrixB_36_26;
  reg        [7:0]    _zz_io_MatrixB_36_27;
  reg        [7:0]    _zz_io_MatrixB_36_28;
  reg        [7:0]    _zz_io_MatrixB_36_29;
  reg        [7:0]    _zz_io_MatrixB_36_30;
  reg        [7:0]    _zz_io_MatrixB_36_31;
  reg        [7:0]    _zz_io_MatrixB_36_32;
  reg        [7:0]    _zz_io_MatrixB_36_33;
  reg        [7:0]    _zz_io_MatrixB_36_34;
  reg        [7:0]    _zz_io_MatrixB_36_35;
  reg                 _zz_io_B_Valid_36;
  reg                 _zz_io_B_Valid_36_1;
  reg                 _zz_io_B_Valid_36_2;
  reg                 _zz_io_B_Valid_36_3;
  reg                 _zz_io_B_Valid_36_4;
  reg                 _zz_io_B_Valid_36_5;
  reg                 _zz_io_B_Valid_36_6;
  reg                 _zz_io_B_Valid_36_7;
  reg                 _zz_io_B_Valid_36_8;
  reg                 _zz_io_B_Valid_36_9;
  reg                 _zz_io_B_Valid_36_10;
  reg                 _zz_io_B_Valid_36_11;
  reg                 _zz_io_B_Valid_36_12;
  reg                 _zz_io_B_Valid_36_13;
  reg                 _zz_io_B_Valid_36_14;
  reg                 _zz_io_B_Valid_36_15;
  reg                 _zz_io_B_Valid_36_16;
  reg                 _zz_io_B_Valid_36_17;
  reg                 _zz_io_B_Valid_36_18;
  reg                 _zz_io_B_Valid_36_19;
  reg                 _zz_io_B_Valid_36_20;
  reg                 _zz_io_B_Valid_36_21;
  reg                 _zz_io_B_Valid_36_22;
  reg                 _zz_io_B_Valid_36_23;
  reg                 _zz_io_B_Valid_36_24;
  reg                 _zz_io_B_Valid_36_25;
  reg                 _zz_io_B_Valid_36_26;
  reg                 _zz_io_B_Valid_36_27;
  reg                 _zz_io_B_Valid_36_28;
  reg                 _zz_io_B_Valid_36_29;
  reg                 _zz_io_B_Valid_36_30;
  reg                 _zz_io_B_Valid_36_31;
  reg                 _zz_io_B_Valid_36_32;
  reg                 _zz_io_B_Valid_36_33;
  reg                 _zz_io_B_Valid_36_34;
  reg                 _zz_io_B_Valid_36_35;
  reg        [7:0]    _zz_io_MatrixB_37;
  reg        [7:0]    _zz_io_MatrixB_37_1;
  reg        [7:0]    _zz_io_MatrixB_37_2;
  reg        [7:0]    _zz_io_MatrixB_37_3;
  reg        [7:0]    _zz_io_MatrixB_37_4;
  reg        [7:0]    _zz_io_MatrixB_37_5;
  reg        [7:0]    _zz_io_MatrixB_37_6;
  reg        [7:0]    _zz_io_MatrixB_37_7;
  reg        [7:0]    _zz_io_MatrixB_37_8;
  reg        [7:0]    _zz_io_MatrixB_37_9;
  reg        [7:0]    _zz_io_MatrixB_37_10;
  reg        [7:0]    _zz_io_MatrixB_37_11;
  reg        [7:0]    _zz_io_MatrixB_37_12;
  reg        [7:0]    _zz_io_MatrixB_37_13;
  reg        [7:0]    _zz_io_MatrixB_37_14;
  reg        [7:0]    _zz_io_MatrixB_37_15;
  reg        [7:0]    _zz_io_MatrixB_37_16;
  reg        [7:0]    _zz_io_MatrixB_37_17;
  reg        [7:0]    _zz_io_MatrixB_37_18;
  reg        [7:0]    _zz_io_MatrixB_37_19;
  reg        [7:0]    _zz_io_MatrixB_37_20;
  reg        [7:0]    _zz_io_MatrixB_37_21;
  reg        [7:0]    _zz_io_MatrixB_37_22;
  reg        [7:0]    _zz_io_MatrixB_37_23;
  reg        [7:0]    _zz_io_MatrixB_37_24;
  reg        [7:0]    _zz_io_MatrixB_37_25;
  reg        [7:0]    _zz_io_MatrixB_37_26;
  reg        [7:0]    _zz_io_MatrixB_37_27;
  reg        [7:0]    _zz_io_MatrixB_37_28;
  reg        [7:0]    _zz_io_MatrixB_37_29;
  reg        [7:0]    _zz_io_MatrixB_37_30;
  reg        [7:0]    _zz_io_MatrixB_37_31;
  reg        [7:0]    _zz_io_MatrixB_37_32;
  reg        [7:0]    _zz_io_MatrixB_37_33;
  reg        [7:0]    _zz_io_MatrixB_37_34;
  reg        [7:0]    _zz_io_MatrixB_37_35;
  reg        [7:0]    _zz_io_MatrixB_37_36;
  reg                 _zz_io_B_Valid_37;
  reg                 _zz_io_B_Valid_37_1;
  reg                 _zz_io_B_Valid_37_2;
  reg                 _zz_io_B_Valid_37_3;
  reg                 _zz_io_B_Valid_37_4;
  reg                 _zz_io_B_Valid_37_5;
  reg                 _zz_io_B_Valid_37_6;
  reg                 _zz_io_B_Valid_37_7;
  reg                 _zz_io_B_Valid_37_8;
  reg                 _zz_io_B_Valid_37_9;
  reg                 _zz_io_B_Valid_37_10;
  reg                 _zz_io_B_Valid_37_11;
  reg                 _zz_io_B_Valid_37_12;
  reg                 _zz_io_B_Valid_37_13;
  reg                 _zz_io_B_Valid_37_14;
  reg                 _zz_io_B_Valid_37_15;
  reg                 _zz_io_B_Valid_37_16;
  reg                 _zz_io_B_Valid_37_17;
  reg                 _zz_io_B_Valid_37_18;
  reg                 _zz_io_B_Valid_37_19;
  reg                 _zz_io_B_Valid_37_20;
  reg                 _zz_io_B_Valid_37_21;
  reg                 _zz_io_B_Valid_37_22;
  reg                 _zz_io_B_Valid_37_23;
  reg                 _zz_io_B_Valid_37_24;
  reg                 _zz_io_B_Valid_37_25;
  reg                 _zz_io_B_Valid_37_26;
  reg                 _zz_io_B_Valid_37_27;
  reg                 _zz_io_B_Valid_37_28;
  reg                 _zz_io_B_Valid_37_29;
  reg                 _zz_io_B_Valid_37_30;
  reg                 _zz_io_B_Valid_37_31;
  reg                 _zz_io_B_Valid_37_32;
  reg                 _zz_io_B_Valid_37_33;
  reg                 _zz_io_B_Valid_37_34;
  reg                 _zz_io_B_Valid_37_35;
  reg                 _zz_io_B_Valid_37_36;
  reg        [7:0]    _zz_io_MatrixB_38;
  reg        [7:0]    _zz_io_MatrixB_38_1;
  reg        [7:0]    _zz_io_MatrixB_38_2;
  reg        [7:0]    _zz_io_MatrixB_38_3;
  reg        [7:0]    _zz_io_MatrixB_38_4;
  reg        [7:0]    _zz_io_MatrixB_38_5;
  reg        [7:0]    _zz_io_MatrixB_38_6;
  reg        [7:0]    _zz_io_MatrixB_38_7;
  reg        [7:0]    _zz_io_MatrixB_38_8;
  reg        [7:0]    _zz_io_MatrixB_38_9;
  reg        [7:0]    _zz_io_MatrixB_38_10;
  reg        [7:0]    _zz_io_MatrixB_38_11;
  reg        [7:0]    _zz_io_MatrixB_38_12;
  reg        [7:0]    _zz_io_MatrixB_38_13;
  reg        [7:0]    _zz_io_MatrixB_38_14;
  reg        [7:0]    _zz_io_MatrixB_38_15;
  reg        [7:0]    _zz_io_MatrixB_38_16;
  reg        [7:0]    _zz_io_MatrixB_38_17;
  reg        [7:0]    _zz_io_MatrixB_38_18;
  reg        [7:0]    _zz_io_MatrixB_38_19;
  reg        [7:0]    _zz_io_MatrixB_38_20;
  reg        [7:0]    _zz_io_MatrixB_38_21;
  reg        [7:0]    _zz_io_MatrixB_38_22;
  reg        [7:0]    _zz_io_MatrixB_38_23;
  reg        [7:0]    _zz_io_MatrixB_38_24;
  reg        [7:0]    _zz_io_MatrixB_38_25;
  reg        [7:0]    _zz_io_MatrixB_38_26;
  reg        [7:0]    _zz_io_MatrixB_38_27;
  reg        [7:0]    _zz_io_MatrixB_38_28;
  reg        [7:0]    _zz_io_MatrixB_38_29;
  reg        [7:0]    _zz_io_MatrixB_38_30;
  reg        [7:0]    _zz_io_MatrixB_38_31;
  reg        [7:0]    _zz_io_MatrixB_38_32;
  reg        [7:0]    _zz_io_MatrixB_38_33;
  reg        [7:0]    _zz_io_MatrixB_38_34;
  reg        [7:0]    _zz_io_MatrixB_38_35;
  reg        [7:0]    _zz_io_MatrixB_38_36;
  reg        [7:0]    _zz_io_MatrixB_38_37;
  reg                 _zz_io_B_Valid_38;
  reg                 _zz_io_B_Valid_38_1;
  reg                 _zz_io_B_Valid_38_2;
  reg                 _zz_io_B_Valid_38_3;
  reg                 _zz_io_B_Valid_38_4;
  reg                 _zz_io_B_Valid_38_5;
  reg                 _zz_io_B_Valid_38_6;
  reg                 _zz_io_B_Valid_38_7;
  reg                 _zz_io_B_Valid_38_8;
  reg                 _zz_io_B_Valid_38_9;
  reg                 _zz_io_B_Valid_38_10;
  reg                 _zz_io_B_Valid_38_11;
  reg                 _zz_io_B_Valid_38_12;
  reg                 _zz_io_B_Valid_38_13;
  reg                 _zz_io_B_Valid_38_14;
  reg                 _zz_io_B_Valid_38_15;
  reg                 _zz_io_B_Valid_38_16;
  reg                 _zz_io_B_Valid_38_17;
  reg                 _zz_io_B_Valid_38_18;
  reg                 _zz_io_B_Valid_38_19;
  reg                 _zz_io_B_Valid_38_20;
  reg                 _zz_io_B_Valid_38_21;
  reg                 _zz_io_B_Valid_38_22;
  reg                 _zz_io_B_Valid_38_23;
  reg                 _zz_io_B_Valid_38_24;
  reg                 _zz_io_B_Valid_38_25;
  reg                 _zz_io_B_Valid_38_26;
  reg                 _zz_io_B_Valid_38_27;
  reg                 _zz_io_B_Valid_38_28;
  reg                 _zz_io_B_Valid_38_29;
  reg                 _zz_io_B_Valid_38_30;
  reg                 _zz_io_B_Valid_38_31;
  reg                 _zz_io_B_Valid_38_32;
  reg                 _zz_io_B_Valid_38_33;
  reg                 _zz_io_B_Valid_38_34;
  reg                 _zz_io_B_Valid_38_35;
  reg                 _zz_io_B_Valid_38_36;
  reg                 _zz_io_B_Valid_38_37;
  reg        [7:0]    _zz_io_MatrixB_39;
  reg        [7:0]    _zz_io_MatrixB_39_1;
  reg        [7:0]    _zz_io_MatrixB_39_2;
  reg        [7:0]    _zz_io_MatrixB_39_3;
  reg        [7:0]    _zz_io_MatrixB_39_4;
  reg        [7:0]    _zz_io_MatrixB_39_5;
  reg        [7:0]    _zz_io_MatrixB_39_6;
  reg        [7:0]    _zz_io_MatrixB_39_7;
  reg        [7:0]    _zz_io_MatrixB_39_8;
  reg        [7:0]    _zz_io_MatrixB_39_9;
  reg        [7:0]    _zz_io_MatrixB_39_10;
  reg        [7:0]    _zz_io_MatrixB_39_11;
  reg        [7:0]    _zz_io_MatrixB_39_12;
  reg        [7:0]    _zz_io_MatrixB_39_13;
  reg        [7:0]    _zz_io_MatrixB_39_14;
  reg        [7:0]    _zz_io_MatrixB_39_15;
  reg        [7:0]    _zz_io_MatrixB_39_16;
  reg        [7:0]    _zz_io_MatrixB_39_17;
  reg        [7:0]    _zz_io_MatrixB_39_18;
  reg        [7:0]    _zz_io_MatrixB_39_19;
  reg        [7:0]    _zz_io_MatrixB_39_20;
  reg        [7:0]    _zz_io_MatrixB_39_21;
  reg        [7:0]    _zz_io_MatrixB_39_22;
  reg        [7:0]    _zz_io_MatrixB_39_23;
  reg        [7:0]    _zz_io_MatrixB_39_24;
  reg        [7:0]    _zz_io_MatrixB_39_25;
  reg        [7:0]    _zz_io_MatrixB_39_26;
  reg        [7:0]    _zz_io_MatrixB_39_27;
  reg        [7:0]    _zz_io_MatrixB_39_28;
  reg        [7:0]    _zz_io_MatrixB_39_29;
  reg        [7:0]    _zz_io_MatrixB_39_30;
  reg        [7:0]    _zz_io_MatrixB_39_31;
  reg        [7:0]    _zz_io_MatrixB_39_32;
  reg        [7:0]    _zz_io_MatrixB_39_33;
  reg        [7:0]    _zz_io_MatrixB_39_34;
  reg        [7:0]    _zz_io_MatrixB_39_35;
  reg        [7:0]    _zz_io_MatrixB_39_36;
  reg        [7:0]    _zz_io_MatrixB_39_37;
  reg        [7:0]    _zz_io_MatrixB_39_38;
  reg                 _zz_io_B_Valid_39;
  reg                 _zz_io_B_Valid_39_1;
  reg                 _zz_io_B_Valid_39_2;
  reg                 _zz_io_B_Valid_39_3;
  reg                 _zz_io_B_Valid_39_4;
  reg                 _zz_io_B_Valid_39_5;
  reg                 _zz_io_B_Valid_39_6;
  reg                 _zz_io_B_Valid_39_7;
  reg                 _zz_io_B_Valid_39_8;
  reg                 _zz_io_B_Valid_39_9;
  reg                 _zz_io_B_Valid_39_10;
  reg                 _zz_io_B_Valid_39_11;
  reg                 _zz_io_B_Valid_39_12;
  reg                 _zz_io_B_Valid_39_13;
  reg                 _zz_io_B_Valid_39_14;
  reg                 _zz_io_B_Valid_39_15;
  reg                 _zz_io_B_Valid_39_16;
  reg                 _zz_io_B_Valid_39_17;
  reg                 _zz_io_B_Valid_39_18;
  reg                 _zz_io_B_Valid_39_19;
  reg                 _zz_io_B_Valid_39_20;
  reg                 _zz_io_B_Valid_39_21;
  reg                 _zz_io_B_Valid_39_22;
  reg                 _zz_io_B_Valid_39_23;
  reg                 _zz_io_B_Valid_39_24;
  reg                 _zz_io_B_Valid_39_25;
  reg                 _zz_io_B_Valid_39_26;
  reg                 _zz_io_B_Valid_39_27;
  reg                 _zz_io_B_Valid_39_28;
  reg                 _zz_io_B_Valid_39_29;
  reg                 _zz_io_B_Valid_39_30;
  reg                 _zz_io_B_Valid_39_31;
  reg                 _zz_io_B_Valid_39_32;
  reg                 _zz_io_B_Valid_39_33;
  reg                 _zz_io_B_Valid_39_34;
  reg                 _zz_io_B_Valid_39_35;
  reg                 _zz_io_B_Valid_39_36;
  reg                 _zz_io_B_Valid_39_37;
  reg                 _zz_io_B_Valid_39_38;
  reg        [7:0]    _zz_io_MatrixB_40;
  reg        [7:0]    _zz_io_MatrixB_40_1;
  reg        [7:0]    _zz_io_MatrixB_40_2;
  reg        [7:0]    _zz_io_MatrixB_40_3;
  reg        [7:0]    _zz_io_MatrixB_40_4;
  reg        [7:0]    _zz_io_MatrixB_40_5;
  reg        [7:0]    _zz_io_MatrixB_40_6;
  reg        [7:0]    _zz_io_MatrixB_40_7;
  reg        [7:0]    _zz_io_MatrixB_40_8;
  reg        [7:0]    _zz_io_MatrixB_40_9;
  reg        [7:0]    _zz_io_MatrixB_40_10;
  reg        [7:0]    _zz_io_MatrixB_40_11;
  reg        [7:0]    _zz_io_MatrixB_40_12;
  reg        [7:0]    _zz_io_MatrixB_40_13;
  reg        [7:0]    _zz_io_MatrixB_40_14;
  reg        [7:0]    _zz_io_MatrixB_40_15;
  reg        [7:0]    _zz_io_MatrixB_40_16;
  reg        [7:0]    _zz_io_MatrixB_40_17;
  reg        [7:0]    _zz_io_MatrixB_40_18;
  reg        [7:0]    _zz_io_MatrixB_40_19;
  reg        [7:0]    _zz_io_MatrixB_40_20;
  reg        [7:0]    _zz_io_MatrixB_40_21;
  reg        [7:0]    _zz_io_MatrixB_40_22;
  reg        [7:0]    _zz_io_MatrixB_40_23;
  reg        [7:0]    _zz_io_MatrixB_40_24;
  reg        [7:0]    _zz_io_MatrixB_40_25;
  reg        [7:0]    _zz_io_MatrixB_40_26;
  reg        [7:0]    _zz_io_MatrixB_40_27;
  reg        [7:0]    _zz_io_MatrixB_40_28;
  reg        [7:0]    _zz_io_MatrixB_40_29;
  reg        [7:0]    _zz_io_MatrixB_40_30;
  reg        [7:0]    _zz_io_MatrixB_40_31;
  reg        [7:0]    _zz_io_MatrixB_40_32;
  reg        [7:0]    _zz_io_MatrixB_40_33;
  reg        [7:0]    _zz_io_MatrixB_40_34;
  reg        [7:0]    _zz_io_MatrixB_40_35;
  reg        [7:0]    _zz_io_MatrixB_40_36;
  reg        [7:0]    _zz_io_MatrixB_40_37;
  reg        [7:0]    _zz_io_MatrixB_40_38;
  reg        [7:0]    _zz_io_MatrixB_40_39;
  reg                 _zz_io_B_Valid_40;
  reg                 _zz_io_B_Valid_40_1;
  reg                 _zz_io_B_Valid_40_2;
  reg                 _zz_io_B_Valid_40_3;
  reg                 _zz_io_B_Valid_40_4;
  reg                 _zz_io_B_Valid_40_5;
  reg                 _zz_io_B_Valid_40_6;
  reg                 _zz_io_B_Valid_40_7;
  reg                 _zz_io_B_Valid_40_8;
  reg                 _zz_io_B_Valid_40_9;
  reg                 _zz_io_B_Valid_40_10;
  reg                 _zz_io_B_Valid_40_11;
  reg                 _zz_io_B_Valid_40_12;
  reg                 _zz_io_B_Valid_40_13;
  reg                 _zz_io_B_Valid_40_14;
  reg                 _zz_io_B_Valid_40_15;
  reg                 _zz_io_B_Valid_40_16;
  reg                 _zz_io_B_Valid_40_17;
  reg                 _zz_io_B_Valid_40_18;
  reg                 _zz_io_B_Valid_40_19;
  reg                 _zz_io_B_Valid_40_20;
  reg                 _zz_io_B_Valid_40_21;
  reg                 _zz_io_B_Valid_40_22;
  reg                 _zz_io_B_Valid_40_23;
  reg                 _zz_io_B_Valid_40_24;
  reg                 _zz_io_B_Valid_40_25;
  reg                 _zz_io_B_Valid_40_26;
  reg                 _zz_io_B_Valid_40_27;
  reg                 _zz_io_B_Valid_40_28;
  reg                 _zz_io_B_Valid_40_29;
  reg                 _zz_io_B_Valid_40_30;
  reg                 _zz_io_B_Valid_40_31;
  reg                 _zz_io_B_Valid_40_32;
  reg                 _zz_io_B_Valid_40_33;
  reg                 _zz_io_B_Valid_40_34;
  reg                 _zz_io_B_Valid_40_35;
  reg                 _zz_io_B_Valid_40_36;
  reg                 _zz_io_B_Valid_40_37;
  reg                 _zz_io_B_Valid_40_38;
  reg                 _zz_io_B_Valid_40_39;
  reg        [7:0]    _zz_io_MatrixB_41;
  reg        [7:0]    _zz_io_MatrixB_41_1;
  reg        [7:0]    _zz_io_MatrixB_41_2;
  reg        [7:0]    _zz_io_MatrixB_41_3;
  reg        [7:0]    _zz_io_MatrixB_41_4;
  reg        [7:0]    _zz_io_MatrixB_41_5;
  reg        [7:0]    _zz_io_MatrixB_41_6;
  reg        [7:0]    _zz_io_MatrixB_41_7;
  reg        [7:0]    _zz_io_MatrixB_41_8;
  reg        [7:0]    _zz_io_MatrixB_41_9;
  reg        [7:0]    _zz_io_MatrixB_41_10;
  reg        [7:0]    _zz_io_MatrixB_41_11;
  reg        [7:0]    _zz_io_MatrixB_41_12;
  reg        [7:0]    _zz_io_MatrixB_41_13;
  reg        [7:0]    _zz_io_MatrixB_41_14;
  reg        [7:0]    _zz_io_MatrixB_41_15;
  reg        [7:0]    _zz_io_MatrixB_41_16;
  reg        [7:0]    _zz_io_MatrixB_41_17;
  reg        [7:0]    _zz_io_MatrixB_41_18;
  reg        [7:0]    _zz_io_MatrixB_41_19;
  reg        [7:0]    _zz_io_MatrixB_41_20;
  reg        [7:0]    _zz_io_MatrixB_41_21;
  reg        [7:0]    _zz_io_MatrixB_41_22;
  reg        [7:0]    _zz_io_MatrixB_41_23;
  reg        [7:0]    _zz_io_MatrixB_41_24;
  reg        [7:0]    _zz_io_MatrixB_41_25;
  reg        [7:0]    _zz_io_MatrixB_41_26;
  reg        [7:0]    _zz_io_MatrixB_41_27;
  reg        [7:0]    _zz_io_MatrixB_41_28;
  reg        [7:0]    _zz_io_MatrixB_41_29;
  reg        [7:0]    _zz_io_MatrixB_41_30;
  reg        [7:0]    _zz_io_MatrixB_41_31;
  reg        [7:0]    _zz_io_MatrixB_41_32;
  reg        [7:0]    _zz_io_MatrixB_41_33;
  reg        [7:0]    _zz_io_MatrixB_41_34;
  reg        [7:0]    _zz_io_MatrixB_41_35;
  reg        [7:0]    _zz_io_MatrixB_41_36;
  reg        [7:0]    _zz_io_MatrixB_41_37;
  reg        [7:0]    _zz_io_MatrixB_41_38;
  reg        [7:0]    _zz_io_MatrixB_41_39;
  reg        [7:0]    _zz_io_MatrixB_41_40;
  reg                 _zz_io_B_Valid_41;
  reg                 _zz_io_B_Valid_41_1;
  reg                 _zz_io_B_Valid_41_2;
  reg                 _zz_io_B_Valid_41_3;
  reg                 _zz_io_B_Valid_41_4;
  reg                 _zz_io_B_Valid_41_5;
  reg                 _zz_io_B_Valid_41_6;
  reg                 _zz_io_B_Valid_41_7;
  reg                 _zz_io_B_Valid_41_8;
  reg                 _zz_io_B_Valid_41_9;
  reg                 _zz_io_B_Valid_41_10;
  reg                 _zz_io_B_Valid_41_11;
  reg                 _zz_io_B_Valid_41_12;
  reg                 _zz_io_B_Valid_41_13;
  reg                 _zz_io_B_Valid_41_14;
  reg                 _zz_io_B_Valid_41_15;
  reg                 _zz_io_B_Valid_41_16;
  reg                 _zz_io_B_Valid_41_17;
  reg                 _zz_io_B_Valid_41_18;
  reg                 _zz_io_B_Valid_41_19;
  reg                 _zz_io_B_Valid_41_20;
  reg                 _zz_io_B_Valid_41_21;
  reg                 _zz_io_B_Valid_41_22;
  reg                 _zz_io_B_Valid_41_23;
  reg                 _zz_io_B_Valid_41_24;
  reg                 _zz_io_B_Valid_41_25;
  reg                 _zz_io_B_Valid_41_26;
  reg                 _zz_io_B_Valid_41_27;
  reg                 _zz_io_B_Valid_41_28;
  reg                 _zz_io_B_Valid_41_29;
  reg                 _zz_io_B_Valid_41_30;
  reg                 _zz_io_B_Valid_41_31;
  reg                 _zz_io_B_Valid_41_32;
  reg                 _zz_io_B_Valid_41_33;
  reg                 _zz_io_B_Valid_41_34;
  reg                 _zz_io_B_Valid_41_35;
  reg                 _zz_io_B_Valid_41_36;
  reg                 _zz_io_B_Valid_41_37;
  reg                 _zz_io_B_Valid_41_38;
  reg                 _zz_io_B_Valid_41_39;
  reg                 _zz_io_B_Valid_41_40;
  reg        [7:0]    _zz_io_MatrixB_42;
  reg        [7:0]    _zz_io_MatrixB_42_1;
  reg        [7:0]    _zz_io_MatrixB_42_2;
  reg        [7:0]    _zz_io_MatrixB_42_3;
  reg        [7:0]    _zz_io_MatrixB_42_4;
  reg        [7:0]    _zz_io_MatrixB_42_5;
  reg        [7:0]    _zz_io_MatrixB_42_6;
  reg        [7:0]    _zz_io_MatrixB_42_7;
  reg        [7:0]    _zz_io_MatrixB_42_8;
  reg        [7:0]    _zz_io_MatrixB_42_9;
  reg        [7:0]    _zz_io_MatrixB_42_10;
  reg        [7:0]    _zz_io_MatrixB_42_11;
  reg        [7:0]    _zz_io_MatrixB_42_12;
  reg        [7:0]    _zz_io_MatrixB_42_13;
  reg        [7:0]    _zz_io_MatrixB_42_14;
  reg        [7:0]    _zz_io_MatrixB_42_15;
  reg        [7:0]    _zz_io_MatrixB_42_16;
  reg        [7:0]    _zz_io_MatrixB_42_17;
  reg        [7:0]    _zz_io_MatrixB_42_18;
  reg        [7:0]    _zz_io_MatrixB_42_19;
  reg        [7:0]    _zz_io_MatrixB_42_20;
  reg        [7:0]    _zz_io_MatrixB_42_21;
  reg        [7:0]    _zz_io_MatrixB_42_22;
  reg        [7:0]    _zz_io_MatrixB_42_23;
  reg        [7:0]    _zz_io_MatrixB_42_24;
  reg        [7:0]    _zz_io_MatrixB_42_25;
  reg        [7:0]    _zz_io_MatrixB_42_26;
  reg        [7:0]    _zz_io_MatrixB_42_27;
  reg        [7:0]    _zz_io_MatrixB_42_28;
  reg        [7:0]    _zz_io_MatrixB_42_29;
  reg        [7:0]    _zz_io_MatrixB_42_30;
  reg        [7:0]    _zz_io_MatrixB_42_31;
  reg        [7:0]    _zz_io_MatrixB_42_32;
  reg        [7:0]    _zz_io_MatrixB_42_33;
  reg        [7:0]    _zz_io_MatrixB_42_34;
  reg        [7:0]    _zz_io_MatrixB_42_35;
  reg        [7:0]    _zz_io_MatrixB_42_36;
  reg        [7:0]    _zz_io_MatrixB_42_37;
  reg        [7:0]    _zz_io_MatrixB_42_38;
  reg        [7:0]    _zz_io_MatrixB_42_39;
  reg        [7:0]    _zz_io_MatrixB_42_40;
  reg        [7:0]    _zz_io_MatrixB_42_41;
  reg                 _zz_io_B_Valid_42;
  reg                 _zz_io_B_Valid_42_1;
  reg                 _zz_io_B_Valid_42_2;
  reg                 _zz_io_B_Valid_42_3;
  reg                 _zz_io_B_Valid_42_4;
  reg                 _zz_io_B_Valid_42_5;
  reg                 _zz_io_B_Valid_42_6;
  reg                 _zz_io_B_Valid_42_7;
  reg                 _zz_io_B_Valid_42_8;
  reg                 _zz_io_B_Valid_42_9;
  reg                 _zz_io_B_Valid_42_10;
  reg                 _zz_io_B_Valid_42_11;
  reg                 _zz_io_B_Valid_42_12;
  reg                 _zz_io_B_Valid_42_13;
  reg                 _zz_io_B_Valid_42_14;
  reg                 _zz_io_B_Valid_42_15;
  reg                 _zz_io_B_Valid_42_16;
  reg                 _zz_io_B_Valid_42_17;
  reg                 _zz_io_B_Valid_42_18;
  reg                 _zz_io_B_Valid_42_19;
  reg                 _zz_io_B_Valid_42_20;
  reg                 _zz_io_B_Valid_42_21;
  reg                 _zz_io_B_Valid_42_22;
  reg                 _zz_io_B_Valid_42_23;
  reg                 _zz_io_B_Valid_42_24;
  reg                 _zz_io_B_Valid_42_25;
  reg                 _zz_io_B_Valid_42_26;
  reg                 _zz_io_B_Valid_42_27;
  reg                 _zz_io_B_Valid_42_28;
  reg                 _zz_io_B_Valid_42_29;
  reg                 _zz_io_B_Valid_42_30;
  reg                 _zz_io_B_Valid_42_31;
  reg                 _zz_io_B_Valid_42_32;
  reg                 _zz_io_B_Valid_42_33;
  reg                 _zz_io_B_Valid_42_34;
  reg                 _zz_io_B_Valid_42_35;
  reg                 _zz_io_B_Valid_42_36;
  reg                 _zz_io_B_Valid_42_37;
  reg                 _zz_io_B_Valid_42_38;
  reg                 _zz_io_B_Valid_42_39;
  reg                 _zz_io_B_Valid_42_40;
  reg                 _zz_io_B_Valid_42_41;
  reg        [7:0]    _zz_io_MatrixB_43;
  reg        [7:0]    _zz_io_MatrixB_43_1;
  reg        [7:0]    _zz_io_MatrixB_43_2;
  reg        [7:0]    _zz_io_MatrixB_43_3;
  reg        [7:0]    _zz_io_MatrixB_43_4;
  reg        [7:0]    _zz_io_MatrixB_43_5;
  reg        [7:0]    _zz_io_MatrixB_43_6;
  reg        [7:0]    _zz_io_MatrixB_43_7;
  reg        [7:0]    _zz_io_MatrixB_43_8;
  reg        [7:0]    _zz_io_MatrixB_43_9;
  reg        [7:0]    _zz_io_MatrixB_43_10;
  reg        [7:0]    _zz_io_MatrixB_43_11;
  reg        [7:0]    _zz_io_MatrixB_43_12;
  reg        [7:0]    _zz_io_MatrixB_43_13;
  reg        [7:0]    _zz_io_MatrixB_43_14;
  reg        [7:0]    _zz_io_MatrixB_43_15;
  reg        [7:0]    _zz_io_MatrixB_43_16;
  reg        [7:0]    _zz_io_MatrixB_43_17;
  reg        [7:0]    _zz_io_MatrixB_43_18;
  reg        [7:0]    _zz_io_MatrixB_43_19;
  reg        [7:0]    _zz_io_MatrixB_43_20;
  reg        [7:0]    _zz_io_MatrixB_43_21;
  reg        [7:0]    _zz_io_MatrixB_43_22;
  reg        [7:0]    _zz_io_MatrixB_43_23;
  reg        [7:0]    _zz_io_MatrixB_43_24;
  reg        [7:0]    _zz_io_MatrixB_43_25;
  reg        [7:0]    _zz_io_MatrixB_43_26;
  reg        [7:0]    _zz_io_MatrixB_43_27;
  reg        [7:0]    _zz_io_MatrixB_43_28;
  reg        [7:0]    _zz_io_MatrixB_43_29;
  reg        [7:0]    _zz_io_MatrixB_43_30;
  reg        [7:0]    _zz_io_MatrixB_43_31;
  reg        [7:0]    _zz_io_MatrixB_43_32;
  reg        [7:0]    _zz_io_MatrixB_43_33;
  reg        [7:0]    _zz_io_MatrixB_43_34;
  reg        [7:0]    _zz_io_MatrixB_43_35;
  reg        [7:0]    _zz_io_MatrixB_43_36;
  reg        [7:0]    _zz_io_MatrixB_43_37;
  reg        [7:0]    _zz_io_MatrixB_43_38;
  reg        [7:0]    _zz_io_MatrixB_43_39;
  reg        [7:0]    _zz_io_MatrixB_43_40;
  reg        [7:0]    _zz_io_MatrixB_43_41;
  reg        [7:0]    _zz_io_MatrixB_43_42;
  reg                 _zz_io_B_Valid_43;
  reg                 _zz_io_B_Valid_43_1;
  reg                 _zz_io_B_Valid_43_2;
  reg                 _zz_io_B_Valid_43_3;
  reg                 _zz_io_B_Valid_43_4;
  reg                 _zz_io_B_Valid_43_5;
  reg                 _zz_io_B_Valid_43_6;
  reg                 _zz_io_B_Valid_43_7;
  reg                 _zz_io_B_Valid_43_8;
  reg                 _zz_io_B_Valid_43_9;
  reg                 _zz_io_B_Valid_43_10;
  reg                 _zz_io_B_Valid_43_11;
  reg                 _zz_io_B_Valid_43_12;
  reg                 _zz_io_B_Valid_43_13;
  reg                 _zz_io_B_Valid_43_14;
  reg                 _zz_io_B_Valid_43_15;
  reg                 _zz_io_B_Valid_43_16;
  reg                 _zz_io_B_Valid_43_17;
  reg                 _zz_io_B_Valid_43_18;
  reg                 _zz_io_B_Valid_43_19;
  reg                 _zz_io_B_Valid_43_20;
  reg                 _zz_io_B_Valid_43_21;
  reg                 _zz_io_B_Valid_43_22;
  reg                 _zz_io_B_Valid_43_23;
  reg                 _zz_io_B_Valid_43_24;
  reg                 _zz_io_B_Valid_43_25;
  reg                 _zz_io_B_Valid_43_26;
  reg                 _zz_io_B_Valid_43_27;
  reg                 _zz_io_B_Valid_43_28;
  reg                 _zz_io_B_Valid_43_29;
  reg                 _zz_io_B_Valid_43_30;
  reg                 _zz_io_B_Valid_43_31;
  reg                 _zz_io_B_Valid_43_32;
  reg                 _zz_io_B_Valid_43_33;
  reg                 _zz_io_B_Valid_43_34;
  reg                 _zz_io_B_Valid_43_35;
  reg                 _zz_io_B_Valid_43_36;
  reg                 _zz_io_B_Valid_43_37;
  reg                 _zz_io_B_Valid_43_38;
  reg                 _zz_io_B_Valid_43_39;
  reg                 _zz_io_B_Valid_43_40;
  reg                 _zz_io_B_Valid_43_41;
  reg                 _zz_io_B_Valid_43_42;
  reg        [7:0]    _zz_io_MatrixB_44;
  reg        [7:0]    _zz_io_MatrixB_44_1;
  reg        [7:0]    _zz_io_MatrixB_44_2;
  reg        [7:0]    _zz_io_MatrixB_44_3;
  reg        [7:0]    _zz_io_MatrixB_44_4;
  reg        [7:0]    _zz_io_MatrixB_44_5;
  reg        [7:0]    _zz_io_MatrixB_44_6;
  reg        [7:0]    _zz_io_MatrixB_44_7;
  reg        [7:0]    _zz_io_MatrixB_44_8;
  reg        [7:0]    _zz_io_MatrixB_44_9;
  reg        [7:0]    _zz_io_MatrixB_44_10;
  reg        [7:0]    _zz_io_MatrixB_44_11;
  reg        [7:0]    _zz_io_MatrixB_44_12;
  reg        [7:0]    _zz_io_MatrixB_44_13;
  reg        [7:0]    _zz_io_MatrixB_44_14;
  reg        [7:0]    _zz_io_MatrixB_44_15;
  reg        [7:0]    _zz_io_MatrixB_44_16;
  reg        [7:0]    _zz_io_MatrixB_44_17;
  reg        [7:0]    _zz_io_MatrixB_44_18;
  reg        [7:0]    _zz_io_MatrixB_44_19;
  reg        [7:0]    _zz_io_MatrixB_44_20;
  reg        [7:0]    _zz_io_MatrixB_44_21;
  reg        [7:0]    _zz_io_MatrixB_44_22;
  reg        [7:0]    _zz_io_MatrixB_44_23;
  reg        [7:0]    _zz_io_MatrixB_44_24;
  reg        [7:0]    _zz_io_MatrixB_44_25;
  reg        [7:0]    _zz_io_MatrixB_44_26;
  reg        [7:0]    _zz_io_MatrixB_44_27;
  reg        [7:0]    _zz_io_MatrixB_44_28;
  reg        [7:0]    _zz_io_MatrixB_44_29;
  reg        [7:0]    _zz_io_MatrixB_44_30;
  reg        [7:0]    _zz_io_MatrixB_44_31;
  reg        [7:0]    _zz_io_MatrixB_44_32;
  reg        [7:0]    _zz_io_MatrixB_44_33;
  reg        [7:0]    _zz_io_MatrixB_44_34;
  reg        [7:0]    _zz_io_MatrixB_44_35;
  reg        [7:0]    _zz_io_MatrixB_44_36;
  reg        [7:0]    _zz_io_MatrixB_44_37;
  reg        [7:0]    _zz_io_MatrixB_44_38;
  reg        [7:0]    _zz_io_MatrixB_44_39;
  reg        [7:0]    _zz_io_MatrixB_44_40;
  reg        [7:0]    _zz_io_MatrixB_44_41;
  reg        [7:0]    _zz_io_MatrixB_44_42;
  reg        [7:0]    _zz_io_MatrixB_44_43;
  reg                 _zz_io_B_Valid_44;
  reg                 _zz_io_B_Valid_44_1;
  reg                 _zz_io_B_Valid_44_2;
  reg                 _zz_io_B_Valid_44_3;
  reg                 _zz_io_B_Valid_44_4;
  reg                 _zz_io_B_Valid_44_5;
  reg                 _zz_io_B_Valid_44_6;
  reg                 _zz_io_B_Valid_44_7;
  reg                 _zz_io_B_Valid_44_8;
  reg                 _zz_io_B_Valid_44_9;
  reg                 _zz_io_B_Valid_44_10;
  reg                 _zz_io_B_Valid_44_11;
  reg                 _zz_io_B_Valid_44_12;
  reg                 _zz_io_B_Valid_44_13;
  reg                 _zz_io_B_Valid_44_14;
  reg                 _zz_io_B_Valid_44_15;
  reg                 _zz_io_B_Valid_44_16;
  reg                 _zz_io_B_Valid_44_17;
  reg                 _zz_io_B_Valid_44_18;
  reg                 _zz_io_B_Valid_44_19;
  reg                 _zz_io_B_Valid_44_20;
  reg                 _zz_io_B_Valid_44_21;
  reg                 _zz_io_B_Valid_44_22;
  reg                 _zz_io_B_Valid_44_23;
  reg                 _zz_io_B_Valid_44_24;
  reg                 _zz_io_B_Valid_44_25;
  reg                 _zz_io_B_Valid_44_26;
  reg                 _zz_io_B_Valid_44_27;
  reg                 _zz_io_B_Valid_44_28;
  reg                 _zz_io_B_Valid_44_29;
  reg                 _zz_io_B_Valid_44_30;
  reg                 _zz_io_B_Valid_44_31;
  reg                 _zz_io_B_Valid_44_32;
  reg                 _zz_io_B_Valid_44_33;
  reg                 _zz_io_B_Valid_44_34;
  reg                 _zz_io_B_Valid_44_35;
  reg                 _zz_io_B_Valid_44_36;
  reg                 _zz_io_B_Valid_44_37;
  reg                 _zz_io_B_Valid_44_38;
  reg                 _zz_io_B_Valid_44_39;
  reg                 _zz_io_B_Valid_44_40;
  reg                 _zz_io_B_Valid_44_41;
  reg                 _zz_io_B_Valid_44_42;
  reg                 _zz_io_B_Valid_44_43;
  reg        [7:0]    _zz_io_MatrixB_45;
  reg        [7:0]    _zz_io_MatrixB_45_1;
  reg        [7:0]    _zz_io_MatrixB_45_2;
  reg        [7:0]    _zz_io_MatrixB_45_3;
  reg        [7:0]    _zz_io_MatrixB_45_4;
  reg        [7:0]    _zz_io_MatrixB_45_5;
  reg        [7:0]    _zz_io_MatrixB_45_6;
  reg        [7:0]    _zz_io_MatrixB_45_7;
  reg        [7:0]    _zz_io_MatrixB_45_8;
  reg        [7:0]    _zz_io_MatrixB_45_9;
  reg        [7:0]    _zz_io_MatrixB_45_10;
  reg        [7:0]    _zz_io_MatrixB_45_11;
  reg        [7:0]    _zz_io_MatrixB_45_12;
  reg        [7:0]    _zz_io_MatrixB_45_13;
  reg        [7:0]    _zz_io_MatrixB_45_14;
  reg        [7:0]    _zz_io_MatrixB_45_15;
  reg        [7:0]    _zz_io_MatrixB_45_16;
  reg        [7:0]    _zz_io_MatrixB_45_17;
  reg        [7:0]    _zz_io_MatrixB_45_18;
  reg        [7:0]    _zz_io_MatrixB_45_19;
  reg        [7:0]    _zz_io_MatrixB_45_20;
  reg        [7:0]    _zz_io_MatrixB_45_21;
  reg        [7:0]    _zz_io_MatrixB_45_22;
  reg        [7:0]    _zz_io_MatrixB_45_23;
  reg        [7:0]    _zz_io_MatrixB_45_24;
  reg        [7:0]    _zz_io_MatrixB_45_25;
  reg        [7:0]    _zz_io_MatrixB_45_26;
  reg        [7:0]    _zz_io_MatrixB_45_27;
  reg        [7:0]    _zz_io_MatrixB_45_28;
  reg        [7:0]    _zz_io_MatrixB_45_29;
  reg        [7:0]    _zz_io_MatrixB_45_30;
  reg        [7:0]    _zz_io_MatrixB_45_31;
  reg        [7:0]    _zz_io_MatrixB_45_32;
  reg        [7:0]    _zz_io_MatrixB_45_33;
  reg        [7:0]    _zz_io_MatrixB_45_34;
  reg        [7:0]    _zz_io_MatrixB_45_35;
  reg        [7:0]    _zz_io_MatrixB_45_36;
  reg        [7:0]    _zz_io_MatrixB_45_37;
  reg        [7:0]    _zz_io_MatrixB_45_38;
  reg        [7:0]    _zz_io_MatrixB_45_39;
  reg        [7:0]    _zz_io_MatrixB_45_40;
  reg        [7:0]    _zz_io_MatrixB_45_41;
  reg        [7:0]    _zz_io_MatrixB_45_42;
  reg        [7:0]    _zz_io_MatrixB_45_43;
  reg        [7:0]    _zz_io_MatrixB_45_44;
  reg                 _zz_io_B_Valid_45;
  reg                 _zz_io_B_Valid_45_1;
  reg                 _zz_io_B_Valid_45_2;
  reg                 _zz_io_B_Valid_45_3;
  reg                 _zz_io_B_Valid_45_4;
  reg                 _zz_io_B_Valid_45_5;
  reg                 _zz_io_B_Valid_45_6;
  reg                 _zz_io_B_Valid_45_7;
  reg                 _zz_io_B_Valid_45_8;
  reg                 _zz_io_B_Valid_45_9;
  reg                 _zz_io_B_Valid_45_10;
  reg                 _zz_io_B_Valid_45_11;
  reg                 _zz_io_B_Valid_45_12;
  reg                 _zz_io_B_Valid_45_13;
  reg                 _zz_io_B_Valid_45_14;
  reg                 _zz_io_B_Valid_45_15;
  reg                 _zz_io_B_Valid_45_16;
  reg                 _zz_io_B_Valid_45_17;
  reg                 _zz_io_B_Valid_45_18;
  reg                 _zz_io_B_Valid_45_19;
  reg                 _zz_io_B_Valid_45_20;
  reg                 _zz_io_B_Valid_45_21;
  reg                 _zz_io_B_Valid_45_22;
  reg                 _zz_io_B_Valid_45_23;
  reg                 _zz_io_B_Valid_45_24;
  reg                 _zz_io_B_Valid_45_25;
  reg                 _zz_io_B_Valid_45_26;
  reg                 _zz_io_B_Valid_45_27;
  reg                 _zz_io_B_Valid_45_28;
  reg                 _zz_io_B_Valid_45_29;
  reg                 _zz_io_B_Valid_45_30;
  reg                 _zz_io_B_Valid_45_31;
  reg                 _zz_io_B_Valid_45_32;
  reg                 _zz_io_B_Valid_45_33;
  reg                 _zz_io_B_Valid_45_34;
  reg                 _zz_io_B_Valid_45_35;
  reg                 _zz_io_B_Valid_45_36;
  reg                 _zz_io_B_Valid_45_37;
  reg                 _zz_io_B_Valid_45_38;
  reg                 _zz_io_B_Valid_45_39;
  reg                 _zz_io_B_Valid_45_40;
  reg                 _zz_io_B_Valid_45_41;
  reg                 _zz_io_B_Valid_45_42;
  reg                 _zz_io_B_Valid_45_43;
  reg                 _zz_io_B_Valid_45_44;
  reg        [7:0]    _zz_io_MatrixB_46;
  reg        [7:0]    _zz_io_MatrixB_46_1;
  reg        [7:0]    _zz_io_MatrixB_46_2;
  reg        [7:0]    _zz_io_MatrixB_46_3;
  reg        [7:0]    _zz_io_MatrixB_46_4;
  reg        [7:0]    _zz_io_MatrixB_46_5;
  reg        [7:0]    _zz_io_MatrixB_46_6;
  reg        [7:0]    _zz_io_MatrixB_46_7;
  reg        [7:0]    _zz_io_MatrixB_46_8;
  reg        [7:0]    _zz_io_MatrixB_46_9;
  reg        [7:0]    _zz_io_MatrixB_46_10;
  reg        [7:0]    _zz_io_MatrixB_46_11;
  reg        [7:0]    _zz_io_MatrixB_46_12;
  reg        [7:0]    _zz_io_MatrixB_46_13;
  reg        [7:0]    _zz_io_MatrixB_46_14;
  reg        [7:0]    _zz_io_MatrixB_46_15;
  reg        [7:0]    _zz_io_MatrixB_46_16;
  reg        [7:0]    _zz_io_MatrixB_46_17;
  reg        [7:0]    _zz_io_MatrixB_46_18;
  reg        [7:0]    _zz_io_MatrixB_46_19;
  reg        [7:0]    _zz_io_MatrixB_46_20;
  reg        [7:0]    _zz_io_MatrixB_46_21;
  reg        [7:0]    _zz_io_MatrixB_46_22;
  reg        [7:0]    _zz_io_MatrixB_46_23;
  reg        [7:0]    _zz_io_MatrixB_46_24;
  reg        [7:0]    _zz_io_MatrixB_46_25;
  reg        [7:0]    _zz_io_MatrixB_46_26;
  reg        [7:0]    _zz_io_MatrixB_46_27;
  reg        [7:0]    _zz_io_MatrixB_46_28;
  reg        [7:0]    _zz_io_MatrixB_46_29;
  reg        [7:0]    _zz_io_MatrixB_46_30;
  reg        [7:0]    _zz_io_MatrixB_46_31;
  reg        [7:0]    _zz_io_MatrixB_46_32;
  reg        [7:0]    _zz_io_MatrixB_46_33;
  reg        [7:0]    _zz_io_MatrixB_46_34;
  reg        [7:0]    _zz_io_MatrixB_46_35;
  reg        [7:0]    _zz_io_MatrixB_46_36;
  reg        [7:0]    _zz_io_MatrixB_46_37;
  reg        [7:0]    _zz_io_MatrixB_46_38;
  reg        [7:0]    _zz_io_MatrixB_46_39;
  reg        [7:0]    _zz_io_MatrixB_46_40;
  reg        [7:0]    _zz_io_MatrixB_46_41;
  reg        [7:0]    _zz_io_MatrixB_46_42;
  reg        [7:0]    _zz_io_MatrixB_46_43;
  reg        [7:0]    _zz_io_MatrixB_46_44;
  reg        [7:0]    _zz_io_MatrixB_46_45;
  reg                 _zz_io_B_Valid_46;
  reg                 _zz_io_B_Valid_46_1;
  reg                 _zz_io_B_Valid_46_2;
  reg                 _zz_io_B_Valid_46_3;
  reg                 _zz_io_B_Valid_46_4;
  reg                 _zz_io_B_Valid_46_5;
  reg                 _zz_io_B_Valid_46_6;
  reg                 _zz_io_B_Valid_46_7;
  reg                 _zz_io_B_Valid_46_8;
  reg                 _zz_io_B_Valid_46_9;
  reg                 _zz_io_B_Valid_46_10;
  reg                 _zz_io_B_Valid_46_11;
  reg                 _zz_io_B_Valid_46_12;
  reg                 _zz_io_B_Valid_46_13;
  reg                 _zz_io_B_Valid_46_14;
  reg                 _zz_io_B_Valid_46_15;
  reg                 _zz_io_B_Valid_46_16;
  reg                 _zz_io_B_Valid_46_17;
  reg                 _zz_io_B_Valid_46_18;
  reg                 _zz_io_B_Valid_46_19;
  reg                 _zz_io_B_Valid_46_20;
  reg                 _zz_io_B_Valid_46_21;
  reg                 _zz_io_B_Valid_46_22;
  reg                 _zz_io_B_Valid_46_23;
  reg                 _zz_io_B_Valid_46_24;
  reg                 _zz_io_B_Valid_46_25;
  reg                 _zz_io_B_Valid_46_26;
  reg                 _zz_io_B_Valid_46_27;
  reg                 _zz_io_B_Valid_46_28;
  reg                 _zz_io_B_Valid_46_29;
  reg                 _zz_io_B_Valid_46_30;
  reg                 _zz_io_B_Valid_46_31;
  reg                 _zz_io_B_Valid_46_32;
  reg                 _zz_io_B_Valid_46_33;
  reg                 _zz_io_B_Valid_46_34;
  reg                 _zz_io_B_Valid_46_35;
  reg                 _zz_io_B_Valid_46_36;
  reg                 _zz_io_B_Valid_46_37;
  reg                 _zz_io_B_Valid_46_38;
  reg                 _zz_io_B_Valid_46_39;
  reg                 _zz_io_B_Valid_46_40;
  reg                 _zz_io_B_Valid_46_41;
  reg                 _zz_io_B_Valid_46_42;
  reg                 _zz_io_B_Valid_46_43;
  reg                 _zz_io_B_Valid_46_44;
  reg                 _zz_io_B_Valid_46_45;
  reg        [7:0]    _zz_io_MatrixB_47;
  reg        [7:0]    _zz_io_MatrixB_47_1;
  reg        [7:0]    _zz_io_MatrixB_47_2;
  reg        [7:0]    _zz_io_MatrixB_47_3;
  reg        [7:0]    _zz_io_MatrixB_47_4;
  reg        [7:0]    _zz_io_MatrixB_47_5;
  reg        [7:0]    _zz_io_MatrixB_47_6;
  reg        [7:0]    _zz_io_MatrixB_47_7;
  reg        [7:0]    _zz_io_MatrixB_47_8;
  reg        [7:0]    _zz_io_MatrixB_47_9;
  reg        [7:0]    _zz_io_MatrixB_47_10;
  reg        [7:0]    _zz_io_MatrixB_47_11;
  reg        [7:0]    _zz_io_MatrixB_47_12;
  reg        [7:0]    _zz_io_MatrixB_47_13;
  reg        [7:0]    _zz_io_MatrixB_47_14;
  reg        [7:0]    _zz_io_MatrixB_47_15;
  reg        [7:0]    _zz_io_MatrixB_47_16;
  reg        [7:0]    _zz_io_MatrixB_47_17;
  reg        [7:0]    _zz_io_MatrixB_47_18;
  reg        [7:0]    _zz_io_MatrixB_47_19;
  reg        [7:0]    _zz_io_MatrixB_47_20;
  reg        [7:0]    _zz_io_MatrixB_47_21;
  reg        [7:0]    _zz_io_MatrixB_47_22;
  reg        [7:0]    _zz_io_MatrixB_47_23;
  reg        [7:0]    _zz_io_MatrixB_47_24;
  reg        [7:0]    _zz_io_MatrixB_47_25;
  reg        [7:0]    _zz_io_MatrixB_47_26;
  reg        [7:0]    _zz_io_MatrixB_47_27;
  reg        [7:0]    _zz_io_MatrixB_47_28;
  reg        [7:0]    _zz_io_MatrixB_47_29;
  reg        [7:0]    _zz_io_MatrixB_47_30;
  reg        [7:0]    _zz_io_MatrixB_47_31;
  reg        [7:0]    _zz_io_MatrixB_47_32;
  reg        [7:0]    _zz_io_MatrixB_47_33;
  reg        [7:0]    _zz_io_MatrixB_47_34;
  reg        [7:0]    _zz_io_MatrixB_47_35;
  reg        [7:0]    _zz_io_MatrixB_47_36;
  reg        [7:0]    _zz_io_MatrixB_47_37;
  reg        [7:0]    _zz_io_MatrixB_47_38;
  reg        [7:0]    _zz_io_MatrixB_47_39;
  reg        [7:0]    _zz_io_MatrixB_47_40;
  reg        [7:0]    _zz_io_MatrixB_47_41;
  reg        [7:0]    _zz_io_MatrixB_47_42;
  reg        [7:0]    _zz_io_MatrixB_47_43;
  reg        [7:0]    _zz_io_MatrixB_47_44;
  reg        [7:0]    _zz_io_MatrixB_47_45;
  reg        [7:0]    _zz_io_MatrixB_47_46;
  reg                 _zz_io_B_Valid_47;
  reg                 _zz_io_B_Valid_47_1;
  reg                 _zz_io_B_Valid_47_2;
  reg                 _zz_io_B_Valid_47_3;
  reg                 _zz_io_B_Valid_47_4;
  reg                 _zz_io_B_Valid_47_5;
  reg                 _zz_io_B_Valid_47_6;
  reg                 _zz_io_B_Valid_47_7;
  reg                 _zz_io_B_Valid_47_8;
  reg                 _zz_io_B_Valid_47_9;
  reg                 _zz_io_B_Valid_47_10;
  reg                 _zz_io_B_Valid_47_11;
  reg                 _zz_io_B_Valid_47_12;
  reg                 _zz_io_B_Valid_47_13;
  reg                 _zz_io_B_Valid_47_14;
  reg                 _zz_io_B_Valid_47_15;
  reg                 _zz_io_B_Valid_47_16;
  reg                 _zz_io_B_Valid_47_17;
  reg                 _zz_io_B_Valid_47_18;
  reg                 _zz_io_B_Valid_47_19;
  reg                 _zz_io_B_Valid_47_20;
  reg                 _zz_io_B_Valid_47_21;
  reg                 _zz_io_B_Valid_47_22;
  reg                 _zz_io_B_Valid_47_23;
  reg                 _zz_io_B_Valid_47_24;
  reg                 _zz_io_B_Valid_47_25;
  reg                 _zz_io_B_Valid_47_26;
  reg                 _zz_io_B_Valid_47_27;
  reg                 _zz_io_B_Valid_47_28;
  reg                 _zz_io_B_Valid_47_29;
  reg                 _zz_io_B_Valid_47_30;
  reg                 _zz_io_B_Valid_47_31;
  reg                 _zz_io_B_Valid_47_32;
  reg                 _zz_io_B_Valid_47_33;
  reg                 _zz_io_B_Valid_47_34;
  reg                 _zz_io_B_Valid_47_35;
  reg                 _zz_io_B_Valid_47_36;
  reg                 _zz_io_B_Valid_47_37;
  reg                 _zz_io_B_Valid_47_38;
  reg                 _zz_io_B_Valid_47_39;
  reg                 _zz_io_B_Valid_47_40;
  reg                 _zz_io_B_Valid_47_41;
  reg                 _zz_io_B_Valid_47_42;
  reg                 _zz_io_B_Valid_47_43;
  reg                 _zz_io_B_Valid_47_44;
  reg                 _zz_io_B_Valid_47_45;
  reg                 _zz_io_B_Valid_47_46;
  reg        [7:0]    _zz_io_MatrixB_48;
  reg        [7:0]    _zz_io_MatrixB_48_1;
  reg        [7:0]    _zz_io_MatrixB_48_2;
  reg        [7:0]    _zz_io_MatrixB_48_3;
  reg        [7:0]    _zz_io_MatrixB_48_4;
  reg        [7:0]    _zz_io_MatrixB_48_5;
  reg        [7:0]    _zz_io_MatrixB_48_6;
  reg        [7:0]    _zz_io_MatrixB_48_7;
  reg        [7:0]    _zz_io_MatrixB_48_8;
  reg        [7:0]    _zz_io_MatrixB_48_9;
  reg        [7:0]    _zz_io_MatrixB_48_10;
  reg        [7:0]    _zz_io_MatrixB_48_11;
  reg        [7:0]    _zz_io_MatrixB_48_12;
  reg        [7:0]    _zz_io_MatrixB_48_13;
  reg        [7:0]    _zz_io_MatrixB_48_14;
  reg        [7:0]    _zz_io_MatrixB_48_15;
  reg        [7:0]    _zz_io_MatrixB_48_16;
  reg        [7:0]    _zz_io_MatrixB_48_17;
  reg        [7:0]    _zz_io_MatrixB_48_18;
  reg        [7:0]    _zz_io_MatrixB_48_19;
  reg        [7:0]    _zz_io_MatrixB_48_20;
  reg        [7:0]    _zz_io_MatrixB_48_21;
  reg        [7:0]    _zz_io_MatrixB_48_22;
  reg        [7:0]    _zz_io_MatrixB_48_23;
  reg        [7:0]    _zz_io_MatrixB_48_24;
  reg        [7:0]    _zz_io_MatrixB_48_25;
  reg        [7:0]    _zz_io_MatrixB_48_26;
  reg        [7:0]    _zz_io_MatrixB_48_27;
  reg        [7:0]    _zz_io_MatrixB_48_28;
  reg        [7:0]    _zz_io_MatrixB_48_29;
  reg        [7:0]    _zz_io_MatrixB_48_30;
  reg        [7:0]    _zz_io_MatrixB_48_31;
  reg        [7:0]    _zz_io_MatrixB_48_32;
  reg        [7:0]    _zz_io_MatrixB_48_33;
  reg        [7:0]    _zz_io_MatrixB_48_34;
  reg        [7:0]    _zz_io_MatrixB_48_35;
  reg        [7:0]    _zz_io_MatrixB_48_36;
  reg        [7:0]    _zz_io_MatrixB_48_37;
  reg        [7:0]    _zz_io_MatrixB_48_38;
  reg        [7:0]    _zz_io_MatrixB_48_39;
  reg        [7:0]    _zz_io_MatrixB_48_40;
  reg        [7:0]    _zz_io_MatrixB_48_41;
  reg        [7:0]    _zz_io_MatrixB_48_42;
  reg        [7:0]    _zz_io_MatrixB_48_43;
  reg        [7:0]    _zz_io_MatrixB_48_44;
  reg        [7:0]    _zz_io_MatrixB_48_45;
  reg        [7:0]    _zz_io_MatrixB_48_46;
  reg        [7:0]    _zz_io_MatrixB_48_47;
  reg                 _zz_io_B_Valid_48;
  reg                 _zz_io_B_Valid_48_1;
  reg                 _zz_io_B_Valid_48_2;
  reg                 _zz_io_B_Valid_48_3;
  reg                 _zz_io_B_Valid_48_4;
  reg                 _zz_io_B_Valid_48_5;
  reg                 _zz_io_B_Valid_48_6;
  reg                 _zz_io_B_Valid_48_7;
  reg                 _zz_io_B_Valid_48_8;
  reg                 _zz_io_B_Valid_48_9;
  reg                 _zz_io_B_Valid_48_10;
  reg                 _zz_io_B_Valid_48_11;
  reg                 _zz_io_B_Valid_48_12;
  reg                 _zz_io_B_Valid_48_13;
  reg                 _zz_io_B_Valid_48_14;
  reg                 _zz_io_B_Valid_48_15;
  reg                 _zz_io_B_Valid_48_16;
  reg                 _zz_io_B_Valid_48_17;
  reg                 _zz_io_B_Valid_48_18;
  reg                 _zz_io_B_Valid_48_19;
  reg                 _zz_io_B_Valid_48_20;
  reg                 _zz_io_B_Valid_48_21;
  reg                 _zz_io_B_Valid_48_22;
  reg                 _zz_io_B_Valid_48_23;
  reg                 _zz_io_B_Valid_48_24;
  reg                 _zz_io_B_Valid_48_25;
  reg                 _zz_io_B_Valid_48_26;
  reg                 _zz_io_B_Valid_48_27;
  reg                 _zz_io_B_Valid_48_28;
  reg                 _zz_io_B_Valid_48_29;
  reg                 _zz_io_B_Valid_48_30;
  reg                 _zz_io_B_Valid_48_31;
  reg                 _zz_io_B_Valid_48_32;
  reg                 _zz_io_B_Valid_48_33;
  reg                 _zz_io_B_Valid_48_34;
  reg                 _zz_io_B_Valid_48_35;
  reg                 _zz_io_B_Valid_48_36;
  reg                 _zz_io_B_Valid_48_37;
  reg                 _zz_io_B_Valid_48_38;
  reg                 _zz_io_B_Valid_48_39;
  reg                 _zz_io_B_Valid_48_40;
  reg                 _zz_io_B_Valid_48_41;
  reg                 _zz_io_B_Valid_48_42;
  reg                 _zz_io_B_Valid_48_43;
  reg                 _zz_io_B_Valid_48_44;
  reg                 _zz_io_B_Valid_48_45;
  reg                 _zz_io_B_Valid_48_46;
  reg                 _zz_io_B_Valid_48_47;
  reg        [7:0]    _zz_io_MatrixB_49;
  reg        [7:0]    _zz_io_MatrixB_49_1;
  reg        [7:0]    _zz_io_MatrixB_49_2;
  reg        [7:0]    _zz_io_MatrixB_49_3;
  reg        [7:0]    _zz_io_MatrixB_49_4;
  reg        [7:0]    _zz_io_MatrixB_49_5;
  reg        [7:0]    _zz_io_MatrixB_49_6;
  reg        [7:0]    _zz_io_MatrixB_49_7;
  reg        [7:0]    _zz_io_MatrixB_49_8;
  reg        [7:0]    _zz_io_MatrixB_49_9;
  reg        [7:0]    _zz_io_MatrixB_49_10;
  reg        [7:0]    _zz_io_MatrixB_49_11;
  reg        [7:0]    _zz_io_MatrixB_49_12;
  reg        [7:0]    _zz_io_MatrixB_49_13;
  reg        [7:0]    _zz_io_MatrixB_49_14;
  reg        [7:0]    _zz_io_MatrixB_49_15;
  reg        [7:0]    _zz_io_MatrixB_49_16;
  reg        [7:0]    _zz_io_MatrixB_49_17;
  reg        [7:0]    _zz_io_MatrixB_49_18;
  reg        [7:0]    _zz_io_MatrixB_49_19;
  reg        [7:0]    _zz_io_MatrixB_49_20;
  reg        [7:0]    _zz_io_MatrixB_49_21;
  reg        [7:0]    _zz_io_MatrixB_49_22;
  reg        [7:0]    _zz_io_MatrixB_49_23;
  reg        [7:0]    _zz_io_MatrixB_49_24;
  reg        [7:0]    _zz_io_MatrixB_49_25;
  reg        [7:0]    _zz_io_MatrixB_49_26;
  reg        [7:0]    _zz_io_MatrixB_49_27;
  reg        [7:0]    _zz_io_MatrixB_49_28;
  reg        [7:0]    _zz_io_MatrixB_49_29;
  reg        [7:0]    _zz_io_MatrixB_49_30;
  reg        [7:0]    _zz_io_MatrixB_49_31;
  reg        [7:0]    _zz_io_MatrixB_49_32;
  reg        [7:0]    _zz_io_MatrixB_49_33;
  reg        [7:0]    _zz_io_MatrixB_49_34;
  reg        [7:0]    _zz_io_MatrixB_49_35;
  reg        [7:0]    _zz_io_MatrixB_49_36;
  reg        [7:0]    _zz_io_MatrixB_49_37;
  reg        [7:0]    _zz_io_MatrixB_49_38;
  reg        [7:0]    _zz_io_MatrixB_49_39;
  reg        [7:0]    _zz_io_MatrixB_49_40;
  reg        [7:0]    _zz_io_MatrixB_49_41;
  reg        [7:0]    _zz_io_MatrixB_49_42;
  reg        [7:0]    _zz_io_MatrixB_49_43;
  reg        [7:0]    _zz_io_MatrixB_49_44;
  reg        [7:0]    _zz_io_MatrixB_49_45;
  reg        [7:0]    _zz_io_MatrixB_49_46;
  reg        [7:0]    _zz_io_MatrixB_49_47;
  reg        [7:0]    _zz_io_MatrixB_49_48;
  reg                 _zz_io_B_Valid_49;
  reg                 _zz_io_B_Valid_49_1;
  reg                 _zz_io_B_Valid_49_2;
  reg                 _zz_io_B_Valid_49_3;
  reg                 _zz_io_B_Valid_49_4;
  reg                 _zz_io_B_Valid_49_5;
  reg                 _zz_io_B_Valid_49_6;
  reg                 _zz_io_B_Valid_49_7;
  reg                 _zz_io_B_Valid_49_8;
  reg                 _zz_io_B_Valid_49_9;
  reg                 _zz_io_B_Valid_49_10;
  reg                 _zz_io_B_Valid_49_11;
  reg                 _zz_io_B_Valid_49_12;
  reg                 _zz_io_B_Valid_49_13;
  reg                 _zz_io_B_Valid_49_14;
  reg                 _zz_io_B_Valid_49_15;
  reg                 _zz_io_B_Valid_49_16;
  reg                 _zz_io_B_Valid_49_17;
  reg                 _zz_io_B_Valid_49_18;
  reg                 _zz_io_B_Valid_49_19;
  reg                 _zz_io_B_Valid_49_20;
  reg                 _zz_io_B_Valid_49_21;
  reg                 _zz_io_B_Valid_49_22;
  reg                 _zz_io_B_Valid_49_23;
  reg                 _zz_io_B_Valid_49_24;
  reg                 _zz_io_B_Valid_49_25;
  reg                 _zz_io_B_Valid_49_26;
  reg                 _zz_io_B_Valid_49_27;
  reg                 _zz_io_B_Valid_49_28;
  reg                 _zz_io_B_Valid_49_29;
  reg                 _zz_io_B_Valid_49_30;
  reg                 _zz_io_B_Valid_49_31;
  reg                 _zz_io_B_Valid_49_32;
  reg                 _zz_io_B_Valid_49_33;
  reg                 _zz_io_B_Valid_49_34;
  reg                 _zz_io_B_Valid_49_35;
  reg                 _zz_io_B_Valid_49_36;
  reg                 _zz_io_B_Valid_49_37;
  reg                 _zz_io_B_Valid_49_38;
  reg                 _zz_io_B_Valid_49_39;
  reg                 _zz_io_B_Valid_49_40;
  reg                 _zz_io_B_Valid_49_41;
  reg                 _zz_io_B_Valid_49_42;
  reg                 _zz_io_B_Valid_49_43;
  reg                 _zz_io_B_Valid_49_44;
  reg                 _zz_io_B_Valid_49_45;
  reg                 _zz_io_B_Valid_49_46;
  reg                 _zz_io_B_Valid_49_47;
  reg                 _zz_io_B_Valid_49_48;
  reg        [7:0]    _zz_io_MatrixB_50;
  reg        [7:0]    _zz_io_MatrixB_50_1;
  reg        [7:0]    _zz_io_MatrixB_50_2;
  reg        [7:0]    _zz_io_MatrixB_50_3;
  reg        [7:0]    _zz_io_MatrixB_50_4;
  reg        [7:0]    _zz_io_MatrixB_50_5;
  reg        [7:0]    _zz_io_MatrixB_50_6;
  reg        [7:0]    _zz_io_MatrixB_50_7;
  reg        [7:0]    _zz_io_MatrixB_50_8;
  reg        [7:0]    _zz_io_MatrixB_50_9;
  reg        [7:0]    _zz_io_MatrixB_50_10;
  reg        [7:0]    _zz_io_MatrixB_50_11;
  reg        [7:0]    _zz_io_MatrixB_50_12;
  reg        [7:0]    _zz_io_MatrixB_50_13;
  reg        [7:0]    _zz_io_MatrixB_50_14;
  reg        [7:0]    _zz_io_MatrixB_50_15;
  reg        [7:0]    _zz_io_MatrixB_50_16;
  reg        [7:0]    _zz_io_MatrixB_50_17;
  reg        [7:0]    _zz_io_MatrixB_50_18;
  reg        [7:0]    _zz_io_MatrixB_50_19;
  reg        [7:0]    _zz_io_MatrixB_50_20;
  reg        [7:0]    _zz_io_MatrixB_50_21;
  reg        [7:0]    _zz_io_MatrixB_50_22;
  reg        [7:0]    _zz_io_MatrixB_50_23;
  reg        [7:0]    _zz_io_MatrixB_50_24;
  reg        [7:0]    _zz_io_MatrixB_50_25;
  reg        [7:0]    _zz_io_MatrixB_50_26;
  reg        [7:0]    _zz_io_MatrixB_50_27;
  reg        [7:0]    _zz_io_MatrixB_50_28;
  reg        [7:0]    _zz_io_MatrixB_50_29;
  reg        [7:0]    _zz_io_MatrixB_50_30;
  reg        [7:0]    _zz_io_MatrixB_50_31;
  reg        [7:0]    _zz_io_MatrixB_50_32;
  reg        [7:0]    _zz_io_MatrixB_50_33;
  reg        [7:0]    _zz_io_MatrixB_50_34;
  reg        [7:0]    _zz_io_MatrixB_50_35;
  reg        [7:0]    _zz_io_MatrixB_50_36;
  reg        [7:0]    _zz_io_MatrixB_50_37;
  reg        [7:0]    _zz_io_MatrixB_50_38;
  reg        [7:0]    _zz_io_MatrixB_50_39;
  reg        [7:0]    _zz_io_MatrixB_50_40;
  reg        [7:0]    _zz_io_MatrixB_50_41;
  reg        [7:0]    _zz_io_MatrixB_50_42;
  reg        [7:0]    _zz_io_MatrixB_50_43;
  reg        [7:0]    _zz_io_MatrixB_50_44;
  reg        [7:0]    _zz_io_MatrixB_50_45;
  reg        [7:0]    _zz_io_MatrixB_50_46;
  reg        [7:0]    _zz_io_MatrixB_50_47;
  reg        [7:0]    _zz_io_MatrixB_50_48;
  reg        [7:0]    _zz_io_MatrixB_50_49;
  reg                 _zz_io_B_Valid_50;
  reg                 _zz_io_B_Valid_50_1;
  reg                 _zz_io_B_Valid_50_2;
  reg                 _zz_io_B_Valid_50_3;
  reg                 _zz_io_B_Valid_50_4;
  reg                 _zz_io_B_Valid_50_5;
  reg                 _zz_io_B_Valid_50_6;
  reg                 _zz_io_B_Valid_50_7;
  reg                 _zz_io_B_Valid_50_8;
  reg                 _zz_io_B_Valid_50_9;
  reg                 _zz_io_B_Valid_50_10;
  reg                 _zz_io_B_Valid_50_11;
  reg                 _zz_io_B_Valid_50_12;
  reg                 _zz_io_B_Valid_50_13;
  reg                 _zz_io_B_Valid_50_14;
  reg                 _zz_io_B_Valid_50_15;
  reg                 _zz_io_B_Valid_50_16;
  reg                 _zz_io_B_Valid_50_17;
  reg                 _zz_io_B_Valid_50_18;
  reg                 _zz_io_B_Valid_50_19;
  reg                 _zz_io_B_Valid_50_20;
  reg                 _zz_io_B_Valid_50_21;
  reg                 _zz_io_B_Valid_50_22;
  reg                 _zz_io_B_Valid_50_23;
  reg                 _zz_io_B_Valid_50_24;
  reg                 _zz_io_B_Valid_50_25;
  reg                 _zz_io_B_Valid_50_26;
  reg                 _zz_io_B_Valid_50_27;
  reg                 _zz_io_B_Valid_50_28;
  reg                 _zz_io_B_Valid_50_29;
  reg                 _zz_io_B_Valid_50_30;
  reg                 _zz_io_B_Valid_50_31;
  reg                 _zz_io_B_Valid_50_32;
  reg                 _zz_io_B_Valid_50_33;
  reg                 _zz_io_B_Valid_50_34;
  reg                 _zz_io_B_Valid_50_35;
  reg                 _zz_io_B_Valid_50_36;
  reg                 _zz_io_B_Valid_50_37;
  reg                 _zz_io_B_Valid_50_38;
  reg                 _zz_io_B_Valid_50_39;
  reg                 _zz_io_B_Valid_50_40;
  reg                 _zz_io_B_Valid_50_41;
  reg                 _zz_io_B_Valid_50_42;
  reg                 _zz_io_B_Valid_50_43;
  reg                 _zz_io_B_Valid_50_44;
  reg                 _zz_io_B_Valid_50_45;
  reg                 _zz_io_B_Valid_50_46;
  reg                 _zz_io_B_Valid_50_47;
  reg                 _zz_io_B_Valid_50_48;
  reg                 _zz_io_B_Valid_50_49;
  reg        [7:0]    _zz_io_MatrixB_51;
  reg        [7:0]    _zz_io_MatrixB_51_1;
  reg        [7:0]    _zz_io_MatrixB_51_2;
  reg        [7:0]    _zz_io_MatrixB_51_3;
  reg        [7:0]    _zz_io_MatrixB_51_4;
  reg        [7:0]    _zz_io_MatrixB_51_5;
  reg        [7:0]    _zz_io_MatrixB_51_6;
  reg        [7:0]    _zz_io_MatrixB_51_7;
  reg        [7:0]    _zz_io_MatrixB_51_8;
  reg        [7:0]    _zz_io_MatrixB_51_9;
  reg        [7:0]    _zz_io_MatrixB_51_10;
  reg        [7:0]    _zz_io_MatrixB_51_11;
  reg        [7:0]    _zz_io_MatrixB_51_12;
  reg        [7:0]    _zz_io_MatrixB_51_13;
  reg        [7:0]    _zz_io_MatrixB_51_14;
  reg        [7:0]    _zz_io_MatrixB_51_15;
  reg        [7:0]    _zz_io_MatrixB_51_16;
  reg        [7:0]    _zz_io_MatrixB_51_17;
  reg        [7:0]    _zz_io_MatrixB_51_18;
  reg        [7:0]    _zz_io_MatrixB_51_19;
  reg        [7:0]    _zz_io_MatrixB_51_20;
  reg        [7:0]    _zz_io_MatrixB_51_21;
  reg        [7:0]    _zz_io_MatrixB_51_22;
  reg        [7:0]    _zz_io_MatrixB_51_23;
  reg        [7:0]    _zz_io_MatrixB_51_24;
  reg        [7:0]    _zz_io_MatrixB_51_25;
  reg        [7:0]    _zz_io_MatrixB_51_26;
  reg        [7:0]    _zz_io_MatrixB_51_27;
  reg        [7:0]    _zz_io_MatrixB_51_28;
  reg        [7:0]    _zz_io_MatrixB_51_29;
  reg        [7:0]    _zz_io_MatrixB_51_30;
  reg        [7:0]    _zz_io_MatrixB_51_31;
  reg        [7:0]    _zz_io_MatrixB_51_32;
  reg        [7:0]    _zz_io_MatrixB_51_33;
  reg        [7:0]    _zz_io_MatrixB_51_34;
  reg        [7:0]    _zz_io_MatrixB_51_35;
  reg        [7:0]    _zz_io_MatrixB_51_36;
  reg        [7:0]    _zz_io_MatrixB_51_37;
  reg        [7:0]    _zz_io_MatrixB_51_38;
  reg        [7:0]    _zz_io_MatrixB_51_39;
  reg        [7:0]    _zz_io_MatrixB_51_40;
  reg        [7:0]    _zz_io_MatrixB_51_41;
  reg        [7:0]    _zz_io_MatrixB_51_42;
  reg        [7:0]    _zz_io_MatrixB_51_43;
  reg        [7:0]    _zz_io_MatrixB_51_44;
  reg        [7:0]    _zz_io_MatrixB_51_45;
  reg        [7:0]    _zz_io_MatrixB_51_46;
  reg        [7:0]    _zz_io_MatrixB_51_47;
  reg        [7:0]    _zz_io_MatrixB_51_48;
  reg        [7:0]    _zz_io_MatrixB_51_49;
  reg        [7:0]    _zz_io_MatrixB_51_50;
  reg                 _zz_io_B_Valid_51;
  reg                 _zz_io_B_Valid_51_1;
  reg                 _zz_io_B_Valid_51_2;
  reg                 _zz_io_B_Valid_51_3;
  reg                 _zz_io_B_Valid_51_4;
  reg                 _zz_io_B_Valid_51_5;
  reg                 _zz_io_B_Valid_51_6;
  reg                 _zz_io_B_Valid_51_7;
  reg                 _zz_io_B_Valid_51_8;
  reg                 _zz_io_B_Valid_51_9;
  reg                 _zz_io_B_Valid_51_10;
  reg                 _zz_io_B_Valid_51_11;
  reg                 _zz_io_B_Valid_51_12;
  reg                 _zz_io_B_Valid_51_13;
  reg                 _zz_io_B_Valid_51_14;
  reg                 _zz_io_B_Valid_51_15;
  reg                 _zz_io_B_Valid_51_16;
  reg                 _zz_io_B_Valid_51_17;
  reg                 _zz_io_B_Valid_51_18;
  reg                 _zz_io_B_Valid_51_19;
  reg                 _zz_io_B_Valid_51_20;
  reg                 _zz_io_B_Valid_51_21;
  reg                 _zz_io_B_Valid_51_22;
  reg                 _zz_io_B_Valid_51_23;
  reg                 _zz_io_B_Valid_51_24;
  reg                 _zz_io_B_Valid_51_25;
  reg                 _zz_io_B_Valid_51_26;
  reg                 _zz_io_B_Valid_51_27;
  reg                 _zz_io_B_Valid_51_28;
  reg                 _zz_io_B_Valid_51_29;
  reg                 _zz_io_B_Valid_51_30;
  reg                 _zz_io_B_Valid_51_31;
  reg                 _zz_io_B_Valid_51_32;
  reg                 _zz_io_B_Valid_51_33;
  reg                 _zz_io_B_Valid_51_34;
  reg                 _zz_io_B_Valid_51_35;
  reg                 _zz_io_B_Valid_51_36;
  reg                 _zz_io_B_Valid_51_37;
  reg                 _zz_io_B_Valid_51_38;
  reg                 _zz_io_B_Valid_51_39;
  reg                 _zz_io_B_Valid_51_40;
  reg                 _zz_io_B_Valid_51_41;
  reg                 _zz_io_B_Valid_51_42;
  reg                 _zz_io_B_Valid_51_43;
  reg                 _zz_io_B_Valid_51_44;
  reg                 _zz_io_B_Valid_51_45;
  reg                 _zz_io_B_Valid_51_46;
  reg                 _zz_io_B_Valid_51_47;
  reg                 _zz_io_B_Valid_51_48;
  reg                 _zz_io_B_Valid_51_49;
  reg                 _zz_io_B_Valid_51_50;
  reg        [7:0]    _zz_io_MatrixB_52;
  reg        [7:0]    _zz_io_MatrixB_52_1;
  reg        [7:0]    _zz_io_MatrixB_52_2;
  reg        [7:0]    _zz_io_MatrixB_52_3;
  reg        [7:0]    _zz_io_MatrixB_52_4;
  reg        [7:0]    _zz_io_MatrixB_52_5;
  reg        [7:0]    _zz_io_MatrixB_52_6;
  reg        [7:0]    _zz_io_MatrixB_52_7;
  reg        [7:0]    _zz_io_MatrixB_52_8;
  reg        [7:0]    _zz_io_MatrixB_52_9;
  reg        [7:0]    _zz_io_MatrixB_52_10;
  reg        [7:0]    _zz_io_MatrixB_52_11;
  reg        [7:0]    _zz_io_MatrixB_52_12;
  reg        [7:0]    _zz_io_MatrixB_52_13;
  reg        [7:0]    _zz_io_MatrixB_52_14;
  reg        [7:0]    _zz_io_MatrixB_52_15;
  reg        [7:0]    _zz_io_MatrixB_52_16;
  reg        [7:0]    _zz_io_MatrixB_52_17;
  reg        [7:0]    _zz_io_MatrixB_52_18;
  reg        [7:0]    _zz_io_MatrixB_52_19;
  reg        [7:0]    _zz_io_MatrixB_52_20;
  reg        [7:0]    _zz_io_MatrixB_52_21;
  reg        [7:0]    _zz_io_MatrixB_52_22;
  reg        [7:0]    _zz_io_MatrixB_52_23;
  reg        [7:0]    _zz_io_MatrixB_52_24;
  reg        [7:0]    _zz_io_MatrixB_52_25;
  reg        [7:0]    _zz_io_MatrixB_52_26;
  reg        [7:0]    _zz_io_MatrixB_52_27;
  reg        [7:0]    _zz_io_MatrixB_52_28;
  reg        [7:0]    _zz_io_MatrixB_52_29;
  reg        [7:0]    _zz_io_MatrixB_52_30;
  reg        [7:0]    _zz_io_MatrixB_52_31;
  reg        [7:0]    _zz_io_MatrixB_52_32;
  reg        [7:0]    _zz_io_MatrixB_52_33;
  reg        [7:0]    _zz_io_MatrixB_52_34;
  reg        [7:0]    _zz_io_MatrixB_52_35;
  reg        [7:0]    _zz_io_MatrixB_52_36;
  reg        [7:0]    _zz_io_MatrixB_52_37;
  reg        [7:0]    _zz_io_MatrixB_52_38;
  reg        [7:0]    _zz_io_MatrixB_52_39;
  reg        [7:0]    _zz_io_MatrixB_52_40;
  reg        [7:0]    _zz_io_MatrixB_52_41;
  reg        [7:0]    _zz_io_MatrixB_52_42;
  reg        [7:0]    _zz_io_MatrixB_52_43;
  reg        [7:0]    _zz_io_MatrixB_52_44;
  reg        [7:0]    _zz_io_MatrixB_52_45;
  reg        [7:0]    _zz_io_MatrixB_52_46;
  reg        [7:0]    _zz_io_MatrixB_52_47;
  reg        [7:0]    _zz_io_MatrixB_52_48;
  reg        [7:0]    _zz_io_MatrixB_52_49;
  reg        [7:0]    _zz_io_MatrixB_52_50;
  reg        [7:0]    _zz_io_MatrixB_52_51;
  reg                 _zz_io_B_Valid_52;
  reg                 _zz_io_B_Valid_52_1;
  reg                 _zz_io_B_Valid_52_2;
  reg                 _zz_io_B_Valid_52_3;
  reg                 _zz_io_B_Valid_52_4;
  reg                 _zz_io_B_Valid_52_5;
  reg                 _zz_io_B_Valid_52_6;
  reg                 _zz_io_B_Valid_52_7;
  reg                 _zz_io_B_Valid_52_8;
  reg                 _zz_io_B_Valid_52_9;
  reg                 _zz_io_B_Valid_52_10;
  reg                 _zz_io_B_Valid_52_11;
  reg                 _zz_io_B_Valid_52_12;
  reg                 _zz_io_B_Valid_52_13;
  reg                 _zz_io_B_Valid_52_14;
  reg                 _zz_io_B_Valid_52_15;
  reg                 _zz_io_B_Valid_52_16;
  reg                 _zz_io_B_Valid_52_17;
  reg                 _zz_io_B_Valid_52_18;
  reg                 _zz_io_B_Valid_52_19;
  reg                 _zz_io_B_Valid_52_20;
  reg                 _zz_io_B_Valid_52_21;
  reg                 _zz_io_B_Valid_52_22;
  reg                 _zz_io_B_Valid_52_23;
  reg                 _zz_io_B_Valid_52_24;
  reg                 _zz_io_B_Valid_52_25;
  reg                 _zz_io_B_Valid_52_26;
  reg                 _zz_io_B_Valid_52_27;
  reg                 _zz_io_B_Valid_52_28;
  reg                 _zz_io_B_Valid_52_29;
  reg                 _zz_io_B_Valid_52_30;
  reg                 _zz_io_B_Valid_52_31;
  reg                 _zz_io_B_Valid_52_32;
  reg                 _zz_io_B_Valid_52_33;
  reg                 _zz_io_B_Valid_52_34;
  reg                 _zz_io_B_Valid_52_35;
  reg                 _zz_io_B_Valid_52_36;
  reg                 _zz_io_B_Valid_52_37;
  reg                 _zz_io_B_Valid_52_38;
  reg                 _zz_io_B_Valid_52_39;
  reg                 _zz_io_B_Valid_52_40;
  reg                 _zz_io_B_Valid_52_41;
  reg                 _zz_io_B_Valid_52_42;
  reg                 _zz_io_B_Valid_52_43;
  reg                 _zz_io_B_Valid_52_44;
  reg                 _zz_io_B_Valid_52_45;
  reg                 _zz_io_B_Valid_52_46;
  reg                 _zz_io_B_Valid_52_47;
  reg                 _zz_io_B_Valid_52_48;
  reg                 _zz_io_B_Valid_52_49;
  reg                 _zz_io_B_Valid_52_50;
  reg                 _zz_io_B_Valid_52_51;
  reg        [7:0]    _zz_io_MatrixB_53;
  reg        [7:0]    _zz_io_MatrixB_53_1;
  reg        [7:0]    _zz_io_MatrixB_53_2;
  reg        [7:0]    _zz_io_MatrixB_53_3;
  reg        [7:0]    _zz_io_MatrixB_53_4;
  reg        [7:0]    _zz_io_MatrixB_53_5;
  reg        [7:0]    _zz_io_MatrixB_53_6;
  reg        [7:0]    _zz_io_MatrixB_53_7;
  reg        [7:0]    _zz_io_MatrixB_53_8;
  reg        [7:0]    _zz_io_MatrixB_53_9;
  reg        [7:0]    _zz_io_MatrixB_53_10;
  reg        [7:0]    _zz_io_MatrixB_53_11;
  reg        [7:0]    _zz_io_MatrixB_53_12;
  reg        [7:0]    _zz_io_MatrixB_53_13;
  reg        [7:0]    _zz_io_MatrixB_53_14;
  reg        [7:0]    _zz_io_MatrixB_53_15;
  reg        [7:0]    _zz_io_MatrixB_53_16;
  reg        [7:0]    _zz_io_MatrixB_53_17;
  reg        [7:0]    _zz_io_MatrixB_53_18;
  reg        [7:0]    _zz_io_MatrixB_53_19;
  reg        [7:0]    _zz_io_MatrixB_53_20;
  reg        [7:0]    _zz_io_MatrixB_53_21;
  reg        [7:0]    _zz_io_MatrixB_53_22;
  reg        [7:0]    _zz_io_MatrixB_53_23;
  reg        [7:0]    _zz_io_MatrixB_53_24;
  reg        [7:0]    _zz_io_MatrixB_53_25;
  reg        [7:0]    _zz_io_MatrixB_53_26;
  reg        [7:0]    _zz_io_MatrixB_53_27;
  reg        [7:0]    _zz_io_MatrixB_53_28;
  reg        [7:0]    _zz_io_MatrixB_53_29;
  reg        [7:0]    _zz_io_MatrixB_53_30;
  reg        [7:0]    _zz_io_MatrixB_53_31;
  reg        [7:0]    _zz_io_MatrixB_53_32;
  reg        [7:0]    _zz_io_MatrixB_53_33;
  reg        [7:0]    _zz_io_MatrixB_53_34;
  reg        [7:0]    _zz_io_MatrixB_53_35;
  reg        [7:0]    _zz_io_MatrixB_53_36;
  reg        [7:0]    _zz_io_MatrixB_53_37;
  reg        [7:0]    _zz_io_MatrixB_53_38;
  reg        [7:0]    _zz_io_MatrixB_53_39;
  reg        [7:0]    _zz_io_MatrixB_53_40;
  reg        [7:0]    _zz_io_MatrixB_53_41;
  reg        [7:0]    _zz_io_MatrixB_53_42;
  reg        [7:0]    _zz_io_MatrixB_53_43;
  reg        [7:0]    _zz_io_MatrixB_53_44;
  reg        [7:0]    _zz_io_MatrixB_53_45;
  reg        [7:0]    _zz_io_MatrixB_53_46;
  reg        [7:0]    _zz_io_MatrixB_53_47;
  reg        [7:0]    _zz_io_MatrixB_53_48;
  reg        [7:0]    _zz_io_MatrixB_53_49;
  reg        [7:0]    _zz_io_MatrixB_53_50;
  reg        [7:0]    _zz_io_MatrixB_53_51;
  reg        [7:0]    _zz_io_MatrixB_53_52;
  reg                 _zz_io_B_Valid_53;
  reg                 _zz_io_B_Valid_53_1;
  reg                 _zz_io_B_Valid_53_2;
  reg                 _zz_io_B_Valid_53_3;
  reg                 _zz_io_B_Valid_53_4;
  reg                 _zz_io_B_Valid_53_5;
  reg                 _zz_io_B_Valid_53_6;
  reg                 _zz_io_B_Valid_53_7;
  reg                 _zz_io_B_Valid_53_8;
  reg                 _zz_io_B_Valid_53_9;
  reg                 _zz_io_B_Valid_53_10;
  reg                 _zz_io_B_Valid_53_11;
  reg                 _zz_io_B_Valid_53_12;
  reg                 _zz_io_B_Valid_53_13;
  reg                 _zz_io_B_Valid_53_14;
  reg                 _zz_io_B_Valid_53_15;
  reg                 _zz_io_B_Valid_53_16;
  reg                 _zz_io_B_Valid_53_17;
  reg                 _zz_io_B_Valid_53_18;
  reg                 _zz_io_B_Valid_53_19;
  reg                 _zz_io_B_Valid_53_20;
  reg                 _zz_io_B_Valid_53_21;
  reg                 _zz_io_B_Valid_53_22;
  reg                 _zz_io_B_Valid_53_23;
  reg                 _zz_io_B_Valid_53_24;
  reg                 _zz_io_B_Valid_53_25;
  reg                 _zz_io_B_Valid_53_26;
  reg                 _zz_io_B_Valid_53_27;
  reg                 _zz_io_B_Valid_53_28;
  reg                 _zz_io_B_Valid_53_29;
  reg                 _zz_io_B_Valid_53_30;
  reg                 _zz_io_B_Valid_53_31;
  reg                 _zz_io_B_Valid_53_32;
  reg                 _zz_io_B_Valid_53_33;
  reg                 _zz_io_B_Valid_53_34;
  reg                 _zz_io_B_Valid_53_35;
  reg                 _zz_io_B_Valid_53_36;
  reg                 _zz_io_B_Valid_53_37;
  reg                 _zz_io_B_Valid_53_38;
  reg                 _zz_io_B_Valid_53_39;
  reg                 _zz_io_B_Valid_53_40;
  reg                 _zz_io_B_Valid_53_41;
  reg                 _zz_io_B_Valid_53_42;
  reg                 _zz_io_B_Valid_53_43;
  reg                 _zz_io_B_Valid_53_44;
  reg                 _zz_io_B_Valid_53_45;
  reg                 _zz_io_B_Valid_53_46;
  reg                 _zz_io_B_Valid_53_47;
  reg                 _zz_io_B_Valid_53_48;
  reg                 _zz_io_B_Valid_53_49;
  reg                 _zz_io_B_Valid_53_50;
  reg                 _zz_io_B_Valid_53_51;
  reg                 _zz_io_B_Valid_53_52;
  reg        [7:0]    _zz_io_MatrixB_54;
  reg        [7:0]    _zz_io_MatrixB_54_1;
  reg        [7:0]    _zz_io_MatrixB_54_2;
  reg        [7:0]    _zz_io_MatrixB_54_3;
  reg        [7:0]    _zz_io_MatrixB_54_4;
  reg        [7:0]    _zz_io_MatrixB_54_5;
  reg        [7:0]    _zz_io_MatrixB_54_6;
  reg        [7:0]    _zz_io_MatrixB_54_7;
  reg        [7:0]    _zz_io_MatrixB_54_8;
  reg        [7:0]    _zz_io_MatrixB_54_9;
  reg        [7:0]    _zz_io_MatrixB_54_10;
  reg        [7:0]    _zz_io_MatrixB_54_11;
  reg        [7:0]    _zz_io_MatrixB_54_12;
  reg        [7:0]    _zz_io_MatrixB_54_13;
  reg        [7:0]    _zz_io_MatrixB_54_14;
  reg        [7:0]    _zz_io_MatrixB_54_15;
  reg        [7:0]    _zz_io_MatrixB_54_16;
  reg        [7:0]    _zz_io_MatrixB_54_17;
  reg        [7:0]    _zz_io_MatrixB_54_18;
  reg        [7:0]    _zz_io_MatrixB_54_19;
  reg        [7:0]    _zz_io_MatrixB_54_20;
  reg        [7:0]    _zz_io_MatrixB_54_21;
  reg        [7:0]    _zz_io_MatrixB_54_22;
  reg        [7:0]    _zz_io_MatrixB_54_23;
  reg        [7:0]    _zz_io_MatrixB_54_24;
  reg        [7:0]    _zz_io_MatrixB_54_25;
  reg        [7:0]    _zz_io_MatrixB_54_26;
  reg        [7:0]    _zz_io_MatrixB_54_27;
  reg        [7:0]    _zz_io_MatrixB_54_28;
  reg        [7:0]    _zz_io_MatrixB_54_29;
  reg        [7:0]    _zz_io_MatrixB_54_30;
  reg        [7:0]    _zz_io_MatrixB_54_31;
  reg        [7:0]    _zz_io_MatrixB_54_32;
  reg        [7:0]    _zz_io_MatrixB_54_33;
  reg        [7:0]    _zz_io_MatrixB_54_34;
  reg        [7:0]    _zz_io_MatrixB_54_35;
  reg        [7:0]    _zz_io_MatrixB_54_36;
  reg        [7:0]    _zz_io_MatrixB_54_37;
  reg        [7:0]    _zz_io_MatrixB_54_38;
  reg        [7:0]    _zz_io_MatrixB_54_39;
  reg        [7:0]    _zz_io_MatrixB_54_40;
  reg        [7:0]    _zz_io_MatrixB_54_41;
  reg        [7:0]    _zz_io_MatrixB_54_42;
  reg        [7:0]    _zz_io_MatrixB_54_43;
  reg        [7:0]    _zz_io_MatrixB_54_44;
  reg        [7:0]    _zz_io_MatrixB_54_45;
  reg        [7:0]    _zz_io_MatrixB_54_46;
  reg        [7:0]    _zz_io_MatrixB_54_47;
  reg        [7:0]    _zz_io_MatrixB_54_48;
  reg        [7:0]    _zz_io_MatrixB_54_49;
  reg        [7:0]    _zz_io_MatrixB_54_50;
  reg        [7:0]    _zz_io_MatrixB_54_51;
  reg        [7:0]    _zz_io_MatrixB_54_52;
  reg        [7:0]    _zz_io_MatrixB_54_53;
  reg                 _zz_io_B_Valid_54;
  reg                 _zz_io_B_Valid_54_1;
  reg                 _zz_io_B_Valid_54_2;
  reg                 _zz_io_B_Valid_54_3;
  reg                 _zz_io_B_Valid_54_4;
  reg                 _zz_io_B_Valid_54_5;
  reg                 _zz_io_B_Valid_54_6;
  reg                 _zz_io_B_Valid_54_7;
  reg                 _zz_io_B_Valid_54_8;
  reg                 _zz_io_B_Valid_54_9;
  reg                 _zz_io_B_Valid_54_10;
  reg                 _zz_io_B_Valid_54_11;
  reg                 _zz_io_B_Valid_54_12;
  reg                 _zz_io_B_Valid_54_13;
  reg                 _zz_io_B_Valid_54_14;
  reg                 _zz_io_B_Valid_54_15;
  reg                 _zz_io_B_Valid_54_16;
  reg                 _zz_io_B_Valid_54_17;
  reg                 _zz_io_B_Valid_54_18;
  reg                 _zz_io_B_Valid_54_19;
  reg                 _zz_io_B_Valid_54_20;
  reg                 _zz_io_B_Valid_54_21;
  reg                 _zz_io_B_Valid_54_22;
  reg                 _zz_io_B_Valid_54_23;
  reg                 _zz_io_B_Valid_54_24;
  reg                 _zz_io_B_Valid_54_25;
  reg                 _zz_io_B_Valid_54_26;
  reg                 _zz_io_B_Valid_54_27;
  reg                 _zz_io_B_Valid_54_28;
  reg                 _zz_io_B_Valid_54_29;
  reg                 _zz_io_B_Valid_54_30;
  reg                 _zz_io_B_Valid_54_31;
  reg                 _zz_io_B_Valid_54_32;
  reg                 _zz_io_B_Valid_54_33;
  reg                 _zz_io_B_Valid_54_34;
  reg                 _zz_io_B_Valid_54_35;
  reg                 _zz_io_B_Valid_54_36;
  reg                 _zz_io_B_Valid_54_37;
  reg                 _zz_io_B_Valid_54_38;
  reg                 _zz_io_B_Valid_54_39;
  reg                 _zz_io_B_Valid_54_40;
  reg                 _zz_io_B_Valid_54_41;
  reg                 _zz_io_B_Valid_54_42;
  reg                 _zz_io_B_Valid_54_43;
  reg                 _zz_io_B_Valid_54_44;
  reg                 _zz_io_B_Valid_54_45;
  reg                 _zz_io_B_Valid_54_46;
  reg                 _zz_io_B_Valid_54_47;
  reg                 _zz_io_B_Valid_54_48;
  reg                 _zz_io_B_Valid_54_49;
  reg                 _zz_io_B_Valid_54_50;
  reg                 _zz_io_B_Valid_54_51;
  reg                 _zz_io_B_Valid_54_52;
  reg                 _zz_io_B_Valid_54_53;
  reg        [7:0]    _zz_io_MatrixB_55;
  reg        [7:0]    _zz_io_MatrixB_55_1;
  reg        [7:0]    _zz_io_MatrixB_55_2;
  reg        [7:0]    _zz_io_MatrixB_55_3;
  reg        [7:0]    _zz_io_MatrixB_55_4;
  reg        [7:0]    _zz_io_MatrixB_55_5;
  reg        [7:0]    _zz_io_MatrixB_55_6;
  reg        [7:0]    _zz_io_MatrixB_55_7;
  reg        [7:0]    _zz_io_MatrixB_55_8;
  reg        [7:0]    _zz_io_MatrixB_55_9;
  reg        [7:0]    _zz_io_MatrixB_55_10;
  reg        [7:0]    _zz_io_MatrixB_55_11;
  reg        [7:0]    _zz_io_MatrixB_55_12;
  reg        [7:0]    _zz_io_MatrixB_55_13;
  reg        [7:0]    _zz_io_MatrixB_55_14;
  reg        [7:0]    _zz_io_MatrixB_55_15;
  reg        [7:0]    _zz_io_MatrixB_55_16;
  reg        [7:0]    _zz_io_MatrixB_55_17;
  reg        [7:0]    _zz_io_MatrixB_55_18;
  reg        [7:0]    _zz_io_MatrixB_55_19;
  reg        [7:0]    _zz_io_MatrixB_55_20;
  reg        [7:0]    _zz_io_MatrixB_55_21;
  reg        [7:0]    _zz_io_MatrixB_55_22;
  reg        [7:0]    _zz_io_MatrixB_55_23;
  reg        [7:0]    _zz_io_MatrixB_55_24;
  reg        [7:0]    _zz_io_MatrixB_55_25;
  reg        [7:0]    _zz_io_MatrixB_55_26;
  reg        [7:0]    _zz_io_MatrixB_55_27;
  reg        [7:0]    _zz_io_MatrixB_55_28;
  reg        [7:0]    _zz_io_MatrixB_55_29;
  reg        [7:0]    _zz_io_MatrixB_55_30;
  reg        [7:0]    _zz_io_MatrixB_55_31;
  reg        [7:0]    _zz_io_MatrixB_55_32;
  reg        [7:0]    _zz_io_MatrixB_55_33;
  reg        [7:0]    _zz_io_MatrixB_55_34;
  reg        [7:0]    _zz_io_MatrixB_55_35;
  reg        [7:0]    _zz_io_MatrixB_55_36;
  reg        [7:0]    _zz_io_MatrixB_55_37;
  reg        [7:0]    _zz_io_MatrixB_55_38;
  reg        [7:0]    _zz_io_MatrixB_55_39;
  reg        [7:0]    _zz_io_MatrixB_55_40;
  reg        [7:0]    _zz_io_MatrixB_55_41;
  reg        [7:0]    _zz_io_MatrixB_55_42;
  reg        [7:0]    _zz_io_MatrixB_55_43;
  reg        [7:0]    _zz_io_MatrixB_55_44;
  reg        [7:0]    _zz_io_MatrixB_55_45;
  reg        [7:0]    _zz_io_MatrixB_55_46;
  reg        [7:0]    _zz_io_MatrixB_55_47;
  reg        [7:0]    _zz_io_MatrixB_55_48;
  reg        [7:0]    _zz_io_MatrixB_55_49;
  reg        [7:0]    _zz_io_MatrixB_55_50;
  reg        [7:0]    _zz_io_MatrixB_55_51;
  reg        [7:0]    _zz_io_MatrixB_55_52;
  reg        [7:0]    _zz_io_MatrixB_55_53;
  reg        [7:0]    _zz_io_MatrixB_55_54;
  reg                 _zz_io_B_Valid_55;
  reg                 _zz_io_B_Valid_55_1;
  reg                 _zz_io_B_Valid_55_2;
  reg                 _zz_io_B_Valid_55_3;
  reg                 _zz_io_B_Valid_55_4;
  reg                 _zz_io_B_Valid_55_5;
  reg                 _zz_io_B_Valid_55_6;
  reg                 _zz_io_B_Valid_55_7;
  reg                 _zz_io_B_Valid_55_8;
  reg                 _zz_io_B_Valid_55_9;
  reg                 _zz_io_B_Valid_55_10;
  reg                 _zz_io_B_Valid_55_11;
  reg                 _zz_io_B_Valid_55_12;
  reg                 _zz_io_B_Valid_55_13;
  reg                 _zz_io_B_Valid_55_14;
  reg                 _zz_io_B_Valid_55_15;
  reg                 _zz_io_B_Valid_55_16;
  reg                 _zz_io_B_Valid_55_17;
  reg                 _zz_io_B_Valid_55_18;
  reg                 _zz_io_B_Valid_55_19;
  reg                 _zz_io_B_Valid_55_20;
  reg                 _zz_io_B_Valid_55_21;
  reg                 _zz_io_B_Valid_55_22;
  reg                 _zz_io_B_Valid_55_23;
  reg                 _zz_io_B_Valid_55_24;
  reg                 _zz_io_B_Valid_55_25;
  reg                 _zz_io_B_Valid_55_26;
  reg                 _zz_io_B_Valid_55_27;
  reg                 _zz_io_B_Valid_55_28;
  reg                 _zz_io_B_Valid_55_29;
  reg                 _zz_io_B_Valid_55_30;
  reg                 _zz_io_B_Valid_55_31;
  reg                 _zz_io_B_Valid_55_32;
  reg                 _zz_io_B_Valid_55_33;
  reg                 _zz_io_B_Valid_55_34;
  reg                 _zz_io_B_Valid_55_35;
  reg                 _zz_io_B_Valid_55_36;
  reg                 _zz_io_B_Valid_55_37;
  reg                 _zz_io_B_Valid_55_38;
  reg                 _zz_io_B_Valid_55_39;
  reg                 _zz_io_B_Valid_55_40;
  reg                 _zz_io_B_Valid_55_41;
  reg                 _zz_io_B_Valid_55_42;
  reg                 _zz_io_B_Valid_55_43;
  reg                 _zz_io_B_Valid_55_44;
  reg                 _zz_io_B_Valid_55_45;
  reg                 _zz_io_B_Valid_55_46;
  reg                 _zz_io_B_Valid_55_47;
  reg                 _zz_io_B_Valid_55_48;
  reg                 _zz_io_B_Valid_55_49;
  reg                 _zz_io_B_Valid_55_50;
  reg                 _zz_io_B_Valid_55_51;
  reg                 _zz_io_B_Valid_55_52;
  reg                 _zz_io_B_Valid_55_53;
  reg                 _zz_io_B_Valid_55_54;
  reg        [7:0]    _zz_io_MatrixB_56;
  reg        [7:0]    _zz_io_MatrixB_56_1;
  reg        [7:0]    _zz_io_MatrixB_56_2;
  reg        [7:0]    _zz_io_MatrixB_56_3;
  reg        [7:0]    _zz_io_MatrixB_56_4;
  reg        [7:0]    _zz_io_MatrixB_56_5;
  reg        [7:0]    _zz_io_MatrixB_56_6;
  reg        [7:0]    _zz_io_MatrixB_56_7;
  reg        [7:0]    _zz_io_MatrixB_56_8;
  reg        [7:0]    _zz_io_MatrixB_56_9;
  reg        [7:0]    _zz_io_MatrixB_56_10;
  reg        [7:0]    _zz_io_MatrixB_56_11;
  reg        [7:0]    _zz_io_MatrixB_56_12;
  reg        [7:0]    _zz_io_MatrixB_56_13;
  reg        [7:0]    _zz_io_MatrixB_56_14;
  reg        [7:0]    _zz_io_MatrixB_56_15;
  reg        [7:0]    _zz_io_MatrixB_56_16;
  reg        [7:0]    _zz_io_MatrixB_56_17;
  reg        [7:0]    _zz_io_MatrixB_56_18;
  reg        [7:0]    _zz_io_MatrixB_56_19;
  reg        [7:0]    _zz_io_MatrixB_56_20;
  reg        [7:0]    _zz_io_MatrixB_56_21;
  reg        [7:0]    _zz_io_MatrixB_56_22;
  reg        [7:0]    _zz_io_MatrixB_56_23;
  reg        [7:0]    _zz_io_MatrixB_56_24;
  reg        [7:0]    _zz_io_MatrixB_56_25;
  reg        [7:0]    _zz_io_MatrixB_56_26;
  reg        [7:0]    _zz_io_MatrixB_56_27;
  reg        [7:0]    _zz_io_MatrixB_56_28;
  reg        [7:0]    _zz_io_MatrixB_56_29;
  reg        [7:0]    _zz_io_MatrixB_56_30;
  reg        [7:0]    _zz_io_MatrixB_56_31;
  reg        [7:0]    _zz_io_MatrixB_56_32;
  reg        [7:0]    _zz_io_MatrixB_56_33;
  reg        [7:0]    _zz_io_MatrixB_56_34;
  reg        [7:0]    _zz_io_MatrixB_56_35;
  reg        [7:0]    _zz_io_MatrixB_56_36;
  reg        [7:0]    _zz_io_MatrixB_56_37;
  reg        [7:0]    _zz_io_MatrixB_56_38;
  reg        [7:0]    _zz_io_MatrixB_56_39;
  reg        [7:0]    _zz_io_MatrixB_56_40;
  reg        [7:0]    _zz_io_MatrixB_56_41;
  reg        [7:0]    _zz_io_MatrixB_56_42;
  reg        [7:0]    _zz_io_MatrixB_56_43;
  reg        [7:0]    _zz_io_MatrixB_56_44;
  reg        [7:0]    _zz_io_MatrixB_56_45;
  reg        [7:0]    _zz_io_MatrixB_56_46;
  reg        [7:0]    _zz_io_MatrixB_56_47;
  reg        [7:0]    _zz_io_MatrixB_56_48;
  reg        [7:0]    _zz_io_MatrixB_56_49;
  reg        [7:0]    _zz_io_MatrixB_56_50;
  reg        [7:0]    _zz_io_MatrixB_56_51;
  reg        [7:0]    _zz_io_MatrixB_56_52;
  reg        [7:0]    _zz_io_MatrixB_56_53;
  reg        [7:0]    _zz_io_MatrixB_56_54;
  reg        [7:0]    _zz_io_MatrixB_56_55;
  reg                 _zz_io_B_Valid_56;
  reg                 _zz_io_B_Valid_56_1;
  reg                 _zz_io_B_Valid_56_2;
  reg                 _zz_io_B_Valid_56_3;
  reg                 _zz_io_B_Valid_56_4;
  reg                 _zz_io_B_Valid_56_5;
  reg                 _zz_io_B_Valid_56_6;
  reg                 _zz_io_B_Valid_56_7;
  reg                 _zz_io_B_Valid_56_8;
  reg                 _zz_io_B_Valid_56_9;
  reg                 _zz_io_B_Valid_56_10;
  reg                 _zz_io_B_Valid_56_11;
  reg                 _zz_io_B_Valid_56_12;
  reg                 _zz_io_B_Valid_56_13;
  reg                 _zz_io_B_Valid_56_14;
  reg                 _zz_io_B_Valid_56_15;
  reg                 _zz_io_B_Valid_56_16;
  reg                 _zz_io_B_Valid_56_17;
  reg                 _zz_io_B_Valid_56_18;
  reg                 _zz_io_B_Valid_56_19;
  reg                 _zz_io_B_Valid_56_20;
  reg                 _zz_io_B_Valid_56_21;
  reg                 _zz_io_B_Valid_56_22;
  reg                 _zz_io_B_Valid_56_23;
  reg                 _zz_io_B_Valid_56_24;
  reg                 _zz_io_B_Valid_56_25;
  reg                 _zz_io_B_Valid_56_26;
  reg                 _zz_io_B_Valid_56_27;
  reg                 _zz_io_B_Valid_56_28;
  reg                 _zz_io_B_Valid_56_29;
  reg                 _zz_io_B_Valid_56_30;
  reg                 _zz_io_B_Valid_56_31;
  reg                 _zz_io_B_Valid_56_32;
  reg                 _zz_io_B_Valid_56_33;
  reg                 _zz_io_B_Valid_56_34;
  reg                 _zz_io_B_Valid_56_35;
  reg                 _zz_io_B_Valid_56_36;
  reg                 _zz_io_B_Valid_56_37;
  reg                 _zz_io_B_Valid_56_38;
  reg                 _zz_io_B_Valid_56_39;
  reg                 _zz_io_B_Valid_56_40;
  reg                 _zz_io_B_Valid_56_41;
  reg                 _zz_io_B_Valid_56_42;
  reg                 _zz_io_B_Valid_56_43;
  reg                 _zz_io_B_Valid_56_44;
  reg                 _zz_io_B_Valid_56_45;
  reg                 _zz_io_B_Valid_56_46;
  reg                 _zz_io_B_Valid_56_47;
  reg                 _zz_io_B_Valid_56_48;
  reg                 _zz_io_B_Valid_56_49;
  reg                 _zz_io_B_Valid_56_50;
  reg                 _zz_io_B_Valid_56_51;
  reg                 _zz_io_B_Valid_56_52;
  reg                 _zz_io_B_Valid_56_53;
  reg                 _zz_io_B_Valid_56_54;
  reg                 _zz_io_B_Valid_56_55;
  reg        [7:0]    _zz_io_MatrixB_57;
  reg        [7:0]    _zz_io_MatrixB_57_1;
  reg        [7:0]    _zz_io_MatrixB_57_2;
  reg        [7:0]    _zz_io_MatrixB_57_3;
  reg        [7:0]    _zz_io_MatrixB_57_4;
  reg        [7:0]    _zz_io_MatrixB_57_5;
  reg        [7:0]    _zz_io_MatrixB_57_6;
  reg        [7:0]    _zz_io_MatrixB_57_7;
  reg        [7:0]    _zz_io_MatrixB_57_8;
  reg        [7:0]    _zz_io_MatrixB_57_9;
  reg        [7:0]    _zz_io_MatrixB_57_10;
  reg        [7:0]    _zz_io_MatrixB_57_11;
  reg        [7:0]    _zz_io_MatrixB_57_12;
  reg        [7:0]    _zz_io_MatrixB_57_13;
  reg        [7:0]    _zz_io_MatrixB_57_14;
  reg        [7:0]    _zz_io_MatrixB_57_15;
  reg        [7:0]    _zz_io_MatrixB_57_16;
  reg        [7:0]    _zz_io_MatrixB_57_17;
  reg        [7:0]    _zz_io_MatrixB_57_18;
  reg        [7:0]    _zz_io_MatrixB_57_19;
  reg        [7:0]    _zz_io_MatrixB_57_20;
  reg        [7:0]    _zz_io_MatrixB_57_21;
  reg        [7:0]    _zz_io_MatrixB_57_22;
  reg        [7:0]    _zz_io_MatrixB_57_23;
  reg        [7:0]    _zz_io_MatrixB_57_24;
  reg        [7:0]    _zz_io_MatrixB_57_25;
  reg        [7:0]    _zz_io_MatrixB_57_26;
  reg        [7:0]    _zz_io_MatrixB_57_27;
  reg        [7:0]    _zz_io_MatrixB_57_28;
  reg        [7:0]    _zz_io_MatrixB_57_29;
  reg        [7:0]    _zz_io_MatrixB_57_30;
  reg        [7:0]    _zz_io_MatrixB_57_31;
  reg        [7:0]    _zz_io_MatrixB_57_32;
  reg        [7:0]    _zz_io_MatrixB_57_33;
  reg        [7:0]    _zz_io_MatrixB_57_34;
  reg        [7:0]    _zz_io_MatrixB_57_35;
  reg        [7:0]    _zz_io_MatrixB_57_36;
  reg        [7:0]    _zz_io_MatrixB_57_37;
  reg        [7:0]    _zz_io_MatrixB_57_38;
  reg        [7:0]    _zz_io_MatrixB_57_39;
  reg        [7:0]    _zz_io_MatrixB_57_40;
  reg        [7:0]    _zz_io_MatrixB_57_41;
  reg        [7:0]    _zz_io_MatrixB_57_42;
  reg        [7:0]    _zz_io_MatrixB_57_43;
  reg        [7:0]    _zz_io_MatrixB_57_44;
  reg        [7:0]    _zz_io_MatrixB_57_45;
  reg        [7:0]    _zz_io_MatrixB_57_46;
  reg        [7:0]    _zz_io_MatrixB_57_47;
  reg        [7:0]    _zz_io_MatrixB_57_48;
  reg        [7:0]    _zz_io_MatrixB_57_49;
  reg        [7:0]    _zz_io_MatrixB_57_50;
  reg        [7:0]    _zz_io_MatrixB_57_51;
  reg        [7:0]    _zz_io_MatrixB_57_52;
  reg        [7:0]    _zz_io_MatrixB_57_53;
  reg        [7:0]    _zz_io_MatrixB_57_54;
  reg        [7:0]    _zz_io_MatrixB_57_55;
  reg        [7:0]    _zz_io_MatrixB_57_56;
  reg                 _zz_io_B_Valid_57;
  reg                 _zz_io_B_Valid_57_1;
  reg                 _zz_io_B_Valid_57_2;
  reg                 _zz_io_B_Valid_57_3;
  reg                 _zz_io_B_Valid_57_4;
  reg                 _zz_io_B_Valid_57_5;
  reg                 _zz_io_B_Valid_57_6;
  reg                 _zz_io_B_Valid_57_7;
  reg                 _zz_io_B_Valid_57_8;
  reg                 _zz_io_B_Valid_57_9;
  reg                 _zz_io_B_Valid_57_10;
  reg                 _zz_io_B_Valid_57_11;
  reg                 _zz_io_B_Valid_57_12;
  reg                 _zz_io_B_Valid_57_13;
  reg                 _zz_io_B_Valid_57_14;
  reg                 _zz_io_B_Valid_57_15;
  reg                 _zz_io_B_Valid_57_16;
  reg                 _zz_io_B_Valid_57_17;
  reg                 _zz_io_B_Valid_57_18;
  reg                 _zz_io_B_Valid_57_19;
  reg                 _zz_io_B_Valid_57_20;
  reg                 _zz_io_B_Valid_57_21;
  reg                 _zz_io_B_Valid_57_22;
  reg                 _zz_io_B_Valid_57_23;
  reg                 _zz_io_B_Valid_57_24;
  reg                 _zz_io_B_Valid_57_25;
  reg                 _zz_io_B_Valid_57_26;
  reg                 _zz_io_B_Valid_57_27;
  reg                 _zz_io_B_Valid_57_28;
  reg                 _zz_io_B_Valid_57_29;
  reg                 _zz_io_B_Valid_57_30;
  reg                 _zz_io_B_Valid_57_31;
  reg                 _zz_io_B_Valid_57_32;
  reg                 _zz_io_B_Valid_57_33;
  reg                 _zz_io_B_Valid_57_34;
  reg                 _zz_io_B_Valid_57_35;
  reg                 _zz_io_B_Valid_57_36;
  reg                 _zz_io_B_Valid_57_37;
  reg                 _zz_io_B_Valid_57_38;
  reg                 _zz_io_B_Valid_57_39;
  reg                 _zz_io_B_Valid_57_40;
  reg                 _zz_io_B_Valid_57_41;
  reg                 _zz_io_B_Valid_57_42;
  reg                 _zz_io_B_Valid_57_43;
  reg                 _zz_io_B_Valid_57_44;
  reg                 _zz_io_B_Valid_57_45;
  reg                 _zz_io_B_Valid_57_46;
  reg                 _zz_io_B_Valid_57_47;
  reg                 _zz_io_B_Valid_57_48;
  reg                 _zz_io_B_Valid_57_49;
  reg                 _zz_io_B_Valid_57_50;
  reg                 _zz_io_B_Valid_57_51;
  reg                 _zz_io_B_Valid_57_52;
  reg                 _zz_io_B_Valid_57_53;
  reg                 _zz_io_B_Valid_57_54;
  reg                 _zz_io_B_Valid_57_55;
  reg                 _zz_io_B_Valid_57_56;
  reg        [7:0]    _zz_io_MatrixB_58;
  reg        [7:0]    _zz_io_MatrixB_58_1;
  reg        [7:0]    _zz_io_MatrixB_58_2;
  reg        [7:0]    _zz_io_MatrixB_58_3;
  reg        [7:0]    _zz_io_MatrixB_58_4;
  reg        [7:0]    _zz_io_MatrixB_58_5;
  reg        [7:0]    _zz_io_MatrixB_58_6;
  reg        [7:0]    _zz_io_MatrixB_58_7;
  reg        [7:0]    _zz_io_MatrixB_58_8;
  reg        [7:0]    _zz_io_MatrixB_58_9;
  reg        [7:0]    _zz_io_MatrixB_58_10;
  reg        [7:0]    _zz_io_MatrixB_58_11;
  reg        [7:0]    _zz_io_MatrixB_58_12;
  reg        [7:0]    _zz_io_MatrixB_58_13;
  reg        [7:0]    _zz_io_MatrixB_58_14;
  reg        [7:0]    _zz_io_MatrixB_58_15;
  reg        [7:0]    _zz_io_MatrixB_58_16;
  reg        [7:0]    _zz_io_MatrixB_58_17;
  reg        [7:0]    _zz_io_MatrixB_58_18;
  reg        [7:0]    _zz_io_MatrixB_58_19;
  reg        [7:0]    _zz_io_MatrixB_58_20;
  reg        [7:0]    _zz_io_MatrixB_58_21;
  reg        [7:0]    _zz_io_MatrixB_58_22;
  reg        [7:0]    _zz_io_MatrixB_58_23;
  reg        [7:0]    _zz_io_MatrixB_58_24;
  reg        [7:0]    _zz_io_MatrixB_58_25;
  reg        [7:0]    _zz_io_MatrixB_58_26;
  reg        [7:0]    _zz_io_MatrixB_58_27;
  reg        [7:0]    _zz_io_MatrixB_58_28;
  reg        [7:0]    _zz_io_MatrixB_58_29;
  reg        [7:0]    _zz_io_MatrixB_58_30;
  reg        [7:0]    _zz_io_MatrixB_58_31;
  reg        [7:0]    _zz_io_MatrixB_58_32;
  reg        [7:0]    _zz_io_MatrixB_58_33;
  reg        [7:0]    _zz_io_MatrixB_58_34;
  reg        [7:0]    _zz_io_MatrixB_58_35;
  reg        [7:0]    _zz_io_MatrixB_58_36;
  reg        [7:0]    _zz_io_MatrixB_58_37;
  reg        [7:0]    _zz_io_MatrixB_58_38;
  reg        [7:0]    _zz_io_MatrixB_58_39;
  reg        [7:0]    _zz_io_MatrixB_58_40;
  reg        [7:0]    _zz_io_MatrixB_58_41;
  reg        [7:0]    _zz_io_MatrixB_58_42;
  reg        [7:0]    _zz_io_MatrixB_58_43;
  reg        [7:0]    _zz_io_MatrixB_58_44;
  reg        [7:0]    _zz_io_MatrixB_58_45;
  reg        [7:0]    _zz_io_MatrixB_58_46;
  reg        [7:0]    _zz_io_MatrixB_58_47;
  reg        [7:0]    _zz_io_MatrixB_58_48;
  reg        [7:0]    _zz_io_MatrixB_58_49;
  reg        [7:0]    _zz_io_MatrixB_58_50;
  reg        [7:0]    _zz_io_MatrixB_58_51;
  reg        [7:0]    _zz_io_MatrixB_58_52;
  reg        [7:0]    _zz_io_MatrixB_58_53;
  reg        [7:0]    _zz_io_MatrixB_58_54;
  reg        [7:0]    _zz_io_MatrixB_58_55;
  reg        [7:0]    _zz_io_MatrixB_58_56;
  reg        [7:0]    _zz_io_MatrixB_58_57;
  reg                 _zz_io_B_Valid_58;
  reg                 _zz_io_B_Valid_58_1;
  reg                 _zz_io_B_Valid_58_2;
  reg                 _zz_io_B_Valid_58_3;
  reg                 _zz_io_B_Valid_58_4;
  reg                 _zz_io_B_Valid_58_5;
  reg                 _zz_io_B_Valid_58_6;
  reg                 _zz_io_B_Valid_58_7;
  reg                 _zz_io_B_Valid_58_8;
  reg                 _zz_io_B_Valid_58_9;
  reg                 _zz_io_B_Valid_58_10;
  reg                 _zz_io_B_Valid_58_11;
  reg                 _zz_io_B_Valid_58_12;
  reg                 _zz_io_B_Valid_58_13;
  reg                 _zz_io_B_Valid_58_14;
  reg                 _zz_io_B_Valid_58_15;
  reg                 _zz_io_B_Valid_58_16;
  reg                 _zz_io_B_Valid_58_17;
  reg                 _zz_io_B_Valid_58_18;
  reg                 _zz_io_B_Valid_58_19;
  reg                 _zz_io_B_Valid_58_20;
  reg                 _zz_io_B_Valid_58_21;
  reg                 _zz_io_B_Valid_58_22;
  reg                 _zz_io_B_Valid_58_23;
  reg                 _zz_io_B_Valid_58_24;
  reg                 _zz_io_B_Valid_58_25;
  reg                 _zz_io_B_Valid_58_26;
  reg                 _zz_io_B_Valid_58_27;
  reg                 _zz_io_B_Valid_58_28;
  reg                 _zz_io_B_Valid_58_29;
  reg                 _zz_io_B_Valid_58_30;
  reg                 _zz_io_B_Valid_58_31;
  reg                 _zz_io_B_Valid_58_32;
  reg                 _zz_io_B_Valid_58_33;
  reg                 _zz_io_B_Valid_58_34;
  reg                 _zz_io_B_Valid_58_35;
  reg                 _zz_io_B_Valid_58_36;
  reg                 _zz_io_B_Valid_58_37;
  reg                 _zz_io_B_Valid_58_38;
  reg                 _zz_io_B_Valid_58_39;
  reg                 _zz_io_B_Valid_58_40;
  reg                 _zz_io_B_Valid_58_41;
  reg                 _zz_io_B_Valid_58_42;
  reg                 _zz_io_B_Valid_58_43;
  reg                 _zz_io_B_Valid_58_44;
  reg                 _zz_io_B_Valid_58_45;
  reg                 _zz_io_B_Valid_58_46;
  reg                 _zz_io_B_Valid_58_47;
  reg                 _zz_io_B_Valid_58_48;
  reg                 _zz_io_B_Valid_58_49;
  reg                 _zz_io_B_Valid_58_50;
  reg                 _zz_io_B_Valid_58_51;
  reg                 _zz_io_B_Valid_58_52;
  reg                 _zz_io_B_Valid_58_53;
  reg                 _zz_io_B_Valid_58_54;
  reg                 _zz_io_B_Valid_58_55;
  reg                 _zz_io_B_Valid_58_56;
  reg                 _zz_io_B_Valid_58_57;
  reg        [7:0]    _zz_io_MatrixB_59;
  reg        [7:0]    _zz_io_MatrixB_59_1;
  reg        [7:0]    _zz_io_MatrixB_59_2;
  reg        [7:0]    _zz_io_MatrixB_59_3;
  reg        [7:0]    _zz_io_MatrixB_59_4;
  reg        [7:0]    _zz_io_MatrixB_59_5;
  reg        [7:0]    _zz_io_MatrixB_59_6;
  reg        [7:0]    _zz_io_MatrixB_59_7;
  reg        [7:0]    _zz_io_MatrixB_59_8;
  reg        [7:0]    _zz_io_MatrixB_59_9;
  reg        [7:0]    _zz_io_MatrixB_59_10;
  reg        [7:0]    _zz_io_MatrixB_59_11;
  reg        [7:0]    _zz_io_MatrixB_59_12;
  reg        [7:0]    _zz_io_MatrixB_59_13;
  reg        [7:0]    _zz_io_MatrixB_59_14;
  reg        [7:0]    _zz_io_MatrixB_59_15;
  reg        [7:0]    _zz_io_MatrixB_59_16;
  reg        [7:0]    _zz_io_MatrixB_59_17;
  reg        [7:0]    _zz_io_MatrixB_59_18;
  reg        [7:0]    _zz_io_MatrixB_59_19;
  reg        [7:0]    _zz_io_MatrixB_59_20;
  reg        [7:0]    _zz_io_MatrixB_59_21;
  reg        [7:0]    _zz_io_MatrixB_59_22;
  reg        [7:0]    _zz_io_MatrixB_59_23;
  reg        [7:0]    _zz_io_MatrixB_59_24;
  reg        [7:0]    _zz_io_MatrixB_59_25;
  reg        [7:0]    _zz_io_MatrixB_59_26;
  reg        [7:0]    _zz_io_MatrixB_59_27;
  reg        [7:0]    _zz_io_MatrixB_59_28;
  reg        [7:0]    _zz_io_MatrixB_59_29;
  reg        [7:0]    _zz_io_MatrixB_59_30;
  reg        [7:0]    _zz_io_MatrixB_59_31;
  reg        [7:0]    _zz_io_MatrixB_59_32;
  reg        [7:0]    _zz_io_MatrixB_59_33;
  reg        [7:0]    _zz_io_MatrixB_59_34;
  reg        [7:0]    _zz_io_MatrixB_59_35;
  reg        [7:0]    _zz_io_MatrixB_59_36;
  reg        [7:0]    _zz_io_MatrixB_59_37;
  reg        [7:0]    _zz_io_MatrixB_59_38;
  reg        [7:0]    _zz_io_MatrixB_59_39;
  reg        [7:0]    _zz_io_MatrixB_59_40;
  reg        [7:0]    _zz_io_MatrixB_59_41;
  reg        [7:0]    _zz_io_MatrixB_59_42;
  reg        [7:0]    _zz_io_MatrixB_59_43;
  reg        [7:0]    _zz_io_MatrixB_59_44;
  reg        [7:0]    _zz_io_MatrixB_59_45;
  reg        [7:0]    _zz_io_MatrixB_59_46;
  reg        [7:0]    _zz_io_MatrixB_59_47;
  reg        [7:0]    _zz_io_MatrixB_59_48;
  reg        [7:0]    _zz_io_MatrixB_59_49;
  reg        [7:0]    _zz_io_MatrixB_59_50;
  reg        [7:0]    _zz_io_MatrixB_59_51;
  reg        [7:0]    _zz_io_MatrixB_59_52;
  reg        [7:0]    _zz_io_MatrixB_59_53;
  reg        [7:0]    _zz_io_MatrixB_59_54;
  reg        [7:0]    _zz_io_MatrixB_59_55;
  reg        [7:0]    _zz_io_MatrixB_59_56;
  reg        [7:0]    _zz_io_MatrixB_59_57;
  reg        [7:0]    _zz_io_MatrixB_59_58;
  reg                 _zz_io_B_Valid_59;
  reg                 _zz_io_B_Valid_59_1;
  reg                 _zz_io_B_Valid_59_2;
  reg                 _zz_io_B_Valid_59_3;
  reg                 _zz_io_B_Valid_59_4;
  reg                 _zz_io_B_Valid_59_5;
  reg                 _zz_io_B_Valid_59_6;
  reg                 _zz_io_B_Valid_59_7;
  reg                 _zz_io_B_Valid_59_8;
  reg                 _zz_io_B_Valid_59_9;
  reg                 _zz_io_B_Valid_59_10;
  reg                 _zz_io_B_Valid_59_11;
  reg                 _zz_io_B_Valid_59_12;
  reg                 _zz_io_B_Valid_59_13;
  reg                 _zz_io_B_Valid_59_14;
  reg                 _zz_io_B_Valid_59_15;
  reg                 _zz_io_B_Valid_59_16;
  reg                 _zz_io_B_Valid_59_17;
  reg                 _zz_io_B_Valid_59_18;
  reg                 _zz_io_B_Valid_59_19;
  reg                 _zz_io_B_Valid_59_20;
  reg                 _zz_io_B_Valid_59_21;
  reg                 _zz_io_B_Valid_59_22;
  reg                 _zz_io_B_Valid_59_23;
  reg                 _zz_io_B_Valid_59_24;
  reg                 _zz_io_B_Valid_59_25;
  reg                 _zz_io_B_Valid_59_26;
  reg                 _zz_io_B_Valid_59_27;
  reg                 _zz_io_B_Valid_59_28;
  reg                 _zz_io_B_Valid_59_29;
  reg                 _zz_io_B_Valid_59_30;
  reg                 _zz_io_B_Valid_59_31;
  reg                 _zz_io_B_Valid_59_32;
  reg                 _zz_io_B_Valid_59_33;
  reg                 _zz_io_B_Valid_59_34;
  reg                 _zz_io_B_Valid_59_35;
  reg                 _zz_io_B_Valid_59_36;
  reg                 _zz_io_B_Valid_59_37;
  reg                 _zz_io_B_Valid_59_38;
  reg                 _zz_io_B_Valid_59_39;
  reg                 _zz_io_B_Valid_59_40;
  reg                 _zz_io_B_Valid_59_41;
  reg                 _zz_io_B_Valid_59_42;
  reg                 _zz_io_B_Valid_59_43;
  reg                 _zz_io_B_Valid_59_44;
  reg                 _zz_io_B_Valid_59_45;
  reg                 _zz_io_B_Valid_59_46;
  reg                 _zz_io_B_Valid_59_47;
  reg                 _zz_io_B_Valid_59_48;
  reg                 _zz_io_B_Valid_59_49;
  reg                 _zz_io_B_Valid_59_50;
  reg                 _zz_io_B_Valid_59_51;
  reg                 _zz_io_B_Valid_59_52;
  reg                 _zz_io_B_Valid_59_53;
  reg                 _zz_io_B_Valid_59_54;
  reg                 _zz_io_B_Valid_59_55;
  reg                 _zz_io_B_Valid_59_56;
  reg                 _zz_io_B_Valid_59_57;
  reg                 _zz_io_B_Valid_59_58;
  reg        [7:0]    _zz_io_MatrixB_60;
  reg        [7:0]    _zz_io_MatrixB_60_1;
  reg        [7:0]    _zz_io_MatrixB_60_2;
  reg        [7:0]    _zz_io_MatrixB_60_3;
  reg        [7:0]    _zz_io_MatrixB_60_4;
  reg        [7:0]    _zz_io_MatrixB_60_5;
  reg        [7:0]    _zz_io_MatrixB_60_6;
  reg        [7:0]    _zz_io_MatrixB_60_7;
  reg        [7:0]    _zz_io_MatrixB_60_8;
  reg        [7:0]    _zz_io_MatrixB_60_9;
  reg        [7:0]    _zz_io_MatrixB_60_10;
  reg        [7:0]    _zz_io_MatrixB_60_11;
  reg        [7:0]    _zz_io_MatrixB_60_12;
  reg        [7:0]    _zz_io_MatrixB_60_13;
  reg        [7:0]    _zz_io_MatrixB_60_14;
  reg        [7:0]    _zz_io_MatrixB_60_15;
  reg        [7:0]    _zz_io_MatrixB_60_16;
  reg        [7:0]    _zz_io_MatrixB_60_17;
  reg        [7:0]    _zz_io_MatrixB_60_18;
  reg        [7:0]    _zz_io_MatrixB_60_19;
  reg        [7:0]    _zz_io_MatrixB_60_20;
  reg        [7:0]    _zz_io_MatrixB_60_21;
  reg        [7:0]    _zz_io_MatrixB_60_22;
  reg        [7:0]    _zz_io_MatrixB_60_23;
  reg        [7:0]    _zz_io_MatrixB_60_24;
  reg        [7:0]    _zz_io_MatrixB_60_25;
  reg        [7:0]    _zz_io_MatrixB_60_26;
  reg        [7:0]    _zz_io_MatrixB_60_27;
  reg        [7:0]    _zz_io_MatrixB_60_28;
  reg        [7:0]    _zz_io_MatrixB_60_29;
  reg        [7:0]    _zz_io_MatrixB_60_30;
  reg        [7:0]    _zz_io_MatrixB_60_31;
  reg        [7:0]    _zz_io_MatrixB_60_32;
  reg        [7:0]    _zz_io_MatrixB_60_33;
  reg        [7:0]    _zz_io_MatrixB_60_34;
  reg        [7:0]    _zz_io_MatrixB_60_35;
  reg        [7:0]    _zz_io_MatrixB_60_36;
  reg        [7:0]    _zz_io_MatrixB_60_37;
  reg        [7:0]    _zz_io_MatrixB_60_38;
  reg        [7:0]    _zz_io_MatrixB_60_39;
  reg        [7:0]    _zz_io_MatrixB_60_40;
  reg        [7:0]    _zz_io_MatrixB_60_41;
  reg        [7:0]    _zz_io_MatrixB_60_42;
  reg        [7:0]    _zz_io_MatrixB_60_43;
  reg        [7:0]    _zz_io_MatrixB_60_44;
  reg        [7:0]    _zz_io_MatrixB_60_45;
  reg        [7:0]    _zz_io_MatrixB_60_46;
  reg        [7:0]    _zz_io_MatrixB_60_47;
  reg        [7:0]    _zz_io_MatrixB_60_48;
  reg        [7:0]    _zz_io_MatrixB_60_49;
  reg        [7:0]    _zz_io_MatrixB_60_50;
  reg        [7:0]    _zz_io_MatrixB_60_51;
  reg        [7:0]    _zz_io_MatrixB_60_52;
  reg        [7:0]    _zz_io_MatrixB_60_53;
  reg        [7:0]    _zz_io_MatrixB_60_54;
  reg        [7:0]    _zz_io_MatrixB_60_55;
  reg        [7:0]    _zz_io_MatrixB_60_56;
  reg        [7:0]    _zz_io_MatrixB_60_57;
  reg        [7:0]    _zz_io_MatrixB_60_58;
  reg        [7:0]    _zz_io_MatrixB_60_59;
  reg                 _zz_io_B_Valid_60;
  reg                 _zz_io_B_Valid_60_1;
  reg                 _zz_io_B_Valid_60_2;
  reg                 _zz_io_B_Valid_60_3;
  reg                 _zz_io_B_Valid_60_4;
  reg                 _zz_io_B_Valid_60_5;
  reg                 _zz_io_B_Valid_60_6;
  reg                 _zz_io_B_Valid_60_7;
  reg                 _zz_io_B_Valid_60_8;
  reg                 _zz_io_B_Valid_60_9;
  reg                 _zz_io_B_Valid_60_10;
  reg                 _zz_io_B_Valid_60_11;
  reg                 _zz_io_B_Valid_60_12;
  reg                 _zz_io_B_Valid_60_13;
  reg                 _zz_io_B_Valid_60_14;
  reg                 _zz_io_B_Valid_60_15;
  reg                 _zz_io_B_Valid_60_16;
  reg                 _zz_io_B_Valid_60_17;
  reg                 _zz_io_B_Valid_60_18;
  reg                 _zz_io_B_Valid_60_19;
  reg                 _zz_io_B_Valid_60_20;
  reg                 _zz_io_B_Valid_60_21;
  reg                 _zz_io_B_Valid_60_22;
  reg                 _zz_io_B_Valid_60_23;
  reg                 _zz_io_B_Valid_60_24;
  reg                 _zz_io_B_Valid_60_25;
  reg                 _zz_io_B_Valid_60_26;
  reg                 _zz_io_B_Valid_60_27;
  reg                 _zz_io_B_Valid_60_28;
  reg                 _zz_io_B_Valid_60_29;
  reg                 _zz_io_B_Valid_60_30;
  reg                 _zz_io_B_Valid_60_31;
  reg                 _zz_io_B_Valid_60_32;
  reg                 _zz_io_B_Valid_60_33;
  reg                 _zz_io_B_Valid_60_34;
  reg                 _zz_io_B_Valid_60_35;
  reg                 _zz_io_B_Valid_60_36;
  reg                 _zz_io_B_Valid_60_37;
  reg                 _zz_io_B_Valid_60_38;
  reg                 _zz_io_B_Valid_60_39;
  reg                 _zz_io_B_Valid_60_40;
  reg                 _zz_io_B_Valid_60_41;
  reg                 _zz_io_B_Valid_60_42;
  reg                 _zz_io_B_Valid_60_43;
  reg                 _zz_io_B_Valid_60_44;
  reg                 _zz_io_B_Valid_60_45;
  reg                 _zz_io_B_Valid_60_46;
  reg                 _zz_io_B_Valid_60_47;
  reg                 _zz_io_B_Valid_60_48;
  reg                 _zz_io_B_Valid_60_49;
  reg                 _zz_io_B_Valid_60_50;
  reg                 _zz_io_B_Valid_60_51;
  reg                 _zz_io_B_Valid_60_52;
  reg                 _zz_io_B_Valid_60_53;
  reg                 _zz_io_B_Valid_60_54;
  reg                 _zz_io_B_Valid_60_55;
  reg                 _zz_io_B_Valid_60_56;
  reg                 _zz_io_B_Valid_60_57;
  reg                 _zz_io_B_Valid_60_58;
  reg                 _zz_io_B_Valid_60_59;
  reg        [7:0]    _zz_io_MatrixB_61;
  reg        [7:0]    _zz_io_MatrixB_61_1;
  reg        [7:0]    _zz_io_MatrixB_61_2;
  reg        [7:0]    _zz_io_MatrixB_61_3;
  reg        [7:0]    _zz_io_MatrixB_61_4;
  reg        [7:0]    _zz_io_MatrixB_61_5;
  reg        [7:0]    _zz_io_MatrixB_61_6;
  reg        [7:0]    _zz_io_MatrixB_61_7;
  reg        [7:0]    _zz_io_MatrixB_61_8;
  reg        [7:0]    _zz_io_MatrixB_61_9;
  reg        [7:0]    _zz_io_MatrixB_61_10;
  reg        [7:0]    _zz_io_MatrixB_61_11;
  reg        [7:0]    _zz_io_MatrixB_61_12;
  reg        [7:0]    _zz_io_MatrixB_61_13;
  reg        [7:0]    _zz_io_MatrixB_61_14;
  reg        [7:0]    _zz_io_MatrixB_61_15;
  reg        [7:0]    _zz_io_MatrixB_61_16;
  reg        [7:0]    _zz_io_MatrixB_61_17;
  reg        [7:0]    _zz_io_MatrixB_61_18;
  reg        [7:0]    _zz_io_MatrixB_61_19;
  reg        [7:0]    _zz_io_MatrixB_61_20;
  reg        [7:0]    _zz_io_MatrixB_61_21;
  reg        [7:0]    _zz_io_MatrixB_61_22;
  reg        [7:0]    _zz_io_MatrixB_61_23;
  reg        [7:0]    _zz_io_MatrixB_61_24;
  reg        [7:0]    _zz_io_MatrixB_61_25;
  reg        [7:0]    _zz_io_MatrixB_61_26;
  reg        [7:0]    _zz_io_MatrixB_61_27;
  reg        [7:0]    _zz_io_MatrixB_61_28;
  reg        [7:0]    _zz_io_MatrixB_61_29;
  reg        [7:0]    _zz_io_MatrixB_61_30;
  reg        [7:0]    _zz_io_MatrixB_61_31;
  reg        [7:0]    _zz_io_MatrixB_61_32;
  reg        [7:0]    _zz_io_MatrixB_61_33;
  reg        [7:0]    _zz_io_MatrixB_61_34;
  reg        [7:0]    _zz_io_MatrixB_61_35;
  reg        [7:0]    _zz_io_MatrixB_61_36;
  reg        [7:0]    _zz_io_MatrixB_61_37;
  reg        [7:0]    _zz_io_MatrixB_61_38;
  reg        [7:0]    _zz_io_MatrixB_61_39;
  reg        [7:0]    _zz_io_MatrixB_61_40;
  reg        [7:0]    _zz_io_MatrixB_61_41;
  reg        [7:0]    _zz_io_MatrixB_61_42;
  reg        [7:0]    _zz_io_MatrixB_61_43;
  reg        [7:0]    _zz_io_MatrixB_61_44;
  reg        [7:0]    _zz_io_MatrixB_61_45;
  reg        [7:0]    _zz_io_MatrixB_61_46;
  reg        [7:0]    _zz_io_MatrixB_61_47;
  reg        [7:0]    _zz_io_MatrixB_61_48;
  reg        [7:0]    _zz_io_MatrixB_61_49;
  reg        [7:0]    _zz_io_MatrixB_61_50;
  reg        [7:0]    _zz_io_MatrixB_61_51;
  reg        [7:0]    _zz_io_MatrixB_61_52;
  reg        [7:0]    _zz_io_MatrixB_61_53;
  reg        [7:0]    _zz_io_MatrixB_61_54;
  reg        [7:0]    _zz_io_MatrixB_61_55;
  reg        [7:0]    _zz_io_MatrixB_61_56;
  reg        [7:0]    _zz_io_MatrixB_61_57;
  reg        [7:0]    _zz_io_MatrixB_61_58;
  reg        [7:0]    _zz_io_MatrixB_61_59;
  reg        [7:0]    _zz_io_MatrixB_61_60;
  reg                 _zz_io_B_Valid_61;
  reg                 _zz_io_B_Valid_61_1;
  reg                 _zz_io_B_Valid_61_2;
  reg                 _zz_io_B_Valid_61_3;
  reg                 _zz_io_B_Valid_61_4;
  reg                 _zz_io_B_Valid_61_5;
  reg                 _zz_io_B_Valid_61_6;
  reg                 _zz_io_B_Valid_61_7;
  reg                 _zz_io_B_Valid_61_8;
  reg                 _zz_io_B_Valid_61_9;
  reg                 _zz_io_B_Valid_61_10;
  reg                 _zz_io_B_Valid_61_11;
  reg                 _zz_io_B_Valid_61_12;
  reg                 _zz_io_B_Valid_61_13;
  reg                 _zz_io_B_Valid_61_14;
  reg                 _zz_io_B_Valid_61_15;
  reg                 _zz_io_B_Valid_61_16;
  reg                 _zz_io_B_Valid_61_17;
  reg                 _zz_io_B_Valid_61_18;
  reg                 _zz_io_B_Valid_61_19;
  reg                 _zz_io_B_Valid_61_20;
  reg                 _zz_io_B_Valid_61_21;
  reg                 _zz_io_B_Valid_61_22;
  reg                 _zz_io_B_Valid_61_23;
  reg                 _zz_io_B_Valid_61_24;
  reg                 _zz_io_B_Valid_61_25;
  reg                 _zz_io_B_Valid_61_26;
  reg                 _zz_io_B_Valid_61_27;
  reg                 _zz_io_B_Valid_61_28;
  reg                 _zz_io_B_Valid_61_29;
  reg                 _zz_io_B_Valid_61_30;
  reg                 _zz_io_B_Valid_61_31;
  reg                 _zz_io_B_Valid_61_32;
  reg                 _zz_io_B_Valid_61_33;
  reg                 _zz_io_B_Valid_61_34;
  reg                 _zz_io_B_Valid_61_35;
  reg                 _zz_io_B_Valid_61_36;
  reg                 _zz_io_B_Valid_61_37;
  reg                 _zz_io_B_Valid_61_38;
  reg                 _zz_io_B_Valid_61_39;
  reg                 _zz_io_B_Valid_61_40;
  reg                 _zz_io_B_Valid_61_41;
  reg                 _zz_io_B_Valid_61_42;
  reg                 _zz_io_B_Valid_61_43;
  reg                 _zz_io_B_Valid_61_44;
  reg                 _zz_io_B_Valid_61_45;
  reg                 _zz_io_B_Valid_61_46;
  reg                 _zz_io_B_Valid_61_47;
  reg                 _zz_io_B_Valid_61_48;
  reg                 _zz_io_B_Valid_61_49;
  reg                 _zz_io_B_Valid_61_50;
  reg                 _zz_io_B_Valid_61_51;
  reg                 _zz_io_B_Valid_61_52;
  reg                 _zz_io_B_Valid_61_53;
  reg                 _zz_io_B_Valid_61_54;
  reg                 _zz_io_B_Valid_61_55;
  reg                 _zz_io_B_Valid_61_56;
  reg                 _zz_io_B_Valid_61_57;
  reg                 _zz_io_B_Valid_61_58;
  reg                 _zz_io_B_Valid_61_59;
  reg                 _zz_io_B_Valid_61_60;
  reg        [7:0]    _zz_io_MatrixB_62;
  reg        [7:0]    _zz_io_MatrixB_62_1;
  reg        [7:0]    _zz_io_MatrixB_62_2;
  reg        [7:0]    _zz_io_MatrixB_62_3;
  reg        [7:0]    _zz_io_MatrixB_62_4;
  reg        [7:0]    _zz_io_MatrixB_62_5;
  reg        [7:0]    _zz_io_MatrixB_62_6;
  reg        [7:0]    _zz_io_MatrixB_62_7;
  reg        [7:0]    _zz_io_MatrixB_62_8;
  reg        [7:0]    _zz_io_MatrixB_62_9;
  reg        [7:0]    _zz_io_MatrixB_62_10;
  reg        [7:0]    _zz_io_MatrixB_62_11;
  reg        [7:0]    _zz_io_MatrixB_62_12;
  reg        [7:0]    _zz_io_MatrixB_62_13;
  reg        [7:0]    _zz_io_MatrixB_62_14;
  reg        [7:0]    _zz_io_MatrixB_62_15;
  reg        [7:0]    _zz_io_MatrixB_62_16;
  reg        [7:0]    _zz_io_MatrixB_62_17;
  reg        [7:0]    _zz_io_MatrixB_62_18;
  reg        [7:0]    _zz_io_MatrixB_62_19;
  reg        [7:0]    _zz_io_MatrixB_62_20;
  reg        [7:0]    _zz_io_MatrixB_62_21;
  reg        [7:0]    _zz_io_MatrixB_62_22;
  reg        [7:0]    _zz_io_MatrixB_62_23;
  reg        [7:0]    _zz_io_MatrixB_62_24;
  reg        [7:0]    _zz_io_MatrixB_62_25;
  reg        [7:0]    _zz_io_MatrixB_62_26;
  reg        [7:0]    _zz_io_MatrixB_62_27;
  reg        [7:0]    _zz_io_MatrixB_62_28;
  reg        [7:0]    _zz_io_MatrixB_62_29;
  reg        [7:0]    _zz_io_MatrixB_62_30;
  reg        [7:0]    _zz_io_MatrixB_62_31;
  reg        [7:0]    _zz_io_MatrixB_62_32;
  reg        [7:0]    _zz_io_MatrixB_62_33;
  reg        [7:0]    _zz_io_MatrixB_62_34;
  reg        [7:0]    _zz_io_MatrixB_62_35;
  reg        [7:0]    _zz_io_MatrixB_62_36;
  reg        [7:0]    _zz_io_MatrixB_62_37;
  reg        [7:0]    _zz_io_MatrixB_62_38;
  reg        [7:0]    _zz_io_MatrixB_62_39;
  reg        [7:0]    _zz_io_MatrixB_62_40;
  reg        [7:0]    _zz_io_MatrixB_62_41;
  reg        [7:0]    _zz_io_MatrixB_62_42;
  reg        [7:0]    _zz_io_MatrixB_62_43;
  reg        [7:0]    _zz_io_MatrixB_62_44;
  reg        [7:0]    _zz_io_MatrixB_62_45;
  reg        [7:0]    _zz_io_MatrixB_62_46;
  reg        [7:0]    _zz_io_MatrixB_62_47;
  reg        [7:0]    _zz_io_MatrixB_62_48;
  reg        [7:0]    _zz_io_MatrixB_62_49;
  reg        [7:0]    _zz_io_MatrixB_62_50;
  reg        [7:0]    _zz_io_MatrixB_62_51;
  reg        [7:0]    _zz_io_MatrixB_62_52;
  reg        [7:0]    _zz_io_MatrixB_62_53;
  reg        [7:0]    _zz_io_MatrixB_62_54;
  reg        [7:0]    _zz_io_MatrixB_62_55;
  reg        [7:0]    _zz_io_MatrixB_62_56;
  reg        [7:0]    _zz_io_MatrixB_62_57;
  reg        [7:0]    _zz_io_MatrixB_62_58;
  reg        [7:0]    _zz_io_MatrixB_62_59;
  reg        [7:0]    _zz_io_MatrixB_62_60;
  reg        [7:0]    _zz_io_MatrixB_62_61;
  reg                 _zz_io_B_Valid_62;
  reg                 _zz_io_B_Valid_62_1;
  reg                 _zz_io_B_Valid_62_2;
  reg                 _zz_io_B_Valid_62_3;
  reg                 _zz_io_B_Valid_62_4;
  reg                 _zz_io_B_Valid_62_5;
  reg                 _zz_io_B_Valid_62_6;
  reg                 _zz_io_B_Valid_62_7;
  reg                 _zz_io_B_Valid_62_8;
  reg                 _zz_io_B_Valid_62_9;
  reg                 _zz_io_B_Valid_62_10;
  reg                 _zz_io_B_Valid_62_11;
  reg                 _zz_io_B_Valid_62_12;
  reg                 _zz_io_B_Valid_62_13;
  reg                 _zz_io_B_Valid_62_14;
  reg                 _zz_io_B_Valid_62_15;
  reg                 _zz_io_B_Valid_62_16;
  reg                 _zz_io_B_Valid_62_17;
  reg                 _zz_io_B_Valid_62_18;
  reg                 _zz_io_B_Valid_62_19;
  reg                 _zz_io_B_Valid_62_20;
  reg                 _zz_io_B_Valid_62_21;
  reg                 _zz_io_B_Valid_62_22;
  reg                 _zz_io_B_Valid_62_23;
  reg                 _zz_io_B_Valid_62_24;
  reg                 _zz_io_B_Valid_62_25;
  reg                 _zz_io_B_Valid_62_26;
  reg                 _zz_io_B_Valid_62_27;
  reg                 _zz_io_B_Valid_62_28;
  reg                 _zz_io_B_Valid_62_29;
  reg                 _zz_io_B_Valid_62_30;
  reg                 _zz_io_B_Valid_62_31;
  reg                 _zz_io_B_Valid_62_32;
  reg                 _zz_io_B_Valid_62_33;
  reg                 _zz_io_B_Valid_62_34;
  reg                 _zz_io_B_Valid_62_35;
  reg                 _zz_io_B_Valid_62_36;
  reg                 _zz_io_B_Valid_62_37;
  reg                 _zz_io_B_Valid_62_38;
  reg                 _zz_io_B_Valid_62_39;
  reg                 _zz_io_B_Valid_62_40;
  reg                 _zz_io_B_Valid_62_41;
  reg                 _zz_io_B_Valid_62_42;
  reg                 _zz_io_B_Valid_62_43;
  reg                 _zz_io_B_Valid_62_44;
  reg                 _zz_io_B_Valid_62_45;
  reg                 _zz_io_B_Valid_62_46;
  reg                 _zz_io_B_Valid_62_47;
  reg                 _zz_io_B_Valid_62_48;
  reg                 _zz_io_B_Valid_62_49;
  reg                 _zz_io_B_Valid_62_50;
  reg                 _zz_io_B_Valid_62_51;
  reg                 _zz_io_B_Valid_62_52;
  reg                 _zz_io_B_Valid_62_53;
  reg                 _zz_io_B_Valid_62_54;
  reg                 _zz_io_B_Valid_62_55;
  reg                 _zz_io_B_Valid_62_56;
  reg                 _zz_io_B_Valid_62_57;
  reg                 _zz_io_B_Valid_62_58;
  reg                 _zz_io_B_Valid_62_59;
  reg                 _zz_io_B_Valid_62_60;
  reg                 _zz_io_B_Valid_62_61;
  reg        [7:0]    _zz_io_MatrixB_63;
  reg        [7:0]    _zz_io_MatrixB_63_1;
  reg        [7:0]    _zz_io_MatrixB_63_2;
  reg        [7:0]    _zz_io_MatrixB_63_3;
  reg        [7:0]    _zz_io_MatrixB_63_4;
  reg        [7:0]    _zz_io_MatrixB_63_5;
  reg        [7:0]    _zz_io_MatrixB_63_6;
  reg        [7:0]    _zz_io_MatrixB_63_7;
  reg        [7:0]    _zz_io_MatrixB_63_8;
  reg        [7:0]    _zz_io_MatrixB_63_9;
  reg        [7:0]    _zz_io_MatrixB_63_10;
  reg        [7:0]    _zz_io_MatrixB_63_11;
  reg        [7:0]    _zz_io_MatrixB_63_12;
  reg        [7:0]    _zz_io_MatrixB_63_13;
  reg        [7:0]    _zz_io_MatrixB_63_14;
  reg        [7:0]    _zz_io_MatrixB_63_15;
  reg        [7:0]    _zz_io_MatrixB_63_16;
  reg        [7:0]    _zz_io_MatrixB_63_17;
  reg        [7:0]    _zz_io_MatrixB_63_18;
  reg        [7:0]    _zz_io_MatrixB_63_19;
  reg        [7:0]    _zz_io_MatrixB_63_20;
  reg        [7:0]    _zz_io_MatrixB_63_21;
  reg        [7:0]    _zz_io_MatrixB_63_22;
  reg        [7:0]    _zz_io_MatrixB_63_23;
  reg        [7:0]    _zz_io_MatrixB_63_24;
  reg        [7:0]    _zz_io_MatrixB_63_25;
  reg        [7:0]    _zz_io_MatrixB_63_26;
  reg        [7:0]    _zz_io_MatrixB_63_27;
  reg        [7:0]    _zz_io_MatrixB_63_28;
  reg        [7:0]    _zz_io_MatrixB_63_29;
  reg        [7:0]    _zz_io_MatrixB_63_30;
  reg        [7:0]    _zz_io_MatrixB_63_31;
  reg        [7:0]    _zz_io_MatrixB_63_32;
  reg        [7:0]    _zz_io_MatrixB_63_33;
  reg        [7:0]    _zz_io_MatrixB_63_34;
  reg        [7:0]    _zz_io_MatrixB_63_35;
  reg        [7:0]    _zz_io_MatrixB_63_36;
  reg        [7:0]    _zz_io_MatrixB_63_37;
  reg        [7:0]    _zz_io_MatrixB_63_38;
  reg        [7:0]    _zz_io_MatrixB_63_39;
  reg        [7:0]    _zz_io_MatrixB_63_40;
  reg        [7:0]    _zz_io_MatrixB_63_41;
  reg        [7:0]    _zz_io_MatrixB_63_42;
  reg        [7:0]    _zz_io_MatrixB_63_43;
  reg        [7:0]    _zz_io_MatrixB_63_44;
  reg        [7:0]    _zz_io_MatrixB_63_45;
  reg        [7:0]    _zz_io_MatrixB_63_46;
  reg        [7:0]    _zz_io_MatrixB_63_47;
  reg        [7:0]    _zz_io_MatrixB_63_48;
  reg        [7:0]    _zz_io_MatrixB_63_49;
  reg        [7:0]    _zz_io_MatrixB_63_50;
  reg        [7:0]    _zz_io_MatrixB_63_51;
  reg        [7:0]    _zz_io_MatrixB_63_52;
  reg        [7:0]    _zz_io_MatrixB_63_53;
  reg        [7:0]    _zz_io_MatrixB_63_54;
  reg        [7:0]    _zz_io_MatrixB_63_55;
  reg        [7:0]    _zz_io_MatrixB_63_56;
  reg        [7:0]    _zz_io_MatrixB_63_57;
  reg        [7:0]    _zz_io_MatrixB_63_58;
  reg        [7:0]    _zz_io_MatrixB_63_59;
  reg        [7:0]    _zz_io_MatrixB_63_60;
  reg        [7:0]    _zz_io_MatrixB_63_61;
  reg        [7:0]    _zz_io_MatrixB_63_62;
  reg                 _zz_io_B_Valid_63;
  reg                 _zz_io_B_Valid_63_1;
  reg                 _zz_io_B_Valid_63_2;
  reg                 _zz_io_B_Valid_63_3;
  reg                 _zz_io_B_Valid_63_4;
  reg                 _zz_io_B_Valid_63_5;
  reg                 _zz_io_B_Valid_63_6;
  reg                 _zz_io_B_Valid_63_7;
  reg                 _zz_io_B_Valid_63_8;
  reg                 _zz_io_B_Valid_63_9;
  reg                 _zz_io_B_Valid_63_10;
  reg                 _zz_io_B_Valid_63_11;
  reg                 _zz_io_B_Valid_63_12;
  reg                 _zz_io_B_Valid_63_13;
  reg                 _zz_io_B_Valid_63_14;
  reg                 _zz_io_B_Valid_63_15;
  reg                 _zz_io_B_Valid_63_16;
  reg                 _zz_io_B_Valid_63_17;
  reg                 _zz_io_B_Valid_63_18;
  reg                 _zz_io_B_Valid_63_19;
  reg                 _zz_io_B_Valid_63_20;
  reg                 _zz_io_B_Valid_63_21;
  reg                 _zz_io_B_Valid_63_22;
  reg                 _zz_io_B_Valid_63_23;
  reg                 _zz_io_B_Valid_63_24;
  reg                 _zz_io_B_Valid_63_25;
  reg                 _zz_io_B_Valid_63_26;
  reg                 _zz_io_B_Valid_63_27;
  reg                 _zz_io_B_Valid_63_28;
  reg                 _zz_io_B_Valid_63_29;
  reg                 _zz_io_B_Valid_63_30;
  reg                 _zz_io_B_Valid_63_31;
  reg                 _zz_io_B_Valid_63_32;
  reg                 _zz_io_B_Valid_63_33;
  reg                 _zz_io_B_Valid_63_34;
  reg                 _zz_io_B_Valid_63_35;
  reg                 _zz_io_B_Valid_63_36;
  reg                 _zz_io_B_Valid_63_37;
  reg                 _zz_io_B_Valid_63_38;
  reg                 _zz_io_B_Valid_63_39;
  reg                 _zz_io_B_Valid_63_40;
  reg                 _zz_io_B_Valid_63_41;
  reg                 _zz_io_B_Valid_63_42;
  reg                 _zz_io_B_Valid_63_43;
  reg                 _zz_io_B_Valid_63_44;
  reg                 _zz_io_B_Valid_63_45;
  reg                 _zz_io_B_Valid_63_46;
  reg                 _zz_io_B_Valid_63_47;
  reg                 _zz_io_B_Valid_63_48;
  reg                 _zz_io_B_Valid_63_49;
  reg                 _zz_io_B_Valid_63_50;
  reg                 _zz_io_B_Valid_63_51;
  reg                 _zz_io_B_Valid_63_52;
  reg                 _zz_io_B_Valid_63_53;
  reg                 _zz_io_B_Valid_63_54;
  reg                 _zz_io_B_Valid_63_55;
  reg                 _zz_io_B_Valid_63_56;
  reg                 _zz_io_B_Valid_63_57;
  reg                 _zz_io_B_Valid_63_58;
  reg                 _zz_io_B_Valid_63_59;
  reg                 _zz_io_B_Valid_63_60;
  reg                 _zz_io_B_Valid_63_61;
  reg                 _zz_io_B_Valid_63_62;
  reg                 toplevel_SubModule_WeightCache_Weight_Cached_delay_1;
  reg                 toplevel_SubModule_WeightCache_Weight_Cached_delay_2;
  reg                 toplevel_SubModule_WeightCache_Weight_Cached_delay_3;
  reg                 _zz_start;
  reg                 _zz_start_1;
  reg                 _zz_start_2;
  `ifndef SYNTHESIS
  reg [127:0] Fsm_currentState_string;
  reg [127:0] Fsm_nextState_string;
  `endif


  Compute_DataIn_Switch InputSwitch (
    .Switch               (InputSwitch_Switch[1:0]              ), //i
    .s0_axis_s2mm_tdata   (s_axis_s2mm_tdata[63:0]              ), //i
    .s0_axis_s2mm_tkeep   (s_axis_s2mm_tkeep[7:0]               ), //i
    .s0_axis_s2mm_tlast   (s_axis_s2mm_tlast                    ), //i
    .s0_axis_s2mm_tready  (InputSwitch_s0_axis_s2mm_tready      ), //o
    .s0_axis_s2mm_tvalid  (s_axis_s2mm_tvalid                   ), //i
    .m_0_axis_mm2s_tdata  (InputSwitch_m_0_axis_mm2s_tdata[63:0]), //o
    .m_0_axis_mm2s_tkeep  (InputSwitch_m_0_axis_mm2s_tkeep[7:0] ), //o
    .m_0_axis_mm2s_tlast  (InputSwitch_m_0_axis_mm2s_tlast      ), //o
    .m_0_axis_mm2s_tready (InputSwitch_m_0_axis_mm2s_tready     ), //i
    .m_0_axis_mm2s_tvalid (InputSwitch_m_0_axis_mm2s_tvalid     ), //o
    .m_1_axis_mm2s_tdata  (InputSwitch_m_1_axis_mm2s_tdata[63:0]), //o
    .m_1_axis_mm2s_tkeep  (InputSwitch_m_1_axis_mm2s_tkeep[7:0] ), //o
    .m_1_axis_mm2s_tlast  (InputSwitch_m_1_axis_mm2s_tlast      ), //o
    .m_1_axis_mm2s_tready (SubModule_Img2Col_s_axis_s2mm_tready ), //i
    .m_1_axis_mm2s_tvalid (InputSwitch_m_1_axis_mm2s_tvalid     )  //o
  );
  Img2ColStreamV2 SubModule_Img2Col (
    .mData                          (SubModule_Img2Col_mData[63:0]               ), //o
    .mValid                         (SubModule_Img2Col_mValid[7:0]               ), //o
    .s_axis_s2mm_tdata              (InputSwitch_m_1_axis_mm2s_tdata[63:0]       ), //i
    .s_axis_s2mm_tkeep              (InputSwitch_m_1_axis_mm2s_tkeep[7:0]        ), //i
    .s_axis_s2mm_tlast              (InputSwitch_m_1_axis_mm2s_tlast             ), //i
    .s_axis_s2mm_tready             (SubModule_Img2Col_s_axis_s2mm_tready        ), //o
    .s_axis_s2mm_tvalid             (InputSwitch_m_1_axis_mm2s_tvalid            ), //i
    .start                          (SubModule_Img2Col_start                     ), //i
    .Raddr_Valid                    (SubModule_Img2Col_Raddr_Valid               ), //o
    .LayerEnd                       (SubModule_Img2Col_LayerEnd                  ), //o
    .Stride                         (Img2Col_Stride[4:0]                         ), //i
    .Kernel_Size                    (Img2Col_Kernel_Size[4:0]                    ), //i
    .Window_Size                    (Img2Col_Window_Size[15:0]                   ), //i
    .InFeature_Size                 (Img2Col_InFeature_Size[15:0]                ), //i
    .InFeature_Channel              (Img2Col_InFeature_Channel[15:0]             ), //i
    .OutFeature_Channel             (Img2Col_OutFeature_Channel[15:0]            ), //i
    .OutFeature_Size                (Img2Col_OutFeature_Size[15:0]               ), //i
    .OutCol_Count_Times             (Img2Col_OutCol_Count_Times[15:0]            ), //i
    .InCol_Count_Times              (Img2Col_InCol_Count_Times[15:0]             ), //i
    .OutRow_Count_Times             (Img2Col_OutRow_Count_Times[15:0]            ), //i
    .OutFeature_Channel_Count_Times (Img2Col_OutFeature_Channel_Count_Times[15:0]), //i
    .Sliding_Size                   (Img2Col_Sliding_Size[12:0]                  ), //i
    .clk                            (clk                                         ), //i
    .reset                          (reset                                       )  //i
  );
  SA_3D SubModule_SA_3D (
    .start              (Control_start                           ), //i
    ._zz_io_MatrixA_0   (SubModule_SA_3D__zz_io_MatrixA_0[7:0]   ), //i
    ._zz_io_MatrixA_1   (SubModule_SA_3D__zz_io_MatrixA_1[7:0]   ), //i
    ._zz_io_MatrixA_2   (SubModule_SA_3D__zz_io_MatrixA_2[7:0]   ), //i
    ._zz_io_MatrixA_3   (SubModule_SA_3D__zz_io_MatrixA_3[7:0]   ), //i
    ._zz_io_MatrixA_4   (SubModule_SA_3D__zz_io_MatrixA_4[7:0]   ), //i
    ._zz_io_MatrixA_5   (SubModule_SA_3D__zz_io_MatrixA_5[7:0]   ), //i
    ._zz_io_MatrixA_6   (SubModule_SA_3D__zz_io_MatrixA_6[7:0]   ), //i
    ._zz_io_MatrixA_7   (SubModule_SA_3D__zz_io_MatrixA_7[7:0]   ), //i
    ._zz_io_MatrixB_0   (SubModule_SA_3D__zz_io_MatrixB_0[7:0]   ), //i
    ._zz_io_MatrixB_1   (_zz_io_MatrixB_1[7:0]                   ), //i
    ._zz_io_MatrixB_2   (_zz_io_MatrixB_2_1[7:0]                 ), //i
    ._zz_io_MatrixB_3   (_zz_io_MatrixB_3_2[7:0]                 ), //i
    ._zz_io_MatrixB_4   (_zz_io_MatrixB_4_3[7:0]                 ), //i
    ._zz_io_MatrixB_5   (_zz_io_MatrixB_5_4[7:0]                 ), //i
    ._zz_io_MatrixB_6   (_zz_io_MatrixB_6_5[7:0]                 ), //i
    ._zz_io_MatrixB_7   (_zz_io_MatrixB_7_6[7:0]                 ), //i
    ._zz_io_MatrixB_8   (_zz_io_MatrixB_8_7[7:0]                 ), //i
    ._zz_io_MatrixB_9   (_zz_io_MatrixB_9_8[7:0]                 ), //i
    ._zz_io_MatrixB_10  (_zz_io_MatrixB_10_9[7:0]                ), //i
    ._zz_io_MatrixB_11  (_zz_io_MatrixB_11_10[7:0]               ), //i
    ._zz_io_MatrixB_12  (_zz_io_MatrixB_12_11[7:0]               ), //i
    ._zz_io_MatrixB_13  (_zz_io_MatrixB_13_12[7:0]               ), //i
    ._zz_io_MatrixB_14  (_zz_io_MatrixB_14_13[7:0]               ), //i
    ._zz_io_MatrixB_15  (_zz_io_MatrixB_15_14[7:0]               ), //i
    ._zz_io_MatrixB_16  (_zz_io_MatrixB_16_15[7:0]               ), //i
    ._zz_io_MatrixB_17  (_zz_io_MatrixB_17_16[7:0]               ), //i
    ._zz_io_MatrixB_18  (_zz_io_MatrixB_18_17[7:0]               ), //i
    ._zz_io_MatrixB_19  (_zz_io_MatrixB_19_18[7:0]               ), //i
    ._zz_io_MatrixB_20  (_zz_io_MatrixB_20_19[7:0]               ), //i
    ._zz_io_MatrixB_21  (_zz_io_MatrixB_21_20[7:0]               ), //i
    ._zz_io_MatrixB_22  (_zz_io_MatrixB_22_21[7:0]               ), //i
    ._zz_io_MatrixB_23  (_zz_io_MatrixB_23_22[7:0]               ), //i
    ._zz_io_MatrixB_24  (_zz_io_MatrixB_24_23[7:0]               ), //i
    ._zz_io_MatrixB_25  (_zz_io_MatrixB_25_24[7:0]               ), //i
    ._zz_io_MatrixB_26  (_zz_io_MatrixB_26_25[7:0]               ), //i
    ._zz_io_MatrixB_27  (_zz_io_MatrixB_27_26[7:0]               ), //i
    ._zz_io_MatrixB_28  (_zz_io_MatrixB_28_27[7:0]               ), //i
    ._zz_io_MatrixB_29  (_zz_io_MatrixB_29_28[7:0]               ), //i
    ._zz_io_MatrixB_30  (_zz_io_MatrixB_30_29[7:0]               ), //i
    ._zz_io_MatrixB_31  (_zz_io_MatrixB_31_30[7:0]               ), //i
    ._zz_io_MatrixB_32  (_zz_io_MatrixB_32_31[7:0]               ), //i
    ._zz_io_MatrixB_33  (_zz_io_MatrixB_33_32[7:0]               ), //i
    ._zz_io_MatrixB_34  (_zz_io_MatrixB_34_33[7:0]               ), //i
    ._zz_io_MatrixB_35  (_zz_io_MatrixB_35_34[7:0]               ), //i
    ._zz_io_MatrixB_36  (_zz_io_MatrixB_36_35[7:0]               ), //i
    ._zz_io_MatrixB_37  (_zz_io_MatrixB_37_36[7:0]               ), //i
    ._zz_io_MatrixB_38  (_zz_io_MatrixB_38_37[7:0]               ), //i
    ._zz_io_MatrixB_39  (_zz_io_MatrixB_39_38[7:0]               ), //i
    ._zz_io_MatrixB_40  (_zz_io_MatrixB_40_39[7:0]               ), //i
    ._zz_io_MatrixB_41  (_zz_io_MatrixB_41_40[7:0]               ), //i
    ._zz_io_MatrixB_42  (_zz_io_MatrixB_42_41[7:0]               ), //i
    ._zz_io_MatrixB_43  (_zz_io_MatrixB_43_42[7:0]               ), //i
    ._zz_io_MatrixB_44  (_zz_io_MatrixB_44_43[7:0]               ), //i
    ._zz_io_MatrixB_45  (_zz_io_MatrixB_45_44[7:0]               ), //i
    ._zz_io_MatrixB_46  (_zz_io_MatrixB_46_45[7:0]               ), //i
    ._zz_io_MatrixB_47  (_zz_io_MatrixB_47_46[7:0]               ), //i
    ._zz_io_MatrixB_48  (_zz_io_MatrixB_48_47[7:0]               ), //i
    ._zz_io_MatrixB_49  (_zz_io_MatrixB_49_48[7:0]               ), //i
    ._zz_io_MatrixB_50  (_zz_io_MatrixB_50_49[7:0]               ), //i
    ._zz_io_MatrixB_51  (_zz_io_MatrixB_51_50[7:0]               ), //i
    ._zz_io_MatrixB_52  (_zz_io_MatrixB_52_51[7:0]               ), //i
    ._zz_io_MatrixB_53  (_zz_io_MatrixB_53_52[7:0]               ), //i
    ._zz_io_MatrixB_54  (_zz_io_MatrixB_54_53[7:0]               ), //i
    ._zz_io_MatrixB_55  (_zz_io_MatrixB_55_54[7:0]               ), //i
    ._zz_io_MatrixB_56  (_zz_io_MatrixB_56_55[7:0]               ), //i
    ._zz_io_MatrixB_57  (_zz_io_MatrixB_57_56[7:0]               ), //i
    ._zz_io_MatrixB_58  (_zz_io_MatrixB_58_57[7:0]               ), //i
    ._zz_io_MatrixB_59  (_zz_io_MatrixB_59_58[7:0]               ), //i
    ._zz_io_MatrixB_60  (_zz_io_MatrixB_60_59[7:0]               ), //i
    ._zz_io_MatrixB_61  (_zz_io_MatrixB_61_60[7:0]               ), //i
    ._zz_io_MatrixB_62  (_zz_io_MatrixB_62_61[7:0]               ), //i
    ._zz_io_MatrixB_63  (_zz_io_MatrixB_63_62[7:0]               ), //i
    ._zz_io_A_Valid_0   (SubModule_SA_3D__zz_io_A_Valid_0        ), //i
    ._zz_io_A_Valid_1   (SubModule_SA_3D__zz_io_A_Valid_1        ), //i
    ._zz_io_A_Valid_2   (SubModule_SA_3D__zz_io_A_Valid_2        ), //i
    ._zz_io_A_Valid_3   (SubModule_SA_3D__zz_io_A_Valid_3        ), //i
    ._zz_io_A_Valid_4   (SubModule_SA_3D__zz_io_A_Valid_4        ), //i
    ._zz_io_A_Valid_5   (SubModule_SA_3D__zz_io_A_Valid_5        ), //i
    ._zz_io_A_Valid_6   (SubModule_SA_3D__zz_io_A_Valid_6        ), //i
    ._zz_io_A_Valid_7   (SubModule_SA_3D__zz_io_A_Valid_7        ), //i
    ._zz_io_B_Valid_0   (SubModule_SA_3D__zz_io_B_Valid_0        ), //i
    ._zz_io_B_Valid_1   (_zz_io_B_Valid_1                        ), //i
    ._zz_io_B_Valid_2   (_zz_io_B_Valid_2_1                      ), //i
    ._zz_io_B_Valid_3   (_zz_io_B_Valid_3_2                      ), //i
    ._zz_io_B_Valid_4   (_zz_io_B_Valid_4_3                      ), //i
    ._zz_io_B_Valid_5   (_zz_io_B_Valid_5_4                      ), //i
    ._zz_io_B_Valid_6   (_zz_io_B_Valid_6_5                      ), //i
    ._zz_io_B_Valid_7   (_zz_io_B_Valid_7_6                      ), //i
    ._zz_io_B_Valid_8   (_zz_io_B_Valid_8_7                      ), //i
    ._zz_io_B_Valid_9   (_zz_io_B_Valid_9_8                      ), //i
    ._zz_io_B_Valid_10  (_zz_io_B_Valid_10_9                     ), //i
    ._zz_io_B_Valid_11  (_zz_io_B_Valid_11_10                    ), //i
    ._zz_io_B_Valid_12  (_zz_io_B_Valid_12_11                    ), //i
    ._zz_io_B_Valid_13  (_zz_io_B_Valid_13_12                    ), //i
    ._zz_io_B_Valid_14  (_zz_io_B_Valid_14_13                    ), //i
    ._zz_io_B_Valid_15  (_zz_io_B_Valid_15_14                    ), //i
    ._zz_io_B_Valid_16  (_zz_io_B_Valid_16_15                    ), //i
    ._zz_io_B_Valid_17  (_zz_io_B_Valid_17_16                    ), //i
    ._zz_io_B_Valid_18  (_zz_io_B_Valid_18_17                    ), //i
    ._zz_io_B_Valid_19  (_zz_io_B_Valid_19_18                    ), //i
    ._zz_io_B_Valid_20  (_zz_io_B_Valid_20_19                    ), //i
    ._zz_io_B_Valid_21  (_zz_io_B_Valid_21_20                    ), //i
    ._zz_io_B_Valid_22  (_zz_io_B_Valid_22_21                    ), //i
    ._zz_io_B_Valid_23  (_zz_io_B_Valid_23_22                    ), //i
    ._zz_io_B_Valid_24  (_zz_io_B_Valid_24_23                    ), //i
    ._zz_io_B_Valid_25  (_zz_io_B_Valid_25_24                    ), //i
    ._zz_io_B_Valid_26  (_zz_io_B_Valid_26_25                    ), //i
    ._zz_io_B_Valid_27  (_zz_io_B_Valid_27_26                    ), //i
    ._zz_io_B_Valid_28  (_zz_io_B_Valid_28_27                    ), //i
    ._zz_io_B_Valid_29  (_zz_io_B_Valid_29_28                    ), //i
    ._zz_io_B_Valid_30  (_zz_io_B_Valid_30_29                    ), //i
    ._zz_io_B_Valid_31  (_zz_io_B_Valid_31_30                    ), //i
    ._zz_io_B_Valid_32  (_zz_io_B_Valid_32_31                    ), //i
    ._zz_io_B_Valid_33  (_zz_io_B_Valid_33_32                    ), //i
    ._zz_io_B_Valid_34  (_zz_io_B_Valid_34_33                    ), //i
    ._zz_io_B_Valid_35  (_zz_io_B_Valid_35_34                    ), //i
    ._zz_io_B_Valid_36  (_zz_io_B_Valid_36_35                    ), //i
    ._zz_io_B_Valid_37  (_zz_io_B_Valid_37_36                    ), //i
    ._zz_io_B_Valid_38  (_zz_io_B_Valid_38_37                    ), //i
    ._zz_io_B_Valid_39  (_zz_io_B_Valid_39_38                    ), //i
    ._zz_io_B_Valid_40  (_zz_io_B_Valid_40_39                    ), //i
    ._zz_io_B_Valid_41  (_zz_io_B_Valid_41_40                    ), //i
    ._zz_io_B_Valid_42  (_zz_io_B_Valid_42_41                    ), //i
    ._zz_io_B_Valid_43  (_zz_io_B_Valid_43_42                    ), //i
    ._zz_io_B_Valid_44  (_zz_io_B_Valid_44_43                    ), //i
    ._zz_io_B_Valid_45  (_zz_io_B_Valid_45_44                    ), //i
    ._zz_io_B_Valid_46  (_zz_io_B_Valid_46_45                    ), //i
    ._zz_io_B_Valid_47  (_zz_io_B_Valid_47_46                    ), //i
    ._zz_io_B_Valid_48  (_zz_io_B_Valid_48_47                    ), //i
    ._zz_io_B_Valid_49  (_zz_io_B_Valid_49_48                    ), //i
    ._zz_io_B_Valid_50  (_zz_io_B_Valid_50_49                    ), //i
    ._zz_io_B_Valid_51  (_zz_io_B_Valid_51_50                    ), //i
    ._zz_io_B_Valid_52  (_zz_io_B_Valid_52_51                    ), //i
    ._zz_io_B_Valid_53  (_zz_io_B_Valid_53_52                    ), //i
    ._zz_io_B_Valid_54  (_zz_io_B_Valid_54_53                    ), //i
    ._zz_io_B_Valid_55  (_zz_io_B_Valid_55_54                    ), //i
    ._zz_io_B_Valid_56  (_zz_io_B_Valid_56_55                    ), //i
    ._zz_io_B_Valid_57  (_zz_io_B_Valid_57_56                    ), //i
    ._zz_io_B_Valid_58  (_zz_io_B_Valid_58_57                    ), //i
    ._zz_io_B_Valid_59  (_zz_io_B_Valid_59_58                    ), //i
    ._zz_io_B_Valid_60  (_zz_io_B_Valid_60_59                    ), //i
    ._zz_io_B_Valid_61  (_zz_io_B_Valid_61_60                    ), //i
    ._zz_io_B_Valid_62  (_zz_io_B_Valid_62_61                    ), //i
    ._zz_io_B_Valid_63  (_zz_io_B_Valid_63_62                    ), //i
    ._zz_io_signCount   (SubModule_SA_3D__zz_io_signCount[15:0]  ), //i
    .clk                (clk                                     ), //i
    .Matrix_C_valid_0   (SubModule_SA_3D_Matrix_C_valid_0        ), //o
    .Matrix_C_valid_1   (SubModule_SA_3D_Matrix_C_valid_1        ), //o
    .Matrix_C_valid_2   (SubModule_SA_3D_Matrix_C_valid_2        ), //o
    .Matrix_C_valid_3   (SubModule_SA_3D_Matrix_C_valid_3        ), //o
    .Matrix_C_valid_4   (SubModule_SA_3D_Matrix_C_valid_4        ), //o
    .Matrix_C_valid_5   (SubModule_SA_3D_Matrix_C_valid_5        ), //o
    .Matrix_C_valid_6   (SubModule_SA_3D_Matrix_C_valid_6        ), //o
    .Matrix_C_valid_7   (SubModule_SA_3D_Matrix_C_valid_7        ), //o
    .Matrix_C_payload_0 (SubModule_SA_3D_Matrix_C_payload_0[31:0]), //o
    .Matrix_C_payload_1 (SubModule_SA_3D_Matrix_C_payload_1[31:0]), //o
    .Matrix_C_payload_2 (SubModule_SA_3D_Matrix_C_payload_2[31:0]), //o
    .Matrix_C_payload_3 (SubModule_SA_3D_Matrix_C_payload_3[31:0]), //o
    .Matrix_C_payload_4 (SubModule_SA_3D_Matrix_C_payload_4[31:0]), //o
    .Matrix_C_payload_5 (SubModule_SA_3D_Matrix_C_payload_5[31:0]), //o
    .Matrix_C_payload_6 (SubModule_SA_3D_Matrix_C_payload_6[31:0]), //o
    .Matrix_C_payload_7 (SubModule_SA_3D_Matrix_C_payload_7[31:0]), //o
    .reset              (reset                                   )  //i
  );
  WeightCache_Stream SubModule_WeightCache (
    .s_axis_s2mm_tdata  (InputSwitch_m_0_axis_mm2s_tdata[63:0]       ), //i
    .s_axis_s2mm_tkeep  (InputSwitch_m_0_axis_mm2s_tkeep[7:0]        ), //i
    .s_axis_s2mm_tlast  (InputSwitch_m_0_axis_mm2s_tlast             ), //i
    .s_axis_s2mm_tready (SubModule_WeightCache_s_axis_s2mm_tready    ), //o
    .s_axis_s2mm_tvalid (InputSwitch_m_0_axis_mm2s_tvalid            ), //i
    .start              (_zz_start_2                                 ), //i
    .Matrix_Row         (Img2Col_WeightMatrix_Row[15:0]              ), //i
    .Matrix_Col         (Img2Col_OutFeature_Channel[15:0]            ), //i
    .mData_0            (SubModule_WeightCache_mData_0[7:0]          ), //o
    .mData_1            (SubModule_WeightCache_mData_1[7:0]          ), //o
    .mData_2            (SubModule_WeightCache_mData_2[7:0]          ), //o
    .mData_3            (SubModule_WeightCache_mData_3[7:0]          ), //o
    .mData_4            (SubModule_WeightCache_mData_4[7:0]          ), //o
    .mData_5            (SubModule_WeightCache_mData_5[7:0]          ), //o
    .mData_6            (SubModule_WeightCache_mData_6[7:0]          ), //o
    .mData_7            (SubModule_WeightCache_mData_7[7:0]          ), //o
    .mData_8            (SubModule_WeightCache_mData_8[7:0]          ), //o
    .mData_9            (SubModule_WeightCache_mData_9[7:0]          ), //o
    .mData_10           (SubModule_WeightCache_mData_10[7:0]         ), //o
    .mData_11           (SubModule_WeightCache_mData_11[7:0]         ), //o
    .mData_12           (SubModule_WeightCache_mData_12[7:0]         ), //o
    .mData_13           (SubModule_WeightCache_mData_13[7:0]         ), //o
    .mData_14           (SubModule_WeightCache_mData_14[7:0]         ), //o
    .mData_15           (SubModule_WeightCache_mData_15[7:0]         ), //o
    .mData_16           (SubModule_WeightCache_mData_16[7:0]         ), //o
    .mData_17           (SubModule_WeightCache_mData_17[7:0]         ), //o
    .mData_18           (SubModule_WeightCache_mData_18[7:0]         ), //o
    .mData_19           (SubModule_WeightCache_mData_19[7:0]         ), //o
    .mData_20           (SubModule_WeightCache_mData_20[7:0]         ), //o
    .mData_21           (SubModule_WeightCache_mData_21[7:0]         ), //o
    .mData_22           (SubModule_WeightCache_mData_22[7:0]         ), //o
    .mData_23           (SubModule_WeightCache_mData_23[7:0]         ), //o
    .mData_24           (SubModule_WeightCache_mData_24[7:0]         ), //o
    .mData_25           (SubModule_WeightCache_mData_25[7:0]         ), //o
    .mData_26           (SubModule_WeightCache_mData_26[7:0]         ), //o
    .mData_27           (SubModule_WeightCache_mData_27[7:0]         ), //o
    .mData_28           (SubModule_WeightCache_mData_28[7:0]         ), //o
    .mData_29           (SubModule_WeightCache_mData_29[7:0]         ), //o
    .mData_30           (SubModule_WeightCache_mData_30[7:0]         ), //o
    .mData_31           (SubModule_WeightCache_mData_31[7:0]         ), //o
    .mData_32           (SubModule_WeightCache_mData_32[7:0]         ), //o
    .mData_33           (SubModule_WeightCache_mData_33[7:0]         ), //o
    .mData_34           (SubModule_WeightCache_mData_34[7:0]         ), //o
    .mData_35           (SubModule_WeightCache_mData_35[7:0]         ), //o
    .mData_36           (SubModule_WeightCache_mData_36[7:0]         ), //o
    .mData_37           (SubModule_WeightCache_mData_37[7:0]         ), //o
    .mData_38           (SubModule_WeightCache_mData_38[7:0]         ), //o
    .mData_39           (SubModule_WeightCache_mData_39[7:0]         ), //o
    .mData_40           (SubModule_WeightCache_mData_40[7:0]         ), //o
    .mData_41           (SubModule_WeightCache_mData_41[7:0]         ), //o
    .mData_42           (SubModule_WeightCache_mData_42[7:0]         ), //o
    .mData_43           (SubModule_WeightCache_mData_43[7:0]         ), //o
    .mData_44           (SubModule_WeightCache_mData_44[7:0]         ), //o
    .mData_45           (SubModule_WeightCache_mData_45[7:0]         ), //o
    .mData_46           (SubModule_WeightCache_mData_46[7:0]         ), //o
    .mData_47           (SubModule_WeightCache_mData_47[7:0]         ), //o
    .mData_48           (SubModule_WeightCache_mData_48[7:0]         ), //o
    .mData_49           (SubModule_WeightCache_mData_49[7:0]         ), //o
    .mData_50           (SubModule_WeightCache_mData_50[7:0]         ), //o
    .mData_51           (SubModule_WeightCache_mData_51[7:0]         ), //o
    .mData_52           (SubModule_WeightCache_mData_52[7:0]         ), //o
    .mData_53           (SubModule_WeightCache_mData_53[7:0]         ), //o
    .mData_54           (SubModule_WeightCache_mData_54[7:0]         ), //o
    .mData_55           (SubModule_WeightCache_mData_55[7:0]         ), //o
    .mData_56           (SubModule_WeightCache_mData_56[7:0]         ), //o
    .mData_57           (SubModule_WeightCache_mData_57[7:0]         ), //o
    .mData_58           (SubModule_WeightCache_mData_58[7:0]         ), //o
    .mData_59           (SubModule_WeightCache_mData_59[7:0]         ), //o
    .mData_60           (SubModule_WeightCache_mData_60[7:0]         ), //o
    .mData_61           (SubModule_WeightCache_mData_61[7:0]         ), //o
    .mData_62           (SubModule_WeightCache_mData_62[7:0]         ), //o
    .mData_63           (SubModule_WeightCache_mData_63[7:0]         ), //o
    .Raddr_Valid        (SubModule_Img2Col_Raddr_Valid               ), //i
    .Weight_Cached      (SubModule_WeightCache_Weight_Cached         ), //o
    .LayerEnd           (LayerEnd                                    ), //i
    .MatrixCol_Switch   (SubModule_WeightCache_MatrixCol_Switch[63:0]), //o
    .clk                (clk                                         ), //i
    .reset              (reset                                       )  //i
  );
  ConvArrangeV3 SubModule_DataArrange (
    .sData_0        (SubModule_DataArrange_sData_0[7:0]       ), //i
    .sData_1        (SubModule_DataArrange_sData_1[7:0]       ), //i
    .sData_2        (SubModule_DataArrange_sData_2[7:0]       ), //i
    .sData_3        (SubModule_DataArrange_sData_3[7:0]       ), //i
    .sData_4        (SubModule_DataArrange_sData_4[7:0]       ), //i
    .sData_5        (SubModule_DataArrange_sData_5[7:0]       ), //i
    .sData_6        (SubModule_DataArrange_sData_6[7:0]       ), //i
    .sData_7        (SubModule_DataArrange_sData_7[7:0]       ), //i
    .sReady         (SubModule_DataArrange_sReady             ), //o
    .sValid         (SubModule_DataArrange_sValid[7:0]        ), //i
    .MatrixCol      (Img2Col_OutMatrix_Col[11:0]              ), //i
    .MatrixRow      (Img2Col_OutMatrix_Row[19:0]              ), //i
    .OutChannel     (SubModule_DataArrange_OutChannel[9:0]    ), //i
    .OutFeatureSize (Img2Col_OutFeature_Size[15:0]            ), //i
    .mData_valid    (SubModule_DataArrange_mData_valid        ), //o
    .mData_ready    (m_axis_mm2s_tready                       ), //i
    .mData_payload  (SubModule_DataArrange_mData_payload[63:0]), //o
    .mLast          (SubModule_DataArrange_mLast              ), //o
    .LayerEnd       (SubModule_DataArrange_LayerEnd           ), //o
    .start          (Control_start                            ), //i
    .SwitchConv     (Control_Switch_Conv                      ), //i
    .clk            (clk                                      ), //i
    .reset          (reset                                    )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      TopCtrl_Enum_IDLE : Fsm_currentState_string = "IDLE            ";
      TopCtrl_Enum_INIT : Fsm_currentState_string = "INIT            ";
      TopCtrl_Enum_WEIGHT_CACHE : Fsm_currentState_string = "WEIGHT_CACHE    ";
      TopCtrl_Enum_RECEIVE_PICTURE : Fsm_currentState_string = "RECEIVE_PICTURE ";
      TopCtrl_Enum_RECEIVE_MATRIX : Fsm_currentState_string = "RECEIVE_MATRIX  ";
      TopCtrl_Enum_WAIT_COMPUTE_END : Fsm_currentState_string = "WAIT_COMPUTE_END";
      default : Fsm_currentState_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      TopCtrl_Enum_IDLE : Fsm_nextState_string = "IDLE            ";
      TopCtrl_Enum_INIT : Fsm_nextState_string = "INIT            ";
      TopCtrl_Enum_WEIGHT_CACHE : Fsm_nextState_string = "WEIGHT_CACHE    ";
      TopCtrl_Enum_RECEIVE_PICTURE : Fsm_nextState_string = "RECEIVE_PICTURE ";
      TopCtrl_Enum_RECEIVE_MATRIX : Fsm_nextState_string = "RECEIVE_MATRIX  ";
      TopCtrl_Enum_WAIT_COMPUTE_END : Fsm_nextState_string = "WAIT_COMPUTE_END";
      default : Fsm_nextState_string = "????????????????";
    endcase
  end
  `endif

  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & TopCtrl_Enum_IDLE) == TopCtrl_Enum_IDLE) : begin
        if(Control_start) begin
          Fsm_nextState = TopCtrl_Enum_INIT;
        end else begin
          Fsm_nextState = TopCtrl_Enum_IDLE;
        end
      end
      (((Fsm_currentState) & TopCtrl_Enum_INIT) == TopCtrl_Enum_INIT) : begin
        if(Fsm_Inited) begin
          Fsm_nextState = TopCtrl_Enum_WEIGHT_CACHE;
        end else begin
          Fsm_nextState = TopCtrl_Enum_INIT;
        end
      end
      (((Fsm_currentState) & TopCtrl_Enum_WEIGHT_CACHE) == TopCtrl_Enum_WEIGHT_CACHE) : begin
        if(when_SA3D_Top_l46) begin
          Fsm_nextState = TopCtrl_Enum_RECEIVE_PICTURE;
        end else begin
          if(when_SA3D_Top_l48) begin
            Fsm_nextState = TopCtrl_Enum_RECEIVE_MATRIX;
          end else begin
            Fsm_nextState = TopCtrl_Enum_WEIGHT_CACHE;
          end
        end
      end
      (((Fsm_currentState) & TopCtrl_Enum_RECEIVE_PICTURE) == TopCtrl_Enum_RECEIVE_PICTURE) : begin
        if(Fsm_Picture_Received) begin
          Fsm_nextState = TopCtrl_Enum_WAIT_COMPUTE_END;
        end else begin
          Fsm_nextState = TopCtrl_Enum_RECEIVE_PICTURE;
        end
      end
      (((Fsm_currentState) & TopCtrl_Enum_RECEIVE_MATRIX) == TopCtrl_Enum_RECEIVE_MATRIX) : begin
        if(Fsm_Matrix_Received) begin
          Fsm_nextState = TopCtrl_Enum_WAIT_COMPUTE_END;
        end else begin
          Fsm_nextState = TopCtrl_Enum_RECEIVE_MATRIX;
        end
      end
      default : begin
        if(Fsm_Compute_End) begin
          Fsm_nextState = TopCtrl_Enum_IDLE;
        end else begin
          Fsm_nextState = TopCtrl_Enum_WAIT_COMPUTE_END;
        end
      end
    endcase
  end

  assign when_SA3D_Top_l46 = (Fsm_WeightCached && Fsm_Switch_Conv);
  assign when_SA3D_Top_l48 = (Fsm_WeightCached && (! Fsm_Switch_Conv));
  assign Fsm_Compute_End = LayerEnd;
  assign when_WaCounter_l19 = ((Fsm_currentState & TopCtrl_Enum_INIT) != 6'b000000);
  assign when_WaCounter_l14 = (InitCnt_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l14) begin
      InitCnt_valid = 1'b1;
    end else begin
      InitCnt_valid = 1'b0;
    end
  end

  assign Fsm_Inited = InitCnt_valid;
  assign s_axis_s2mm_tready = InputSwitch_s0_axis_s2mm_tready;
  assign when_SA3D_Top_l131 = ((Fsm_currentState & TopCtrl_Enum_WEIGHT_CACHE) != 6'b000000);
  always @(*) begin
    if(when_SA3D_Top_l131) begin
      InputSwitch_Switch = 2'b00;
    end else begin
      if(Control_Switch_Conv) begin
        InputSwitch_Switch = 2'b01;
      end else begin
        InputSwitch_Switch = 2'b10;
      end
    end
  end

  assign SubModule_SA_3D__zz_io_MatrixA_0 = SubModule_Img2Col_mData[7 : 0];
  assign SubModule_SA_3D__zz_io_A_Valid_0 = SubModule_Img2Col_mValid[0];
  assign SubModule_SA_3D__zz_io_MatrixA_1 = SubModule_Img2Col_mData[15 : 8];
  assign SubModule_SA_3D__zz_io_A_Valid_1 = SubModule_Img2Col_mValid[1];
  assign SubModule_SA_3D__zz_io_MatrixA_2 = SubModule_Img2Col_mData[23 : 16];
  assign SubModule_SA_3D__zz_io_A_Valid_2 = SubModule_Img2Col_mValid[2];
  assign SubModule_SA_3D__zz_io_MatrixA_3 = SubModule_Img2Col_mData[31 : 24];
  assign SubModule_SA_3D__zz_io_A_Valid_3 = SubModule_Img2Col_mValid[3];
  assign SubModule_SA_3D__zz_io_MatrixA_4 = SubModule_Img2Col_mData[39 : 32];
  assign SubModule_SA_3D__zz_io_A_Valid_4 = SubModule_Img2Col_mValid[4];
  assign SubModule_SA_3D__zz_io_MatrixA_5 = SubModule_Img2Col_mData[47 : 40];
  assign SubModule_SA_3D__zz_io_A_Valid_5 = SubModule_Img2Col_mValid[5];
  assign SubModule_SA_3D__zz_io_MatrixA_6 = SubModule_Img2Col_mData[55 : 48];
  assign SubModule_SA_3D__zz_io_A_Valid_6 = SubModule_Img2Col_mValid[6];
  assign SubModule_SA_3D__zz_io_MatrixA_7 = SubModule_Img2Col_mData[63 : 56];
  assign SubModule_SA_3D__zz_io_A_Valid_7 = SubModule_Img2Col_mValid[7];
  assign SubModule_SA_3D__zz_io_signCount = (Img2Col_WeightMatrix_Row - 16'h0001);
  assign SubModule_SA_3D__zz_io_MatrixB_0 = SubModule_WeightCache_mData_0;
  assign SubModule_SA_3D__zz_io_B_Valid_0 = SubModule_WeightCache_MatrixCol_Switch[0];
  assign SubModule_Img2Col_start = (toplevel_SubModule_WeightCache_Weight_Cached_delay_3 && Control_Switch_Conv);
  assign Fsm_Picture_Received = SubModule_Img2Col_LayerEnd;
  assign Fsm_Switch_Conv = Control_Switch_Conv;
  assign Fsm_WeightCached = SubModule_WeightCache_Weight_Cached;
  always @(*) begin
    InputSwitch_m_0_axis_mm2s_tready = SubModule_WeightCache_s_axis_s2mm_tready;
    if(SubModule_WeightCache_s_axis_s2mm_tready) begin
      InputSwitch_m_0_axis_mm2s_tready = SubModule_WeightCache_s_axis_s2mm_tready;
    end else begin
      InputSwitch_m_0_axis_mm2s_tready = 1'b0;
    end
  end

  assign Fsm_Matrix_Received = 1'b0;
  assign SubModule_DataArrange_OutChannel = Img2Col_OutFeature_Channel[9:0];
  assign m_axis_mm2s_tdata = SubModule_DataArrange_mData_payload;
  assign m_axis_mm2s_tlast = SubModule_DataArrange_mLast;
  assign m_axis_mm2s_tvalid = SubModule_DataArrange_mData_valid;
  assign m_axis_mm2s_tkeep = 8'hff;
  assign SubModule_DataArrange_sData_0 = SubModule_SA_3D_Matrix_C_payload_0[7:0];
  always @(*) begin
    SubModule_DataArrange_sValid[0] = SubModule_SA_3D_Matrix_C_valid_0;
    SubModule_DataArrange_sValid[1] = SubModule_SA_3D_Matrix_C_valid_1;
    SubModule_DataArrange_sValid[2] = SubModule_SA_3D_Matrix_C_valid_2;
    SubModule_DataArrange_sValid[3] = SubModule_SA_3D_Matrix_C_valid_3;
    SubModule_DataArrange_sValid[4] = SubModule_SA_3D_Matrix_C_valid_4;
    SubModule_DataArrange_sValid[5] = SubModule_SA_3D_Matrix_C_valid_5;
    SubModule_DataArrange_sValid[6] = SubModule_SA_3D_Matrix_C_valid_6;
    SubModule_DataArrange_sValid[7] = SubModule_SA_3D_Matrix_C_valid_7;
  end

  assign SubModule_DataArrange_sData_1 = SubModule_SA_3D_Matrix_C_payload_1[7:0];
  assign SubModule_DataArrange_sData_2 = SubModule_SA_3D_Matrix_C_payload_2[7:0];
  assign SubModule_DataArrange_sData_3 = SubModule_SA_3D_Matrix_C_payload_3[7:0];
  assign SubModule_DataArrange_sData_4 = SubModule_SA_3D_Matrix_C_payload_4[7:0];
  assign SubModule_DataArrange_sData_5 = SubModule_SA_3D_Matrix_C_payload_5[7:0];
  assign SubModule_DataArrange_sData_6 = SubModule_SA_3D_Matrix_C_payload_6[7:0];
  assign SubModule_DataArrange_sData_7 = SubModule_SA_3D_Matrix_C_payload_7[7:0];
  assign LayerEnd = SubModule_DataArrange_LayerEnd;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= TopCtrl_Enum_IDLE;
      InitCnt_count <= 3'b000;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l19) begin
        InitCnt_count <= (InitCnt_count + 3'b001);
        if(InitCnt_valid) begin
          InitCnt_count <= 3'b000;
        end
      end
    end
  end

  always @(posedge clk) begin
    _zz_io_MatrixB_1 <= SubModule_WeightCache_mData_1;
    _zz_io_B_Valid_1 <= SubModule_WeightCache_MatrixCol_Switch[1];
    _zz_io_MatrixB_2 <= SubModule_WeightCache_mData_2;
    _zz_io_MatrixB_2_1 <= _zz_io_MatrixB_2;
    _zz_io_B_Valid_2 <= SubModule_WeightCache_MatrixCol_Switch[2];
    _zz_io_B_Valid_2_1 <= _zz_io_B_Valid_2;
    _zz_io_MatrixB_3 <= SubModule_WeightCache_mData_3;
    _zz_io_MatrixB_3_1 <= _zz_io_MatrixB_3;
    _zz_io_MatrixB_3_2 <= _zz_io_MatrixB_3_1;
    _zz_io_B_Valid_3 <= SubModule_WeightCache_MatrixCol_Switch[3];
    _zz_io_B_Valid_3_1 <= _zz_io_B_Valid_3;
    _zz_io_B_Valid_3_2 <= _zz_io_B_Valid_3_1;
    _zz_io_MatrixB_4 <= SubModule_WeightCache_mData_4;
    _zz_io_MatrixB_4_1 <= _zz_io_MatrixB_4;
    _zz_io_MatrixB_4_2 <= _zz_io_MatrixB_4_1;
    _zz_io_MatrixB_4_3 <= _zz_io_MatrixB_4_2;
    _zz_io_B_Valid_4 <= SubModule_WeightCache_MatrixCol_Switch[4];
    _zz_io_B_Valid_4_1 <= _zz_io_B_Valid_4;
    _zz_io_B_Valid_4_2 <= _zz_io_B_Valid_4_1;
    _zz_io_B_Valid_4_3 <= _zz_io_B_Valid_4_2;
    _zz_io_MatrixB_5 <= SubModule_WeightCache_mData_5;
    _zz_io_MatrixB_5_1 <= _zz_io_MatrixB_5;
    _zz_io_MatrixB_5_2 <= _zz_io_MatrixB_5_1;
    _zz_io_MatrixB_5_3 <= _zz_io_MatrixB_5_2;
    _zz_io_MatrixB_5_4 <= _zz_io_MatrixB_5_3;
    _zz_io_B_Valid_5 <= SubModule_WeightCache_MatrixCol_Switch[5];
    _zz_io_B_Valid_5_1 <= _zz_io_B_Valid_5;
    _zz_io_B_Valid_5_2 <= _zz_io_B_Valid_5_1;
    _zz_io_B_Valid_5_3 <= _zz_io_B_Valid_5_2;
    _zz_io_B_Valid_5_4 <= _zz_io_B_Valid_5_3;
    _zz_io_MatrixB_6 <= SubModule_WeightCache_mData_6;
    _zz_io_MatrixB_6_1 <= _zz_io_MatrixB_6;
    _zz_io_MatrixB_6_2 <= _zz_io_MatrixB_6_1;
    _zz_io_MatrixB_6_3 <= _zz_io_MatrixB_6_2;
    _zz_io_MatrixB_6_4 <= _zz_io_MatrixB_6_3;
    _zz_io_MatrixB_6_5 <= _zz_io_MatrixB_6_4;
    _zz_io_B_Valid_6 <= SubModule_WeightCache_MatrixCol_Switch[6];
    _zz_io_B_Valid_6_1 <= _zz_io_B_Valid_6;
    _zz_io_B_Valid_6_2 <= _zz_io_B_Valid_6_1;
    _zz_io_B_Valid_6_3 <= _zz_io_B_Valid_6_2;
    _zz_io_B_Valid_6_4 <= _zz_io_B_Valid_6_3;
    _zz_io_B_Valid_6_5 <= _zz_io_B_Valid_6_4;
    _zz_io_MatrixB_7 <= SubModule_WeightCache_mData_7;
    _zz_io_MatrixB_7_1 <= _zz_io_MatrixB_7;
    _zz_io_MatrixB_7_2 <= _zz_io_MatrixB_7_1;
    _zz_io_MatrixB_7_3 <= _zz_io_MatrixB_7_2;
    _zz_io_MatrixB_7_4 <= _zz_io_MatrixB_7_3;
    _zz_io_MatrixB_7_5 <= _zz_io_MatrixB_7_4;
    _zz_io_MatrixB_7_6 <= _zz_io_MatrixB_7_5;
    _zz_io_B_Valid_7 <= SubModule_WeightCache_MatrixCol_Switch[7];
    _zz_io_B_Valid_7_1 <= _zz_io_B_Valid_7;
    _zz_io_B_Valid_7_2 <= _zz_io_B_Valid_7_1;
    _zz_io_B_Valid_7_3 <= _zz_io_B_Valid_7_2;
    _zz_io_B_Valid_7_4 <= _zz_io_B_Valid_7_3;
    _zz_io_B_Valid_7_5 <= _zz_io_B_Valid_7_4;
    _zz_io_B_Valid_7_6 <= _zz_io_B_Valid_7_5;
    _zz_io_MatrixB_8 <= SubModule_WeightCache_mData_8;
    _zz_io_MatrixB_8_1 <= _zz_io_MatrixB_8;
    _zz_io_MatrixB_8_2 <= _zz_io_MatrixB_8_1;
    _zz_io_MatrixB_8_3 <= _zz_io_MatrixB_8_2;
    _zz_io_MatrixB_8_4 <= _zz_io_MatrixB_8_3;
    _zz_io_MatrixB_8_5 <= _zz_io_MatrixB_8_4;
    _zz_io_MatrixB_8_6 <= _zz_io_MatrixB_8_5;
    _zz_io_MatrixB_8_7 <= _zz_io_MatrixB_8_6;
    _zz_io_B_Valid_8 <= SubModule_WeightCache_MatrixCol_Switch[8];
    _zz_io_B_Valid_8_1 <= _zz_io_B_Valid_8;
    _zz_io_B_Valid_8_2 <= _zz_io_B_Valid_8_1;
    _zz_io_B_Valid_8_3 <= _zz_io_B_Valid_8_2;
    _zz_io_B_Valid_8_4 <= _zz_io_B_Valid_8_3;
    _zz_io_B_Valid_8_5 <= _zz_io_B_Valid_8_4;
    _zz_io_B_Valid_8_6 <= _zz_io_B_Valid_8_5;
    _zz_io_B_Valid_8_7 <= _zz_io_B_Valid_8_6;
    _zz_io_MatrixB_9 <= SubModule_WeightCache_mData_9;
    _zz_io_MatrixB_9_1 <= _zz_io_MatrixB_9;
    _zz_io_MatrixB_9_2 <= _zz_io_MatrixB_9_1;
    _zz_io_MatrixB_9_3 <= _zz_io_MatrixB_9_2;
    _zz_io_MatrixB_9_4 <= _zz_io_MatrixB_9_3;
    _zz_io_MatrixB_9_5 <= _zz_io_MatrixB_9_4;
    _zz_io_MatrixB_9_6 <= _zz_io_MatrixB_9_5;
    _zz_io_MatrixB_9_7 <= _zz_io_MatrixB_9_6;
    _zz_io_MatrixB_9_8 <= _zz_io_MatrixB_9_7;
    _zz_io_B_Valid_9 <= SubModule_WeightCache_MatrixCol_Switch[9];
    _zz_io_B_Valid_9_1 <= _zz_io_B_Valid_9;
    _zz_io_B_Valid_9_2 <= _zz_io_B_Valid_9_1;
    _zz_io_B_Valid_9_3 <= _zz_io_B_Valid_9_2;
    _zz_io_B_Valid_9_4 <= _zz_io_B_Valid_9_3;
    _zz_io_B_Valid_9_5 <= _zz_io_B_Valid_9_4;
    _zz_io_B_Valid_9_6 <= _zz_io_B_Valid_9_5;
    _zz_io_B_Valid_9_7 <= _zz_io_B_Valid_9_6;
    _zz_io_B_Valid_9_8 <= _zz_io_B_Valid_9_7;
    _zz_io_MatrixB_10 <= SubModule_WeightCache_mData_10;
    _zz_io_MatrixB_10_1 <= _zz_io_MatrixB_10;
    _zz_io_MatrixB_10_2 <= _zz_io_MatrixB_10_1;
    _zz_io_MatrixB_10_3 <= _zz_io_MatrixB_10_2;
    _zz_io_MatrixB_10_4 <= _zz_io_MatrixB_10_3;
    _zz_io_MatrixB_10_5 <= _zz_io_MatrixB_10_4;
    _zz_io_MatrixB_10_6 <= _zz_io_MatrixB_10_5;
    _zz_io_MatrixB_10_7 <= _zz_io_MatrixB_10_6;
    _zz_io_MatrixB_10_8 <= _zz_io_MatrixB_10_7;
    _zz_io_MatrixB_10_9 <= _zz_io_MatrixB_10_8;
    _zz_io_B_Valid_10 <= SubModule_WeightCache_MatrixCol_Switch[10];
    _zz_io_B_Valid_10_1 <= _zz_io_B_Valid_10;
    _zz_io_B_Valid_10_2 <= _zz_io_B_Valid_10_1;
    _zz_io_B_Valid_10_3 <= _zz_io_B_Valid_10_2;
    _zz_io_B_Valid_10_4 <= _zz_io_B_Valid_10_3;
    _zz_io_B_Valid_10_5 <= _zz_io_B_Valid_10_4;
    _zz_io_B_Valid_10_6 <= _zz_io_B_Valid_10_5;
    _zz_io_B_Valid_10_7 <= _zz_io_B_Valid_10_6;
    _zz_io_B_Valid_10_8 <= _zz_io_B_Valid_10_7;
    _zz_io_B_Valid_10_9 <= _zz_io_B_Valid_10_8;
    _zz_io_MatrixB_11 <= SubModule_WeightCache_mData_11;
    _zz_io_MatrixB_11_1 <= _zz_io_MatrixB_11;
    _zz_io_MatrixB_11_2 <= _zz_io_MatrixB_11_1;
    _zz_io_MatrixB_11_3 <= _zz_io_MatrixB_11_2;
    _zz_io_MatrixB_11_4 <= _zz_io_MatrixB_11_3;
    _zz_io_MatrixB_11_5 <= _zz_io_MatrixB_11_4;
    _zz_io_MatrixB_11_6 <= _zz_io_MatrixB_11_5;
    _zz_io_MatrixB_11_7 <= _zz_io_MatrixB_11_6;
    _zz_io_MatrixB_11_8 <= _zz_io_MatrixB_11_7;
    _zz_io_MatrixB_11_9 <= _zz_io_MatrixB_11_8;
    _zz_io_MatrixB_11_10 <= _zz_io_MatrixB_11_9;
    _zz_io_B_Valid_11 <= SubModule_WeightCache_MatrixCol_Switch[11];
    _zz_io_B_Valid_11_1 <= _zz_io_B_Valid_11;
    _zz_io_B_Valid_11_2 <= _zz_io_B_Valid_11_1;
    _zz_io_B_Valid_11_3 <= _zz_io_B_Valid_11_2;
    _zz_io_B_Valid_11_4 <= _zz_io_B_Valid_11_3;
    _zz_io_B_Valid_11_5 <= _zz_io_B_Valid_11_4;
    _zz_io_B_Valid_11_6 <= _zz_io_B_Valid_11_5;
    _zz_io_B_Valid_11_7 <= _zz_io_B_Valid_11_6;
    _zz_io_B_Valid_11_8 <= _zz_io_B_Valid_11_7;
    _zz_io_B_Valid_11_9 <= _zz_io_B_Valid_11_8;
    _zz_io_B_Valid_11_10 <= _zz_io_B_Valid_11_9;
    _zz_io_MatrixB_12 <= SubModule_WeightCache_mData_12;
    _zz_io_MatrixB_12_1 <= _zz_io_MatrixB_12;
    _zz_io_MatrixB_12_2 <= _zz_io_MatrixB_12_1;
    _zz_io_MatrixB_12_3 <= _zz_io_MatrixB_12_2;
    _zz_io_MatrixB_12_4 <= _zz_io_MatrixB_12_3;
    _zz_io_MatrixB_12_5 <= _zz_io_MatrixB_12_4;
    _zz_io_MatrixB_12_6 <= _zz_io_MatrixB_12_5;
    _zz_io_MatrixB_12_7 <= _zz_io_MatrixB_12_6;
    _zz_io_MatrixB_12_8 <= _zz_io_MatrixB_12_7;
    _zz_io_MatrixB_12_9 <= _zz_io_MatrixB_12_8;
    _zz_io_MatrixB_12_10 <= _zz_io_MatrixB_12_9;
    _zz_io_MatrixB_12_11 <= _zz_io_MatrixB_12_10;
    _zz_io_B_Valid_12 <= SubModule_WeightCache_MatrixCol_Switch[12];
    _zz_io_B_Valid_12_1 <= _zz_io_B_Valid_12;
    _zz_io_B_Valid_12_2 <= _zz_io_B_Valid_12_1;
    _zz_io_B_Valid_12_3 <= _zz_io_B_Valid_12_2;
    _zz_io_B_Valid_12_4 <= _zz_io_B_Valid_12_3;
    _zz_io_B_Valid_12_5 <= _zz_io_B_Valid_12_4;
    _zz_io_B_Valid_12_6 <= _zz_io_B_Valid_12_5;
    _zz_io_B_Valid_12_7 <= _zz_io_B_Valid_12_6;
    _zz_io_B_Valid_12_8 <= _zz_io_B_Valid_12_7;
    _zz_io_B_Valid_12_9 <= _zz_io_B_Valid_12_8;
    _zz_io_B_Valid_12_10 <= _zz_io_B_Valid_12_9;
    _zz_io_B_Valid_12_11 <= _zz_io_B_Valid_12_10;
    _zz_io_MatrixB_13 <= SubModule_WeightCache_mData_13;
    _zz_io_MatrixB_13_1 <= _zz_io_MatrixB_13;
    _zz_io_MatrixB_13_2 <= _zz_io_MatrixB_13_1;
    _zz_io_MatrixB_13_3 <= _zz_io_MatrixB_13_2;
    _zz_io_MatrixB_13_4 <= _zz_io_MatrixB_13_3;
    _zz_io_MatrixB_13_5 <= _zz_io_MatrixB_13_4;
    _zz_io_MatrixB_13_6 <= _zz_io_MatrixB_13_5;
    _zz_io_MatrixB_13_7 <= _zz_io_MatrixB_13_6;
    _zz_io_MatrixB_13_8 <= _zz_io_MatrixB_13_7;
    _zz_io_MatrixB_13_9 <= _zz_io_MatrixB_13_8;
    _zz_io_MatrixB_13_10 <= _zz_io_MatrixB_13_9;
    _zz_io_MatrixB_13_11 <= _zz_io_MatrixB_13_10;
    _zz_io_MatrixB_13_12 <= _zz_io_MatrixB_13_11;
    _zz_io_B_Valid_13 <= SubModule_WeightCache_MatrixCol_Switch[13];
    _zz_io_B_Valid_13_1 <= _zz_io_B_Valid_13;
    _zz_io_B_Valid_13_2 <= _zz_io_B_Valid_13_1;
    _zz_io_B_Valid_13_3 <= _zz_io_B_Valid_13_2;
    _zz_io_B_Valid_13_4 <= _zz_io_B_Valid_13_3;
    _zz_io_B_Valid_13_5 <= _zz_io_B_Valid_13_4;
    _zz_io_B_Valid_13_6 <= _zz_io_B_Valid_13_5;
    _zz_io_B_Valid_13_7 <= _zz_io_B_Valid_13_6;
    _zz_io_B_Valid_13_8 <= _zz_io_B_Valid_13_7;
    _zz_io_B_Valid_13_9 <= _zz_io_B_Valid_13_8;
    _zz_io_B_Valid_13_10 <= _zz_io_B_Valid_13_9;
    _zz_io_B_Valid_13_11 <= _zz_io_B_Valid_13_10;
    _zz_io_B_Valid_13_12 <= _zz_io_B_Valid_13_11;
    _zz_io_MatrixB_14 <= SubModule_WeightCache_mData_14;
    _zz_io_MatrixB_14_1 <= _zz_io_MatrixB_14;
    _zz_io_MatrixB_14_2 <= _zz_io_MatrixB_14_1;
    _zz_io_MatrixB_14_3 <= _zz_io_MatrixB_14_2;
    _zz_io_MatrixB_14_4 <= _zz_io_MatrixB_14_3;
    _zz_io_MatrixB_14_5 <= _zz_io_MatrixB_14_4;
    _zz_io_MatrixB_14_6 <= _zz_io_MatrixB_14_5;
    _zz_io_MatrixB_14_7 <= _zz_io_MatrixB_14_6;
    _zz_io_MatrixB_14_8 <= _zz_io_MatrixB_14_7;
    _zz_io_MatrixB_14_9 <= _zz_io_MatrixB_14_8;
    _zz_io_MatrixB_14_10 <= _zz_io_MatrixB_14_9;
    _zz_io_MatrixB_14_11 <= _zz_io_MatrixB_14_10;
    _zz_io_MatrixB_14_12 <= _zz_io_MatrixB_14_11;
    _zz_io_MatrixB_14_13 <= _zz_io_MatrixB_14_12;
    _zz_io_B_Valid_14 <= SubModule_WeightCache_MatrixCol_Switch[14];
    _zz_io_B_Valid_14_1 <= _zz_io_B_Valid_14;
    _zz_io_B_Valid_14_2 <= _zz_io_B_Valid_14_1;
    _zz_io_B_Valid_14_3 <= _zz_io_B_Valid_14_2;
    _zz_io_B_Valid_14_4 <= _zz_io_B_Valid_14_3;
    _zz_io_B_Valid_14_5 <= _zz_io_B_Valid_14_4;
    _zz_io_B_Valid_14_6 <= _zz_io_B_Valid_14_5;
    _zz_io_B_Valid_14_7 <= _zz_io_B_Valid_14_6;
    _zz_io_B_Valid_14_8 <= _zz_io_B_Valid_14_7;
    _zz_io_B_Valid_14_9 <= _zz_io_B_Valid_14_8;
    _zz_io_B_Valid_14_10 <= _zz_io_B_Valid_14_9;
    _zz_io_B_Valid_14_11 <= _zz_io_B_Valid_14_10;
    _zz_io_B_Valid_14_12 <= _zz_io_B_Valid_14_11;
    _zz_io_B_Valid_14_13 <= _zz_io_B_Valid_14_12;
    _zz_io_MatrixB_15 <= SubModule_WeightCache_mData_15;
    _zz_io_MatrixB_15_1 <= _zz_io_MatrixB_15;
    _zz_io_MatrixB_15_2 <= _zz_io_MatrixB_15_1;
    _zz_io_MatrixB_15_3 <= _zz_io_MatrixB_15_2;
    _zz_io_MatrixB_15_4 <= _zz_io_MatrixB_15_3;
    _zz_io_MatrixB_15_5 <= _zz_io_MatrixB_15_4;
    _zz_io_MatrixB_15_6 <= _zz_io_MatrixB_15_5;
    _zz_io_MatrixB_15_7 <= _zz_io_MatrixB_15_6;
    _zz_io_MatrixB_15_8 <= _zz_io_MatrixB_15_7;
    _zz_io_MatrixB_15_9 <= _zz_io_MatrixB_15_8;
    _zz_io_MatrixB_15_10 <= _zz_io_MatrixB_15_9;
    _zz_io_MatrixB_15_11 <= _zz_io_MatrixB_15_10;
    _zz_io_MatrixB_15_12 <= _zz_io_MatrixB_15_11;
    _zz_io_MatrixB_15_13 <= _zz_io_MatrixB_15_12;
    _zz_io_MatrixB_15_14 <= _zz_io_MatrixB_15_13;
    _zz_io_B_Valid_15 <= SubModule_WeightCache_MatrixCol_Switch[15];
    _zz_io_B_Valid_15_1 <= _zz_io_B_Valid_15;
    _zz_io_B_Valid_15_2 <= _zz_io_B_Valid_15_1;
    _zz_io_B_Valid_15_3 <= _zz_io_B_Valid_15_2;
    _zz_io_B_Valid_15_4 <= _zz_io_B_Valid_15_3;
    _zz_io_B_Valid_15_5 <= _zz_io_B_Valid_15_4;
    _zz_io_B_Valid_15_6 <= _zz_io_B_Valid_15_5;
    _zz_io_B_Valid_15_7 <= _zz_io_B_Valid_15_6;
    _zz_io_B_Valid_15_8 <= _zz_io_B_Valid_15_7;
    _zz_io_B_Valid_15_9 <= _zz_io_B_Valid_15_8;
    _zz_io_B_Valid_15_10 <= _zz_io_B_Valid_15_9;
    _zz_io_B_Valid_15_11 <= _zz_io_B_Valid_15_10;
    _zz_io_B_Valid_15_12 <= _zz_io_B_Valid_15_11;
    _zz_io_B_Valid_15_13 <= _zz_io_B_Valid_15_12;
    _zz_io_B_Valid_15_14 <= _zz_io_B_Valid_15_13;
    _zz_io_MatrixB_16 <= SubModule_WeightCache_mData_16;
    _zz_io_MatrixB_16_1 <= _zz_io_MatrixB_16;
    _zz_io_MatrixB_16_2 <= _zz_io_MatrixB_16_1;
    _zz_io_MatrixB_16_3 <= _zz_io_MatrixB_16_2;
    _zz_io_MatrixB_16_4 <= _zz_io_MatrixB_16_3;
    _zz_io_MatrixB_16_5 <= _zz_io_MatrixB_16_4;
    _zz_io_MatrixB_16_6 <= _zz_io_MatrixB_16_5;
    _zz_io_MatrixB_16_7 <= _zz_io_MatrixB_16_6;
    _zz_io_MatrixB_16_8 <= _zz_io_MatrixB_16_7;
    _zz_io_MatrixB_16_9 <= _zz_io_MatrixB_16_8;
    _zz_io_MatrixB_16_10 <= _zz_io_MatrixB_16_9;
    _zz_io_MatrixB_16_11 <= _zz_io_MatrixB_16_10;
    _zz_io_MatrixB_16_12 <= _zz_io_MatrixB_16_11;
    _zz_io_MatrixB_16_13 <= _zz_io_MatrixB_16_12;
    _zz_io_MatrixB_16_14 <= _zz_io_MatrixB_16_13;
    _zz_io_MatrixB_16_15 <= _zz_io_MatrixB_16_14;
    _zz_io_B_Valid_16 <= SubModule_WeightCache_MatrixCol_Switch[16];
    _zz_io_B_Valid_16_1 <= _zz_io_B_Valid_16;
    _zz_io_B_Valid_16_2 <= _zz_io_B_Valid_16_1;
    _zz_io_B_Valid_16_3 <= _zz_io_B_Valid_16_2;
    _zz_io_B_Valid_16_4 <= _zz_io_B_Valid_16_3;
    _zz_io_B_Valid_16_5 <= _zz_io_B_Valid_16_4;
    _zz_io_B_Valid_16_6 <= _zz_io_B_Valid_16_5;
    _zz_io_B_Valid_16_7 <= _zz_io_B_Valid_16_6;
    _zz_io_B_Valid_16_8 <= _zz_io_B_Valid_16_7;
    _zz_io_B_Valid_16_9 <= _zz_io_B_Valid_16_8;
    _zz_io_B_Valid_16_10 <= _zz_io_B_Valid_16_9;
    _zz_io_B_Valid_16_11 <= _zz_io_B_Valid_16_10;
    _zz_io_B_Valid_16_12 <= _zz_io_B_Valid_16_11;
    _zz_io_B_Valid_16_13 <= _zz_io_B_Valid_16_12;
    _zz_io_B_Valid_16_14 <= _zz_io_B_Valid_16_13;
    _zz_io_B_Valid_16_15 <= _zz_io_B_Valid_16_14;
    _zz_io_MatrixB_17 <= SubModule_WeightCache_mData_17;
    _zz_io_MatrixB_17_1 <= _zz_io_MatrixB_17;
    _zz_io_MatrixB_17_2 <= _zz_io_MatrixB_17_1;
    _zz_io_MatrixB_17_3 <= _zz_io_MatrixB_17_2;
    _zz_io_MatrixB_17_4 <= _zz_io_MatrixB_17_3;
    _zz_io_MatrixB_17_5 <= _zz_io_MatrixB_17_4;
    _zz_io_MatrixB_17_6 <= _zz_io_MatrixB_17_5;
    _zz_io_MatrixB_17_7 <= _zz_io_MatrixB_17_6;
    _zz_io_MatrixB_17_8 <= _zz_io_MatrixB_17_7;
    _zz_io_MatrixB_17_9 <= _zz_io_MatrixB_17_8;
    _zz_io_MatrixB_17_10 <= _zz_io_MatrixB_17_9;
    _zz_io_MatrixB_17_11 <= _zz_io_MatrixB_17_10;
    _zz_io_MatrixB_17_12 <= _zz_io_MatrixB_17_11;
    _zz_io_MatrixB_17_13 <= _zz_io_MatrixB_17_12;
    _zz_io_MatrixB_17_14 <= _zz_io_MatrixB_17_13;
    _zz_io_MatrixB_17_15 <= _zz_io_MatrixB_17_14;
    _zz_io_MatrixB_17_16 <= _zz_io_MatrixB_17_15;
    _zz_io_B_Valid_17 <= SubModule_WeightCache_MatrixCol_Switch[17];
    _zz_io_B_Valid_17_1 <= _zz_io_B_Valid_17;
    _zz_io_B_Valid_17_2 <= _zz_io_B_Valid_17_1;
    _zz_io_B_Valid_17_3 <= _zz_io_B_Valid_17_2;
    _zz_io_B_Valid_17_4 <= _zz_io_B_Valid_17_3;
    _zz_io_B_Valid_17_5 <= _zz_io_B_Valid_17_4;
    _zz_io_B_Valid_17_6 <= _zz_io_B_Valid_17_5;
    _zz_io_B_Valid_17_7 <= _zz_io_B_Valid_17_6;
    _zz_io_B_Valid_17_8 <= _zz_io_B_Valid_17_7;
    _zz_io_B_Valid_17_9 <= _zz_io_B_Valid_17_8;
    _zz_io_B_Valid_17_10 <= _zz_io_B_Valid_17_9;
    _zz_io_B_Valid_17_11 <= _zz_io_B_Valid_17_10;
    _zz_io_B_Valid_17_12 <= _zz_io_B_Valid_17_11;
    _zz_io_B_Valid_17_13 <= _zz_io_B_Valid_17_12;
    _zz_io_B_Valid_17_14 <= _zz_io_B_Valid_17_13;
    _zz_io_B_Valid_17_15 <= _zz_io_B_Valid_17_14;
    _zz_io_B_Valid_17_16 <= _zz_io_B_Valid_17_15;
    _zz_io_MatrixB_18 <= SubModule_WeightCache_mData_18;
    _zz_io_MatrixB_18_1 <= _zz_io_MatrixB_18;
    _zz_io_MatrixB_18_2 <= _zz_io_MatrixB_18_1;
    _zz_io_MatrixB_18_3 <= _zz_io_MatrixB_18_2;
    _zz_io_MatrixB_18_4 <= _zz_io_MatrixB_18_3;
    _zz_io_MatrixB_18_5 <= _zz_io_MatrixB_18_4;
    _zz_io_MatrixB_18_6 <= _zz_io_MatrixB_18_5;
    _zz_io_MatrixB_18_7 <= _zz_io_MatrixB_18_6;
    _zz_io_MatrixB_18_8 <= _zz_io_MatrixB_18_7;
    _zz_io_MatrixB_18_9 <= _zz_io_MatrixB_18_8;
    _zz_io_MatrixB_18_10 <= _zz_io_MatrixB_18_9;
    _zz_io_MatrixB_18_11 <= _zz_io_MatrixB_18_10;
    _zz_io_MatrixB_18_12 <= _zz_io_MatrixB_18_11;
    _zz_io_MatrixB_18_13 <= _zz_io_MatrixB_18_12;
    _zz_io_MatrixB_18_14 <= _zz_io_MatrixB_18_13;
    _zz_io_MatrixB_18_15 <= _zz_io_MatrixB_18_14;
    _zz_io_MatrixB_18_16 <= _zz_io_MatrixB_18_15;
    _zz_io_MatrixB_18_17 <= _zz_io_MatrixB_18_16;
    _zz_io_B_Valid_18 <= SubModule_WeightCache_MatrixCol_Switch[18];
    _zz_io_B_Valid_18_1 <= _zz_io_B_Valid_18;
    _zz_io_B_Valid_18_2 <= _zz_io_B_Valid_18_1;
    _zz_io_B_Valid_18_3 <= _zz_io_B_Valid_18_2;
    _zz_io_B_Valid_18_4 <= _zz_io_B_Valid_18_3;
    _zz_io_B_Valid_18_5 <= _zz_io_B_Valid_18_4;
    _zz_io_B_Valid_18_6 <= _zz_io_B_Valid_18_5;
    _zz_io_B_Valid_18_7 <= _zz_io_B_Valid_18_6;
    _zz_io_B_Valid_18_8 <= _zz_io_B_Valid_18_7;
    _zz_io_B_Valid_18_9 <= _zz_io_B_Valid_18_8;
    _zz_io_B_Valid_18_10 <= _zz_io_B_Valid_18_9;
    _zz_io_B_Valid_18_11 <= _zz_io_B_Valid_18_10;
    _zz_io_B_Valid_18_12 <= _zz_io_B_Valid_18_11;
    _zz_io_B_Valid_18_13 <= _zz_io_B_Valid_18_12;
    _zz_io_B_Valid_18_14 <= _zz_io_B_Valid_18_13;
    _zz_io_B_Valid_18_15 <= _zz_io_B_Valid_18_14;
    _zz_io_B_Valid_18_16 <= _zz_io_B_Valid_18_15;
    _zz_io_B_Valid_18_17 <= _zz_io_B_Valid_18_16;
    _zz_io_MatrixB_19 <= SubModule_WeightCache_mData_19;
    _zz_io_MatrixB_19_1 <= _zz_io_MatrixB_19;
    _zz_io_MatrixB_19_2 <= _zz_io_MatrixB_19_1;
    _zz_io_MatrixB_19_3 <= _zz_io_MatrixB_19_2;
    _zz_io_MatrixB_19_4 <= _zz_io_MatrixB_19_3;
    _zz_io_MatrixB_19_5 <= _zz_io_MatrixB_19_4;
    _zz_io_MatrixB_19_6 <= _zz_io_MatrixB_19_5;
    _zz_io_MatrixB_19_7 <= _zz_io_MatrixB_19_6;
    _zz_io_MatrixB_19_8 <= _zz_io_MatrixB_19_7;
    _zz_io_MatrixB_19_9 <= _zz_io_MatrixB_19_8;
    _zz_io_MatrixB_19_10 <= _zz_io_MatrixB_19_9;
    _zz_io_MatrixB_19_11 <= _zz_io_MatrixB_19_10;
    _zz_io_MatrixB_19_12 <= _zz_io_MatrixB_19_11;
    _zz_io_MatrixB_19_13 <= _zz_io_MatrixB_19_12;
    _zz_io_MatrixB_19_14 <= _zz_io_MatrixB_19_13;
    _zz_io_MatrixB_19_15 <= _zz_io_MatrixB_19_14;
    _zz_io_MatrixB_19_16 <= _zz_io_MatrixB_19_15;
    _zz_io_MatrixB_19_17 <= _zz_io_MatrixB_19_16;
    _zz_io_MatrixB_19_18 <= _zz_io_MatrixB_19_17;
    _zz_io_B_Valid_19 <= SubModule_WeightCache_MatrixCol_Switch[19];
    _zz_io_B_Valid_19_1 <= _zz_io_B_Valid_19;
    _zz_io_B_Valid_19_2 <= _zz_io_B_Valid_19_1;
    _zz_io_B_Valid_19_3 <= _zz_io_B_Valid_19_2;
    _zz_io_B_Valid_19_4 <= _zz_io_B_Valid_19_3;
    _zz_io_B_Valid_19_5 <= _zz_io_B_Valid_19_4;
    _zz_io_B_Valid_19_6 <= _zz_io_B_Valid_19_5;
    _zz_io_B_Valid_19_7 <= _zz_io_B_Valid_19_6;
    _zz_io_B_Valid_19_8 <= _zz_io_B_Valid_19_7;
    _zz_io_B_Valid_19_9 <= _zz_io_B_Valid_19_8;
    _zz_io_B_Valid_19_10 <= _zz_io_B_Valid_19_9;
    _zz_io_B_Valid_19_11 <= _zz_io_B_Valid_19_10;
    _zz_io_B_Valid_19_12 <= _zz_io_B_Valid_19_11;
    _zz_io_B_Valid_19_13 <= _zz_io_B_Valid_19_12;
    _zz_io_B_Valid_19_14 <= _zz_io_B_Valid_19_13;
    _zz_io_B_Valid_19_15 <= _zz_io_B_Valid_19_14;
    _zz_io_B_Valid_19_16 <= _zz_io_B_Valid_19_15;
    _zz_io_B_Valid_19_17 <= _zz_io_B_Valid_19_16;
    _zz_io_B_Valid_19_18 <= _zz_io_B_Valid_19_17;
    _zz_io_MatrixB_20 <= SubModule_WeightCache_mData_20;
    _zz_io_MatrixB_20_1 <= _zz_io_MatrixB_20;
    _zz_io_MatrixB_20_2 <= _zz_io_MatrixB_20_1;
    _zz_io_MatrixB_20_3 <= _zz_io_MatrixB_20_2;
    _zz_io_MatrixB_20_4 <= _zz_io_MatrixB_20_3;
    _zz_io_MatrixB_20_5 <= _zz_io_MatrixB_20_4;
    _zz_io_MatrixB_20_6 <= _zz_io_MatrixB_20_5;
    _zz_io_MatrixB_20_7 <= _zz_io_MatrixB_20_6;
    _zz_io_MatrixB_20_8 <= _zz_io_MatrixB_20_7;
    _zz_io_MatrixB_20_9 <= _zz_io_MatrixB_20_8;
    _zz_io_MatrixB_20_10 <= _zz_io_MatrixB_20_9;
    _zz_io_MatrixB_20_11 <= _zz_io_MatrixB_20_10;
    _zz_io_MatrixB_20_12 <= _zz_io_MatrixB_20_11;
    _zz_io_MatrixB_20_13 <= _zz_io_MatrixB_20_12;
    _zz_io_MatrixB_20_14 <= _zz_io_MatrixB_20_13;
    _zz_io_MatrixB_20_15 <= _zz_io_MatrixB_20_14;
    _zz_io_MatrixB_20_16 <= _zz_io_MatrixB_20_15;
    _zz_io_MatrixB_20_17 <= _zz_io_MatrixB_20_16;
    _zz_io_MatrixB_20_18 <= _zz_io_MatrixB_20_17;
    _zz_io_MatrixB_20_19 <= _zz_io_MatrixB_20_18;
    _zz_io_B_Valid_20 <= SubModule_WeightCache_MatrixCol_Switch[20];
    _zz_io_B_Valid_20_1 <= _zz_io_B_Valid_20;
    _zz_io_B_Valid_20_2 <= _zz_io_B_Valid_20_1;
    _zz_io_B_Valid_20_3 <= _zz_io_B_Valid_20_2;
    _zz_io_B_Valid_20_4 <= _zz_io_B_Valid_20_3;
    _zz_io_B_Valid_20_5 <= _zz_io_B_Valid_20_4;
    _zz_io_B_Valid_20_6 <= _zz_io_B_Valid_20_5;
    _zz_io_B_Valid_20_7 <= _zz_io_B_Valid_20_6;
    _zz_io_B_Valid_20_8 <= _zz_io_B_Valid_20_7;
    _zz_io_B_Valid_20_9 <= _zz_io_B_Valid_20_8;
    _zz_io_B_Valid_20_10 <= _zz_io_B_Valid_20_9;
    _zz_io_B_Valid_20_11 <= _zz_io_B_Valid_20_10;
    _zz_io_B_Valid_20_12 <= _zz_io_B_Valid_20_11;
    _zz_io_B_Valid_20_13 <= _zz_io_B_Valid_20_12;
    _zz_io_B_Valid_20_14 <= _zz_io_B_Valid_20_13;
    _zz_io_B_Valid_20_15 <= _zz_io_B_Valid_20_14;
    _zz_io_B_Valid_20_16 <= _zz_io_B_Valid_20_15;
    _zz_io_B_Valid_20_17 <= _zz_io_B_Valid_20_16;
    _zz_io_B_Valid_20_18 <= _zz_io_B_Valid_20_17;
    _zz_io_B_Valid_20_19 <= _zz_io_B_Valid_20_18;
    _zz_io_MatrixB_21 <= SubModule_WeightCache_mData_21;
    _zz_io_MatrixB_21_1 <= _zz_io_MatrixB_21;
    _zz_io_MatrixB_21_2 <= _zz_io_MatrixB_21_1;
    _zz_io_MatrixB_21_3 <= _zz_io_MatrixB_21_2;
    _zz_io_MatrixB_21_4 <= _zz_io_MatrixB_21_3;
    _zz_io_MatrixB_21_5 <= _zz_io_MatrixB_21_4;
    _zz_io_MatrixB_21_6 <= _zz_io_MatrixB_21_5;
    _zz_io_MatrixB_21_7 <= _zz_io_MatrixB_21_6;
    _zz_io_MatrixB_21_8 <= _zz_io_MatrixB_21_7;
    _zz_io_MatrixB_21_9 <= _zz_io_MatrixB_21_8;
    _zz_io_MatrixB_21_10 <= _zz_io_MatrixB_21_9;
    _zz_io_MatrixB_21_11 <= _zz_io_MatrixB_21_10;
    _zz_io_MatrixB_21_12 <= _zz_io_MatrixB_21_11;
    _zz_io_MatrixB_21_13 <= _zz_io_MatrixB_21_12;
    _zz_io_MatrixB_21_14 <= _zz_io_MatrixB_21_13;
    _zz_io_MatrixB_21_15 <= _zz_io_MatrixB_21_14;
    _zz_io_MatrixB_21_16 <= _zz_io_MatrixB_21_15;
    _zz_io_MatrixB_21_17 <= _zz_io_MatrixB_21_16;
    _zz_io_MatrixB_21_18 <= _zz_io_MatrixB_21_17;
    _zz_io_MatrixB_21_19 <= _zz_io_MatrixB_21_18;
    _zz_io_MatrixB_21_20 <= _zz_io_MatrixB_21_19;
    _zz_io_B_Valid_21 <= SubModule_WeightCache_MatrixCol_Switch[21];
    _zz_io_B_Valid_21_1 <= _zz_io_B_Valid_21;
    _zz_io_B_Valid_21_2 <= _zz_io_B_Valid_21_1;
    _zz_io_B_Valid_21_3 <= _zz_io_B_Valid_21_2;
    _zz_io_B_Valid_21_4 <= _zz_io_B_Valid_21_3;
    _zz_io_B_Valid_21_5 <= _zz_io_B_Valid_21_4;
    _zz_io_B_Valid_21_6 <= _zz_io_B_Valid_21_5;
    _zz_io_B_Valid_21_7 <= _zz_io_B_Valid_21_6;
    _zz_io_B_Valid_21_8 <= _zz_io_B_Valid_21_7;
    _zz_io_B_Valid_21_9 <= _zz_io_B_Valid_21_8;
    _zz_io_B_Valid_21_10 <= _zz_io_B_Valid_21_9;
    _zz_io_B_Valid_21_11 <= _zz_io_B_Valid_21_10;
    _zz_io_B_Valid_21_12 <= _zz_io_B_Valid_21_11;
    _zz_io_B_Valid_21_13 <= _zz_io_B_Valid_21_12;
    _zz_io_B_Valid_21_14 <= _zz_io_B_Valid_21_13;
    _zz_io_B_Valid_21_15 <= _zz_io_B_Valid_21_14;
    _zz_io_B_Valid_21_16 <= _zz_io_B_Valid_21_15;
    _zz_io_B_Valid_21_17 <= _zz_io_B_Valid_21_16;
    _zz_io_B_Valid_21_18 <= _zz_io_B_Valid_21_17;
    _zz_io_B_Valid_21_19 <= _zz_io_B_Valid_21_18;
    _zz_io_B_Valid_21_20 <= _zz_io_B_Valid_21_19;
    _zz_io_MatrixB_22 <= SubModule_WeightCache_mData_22;
    _zz_io_MatrixB_22_1 <= _zz_io_MatrixB_22;
    _zz_io_MatrixB_22_2 <= _zz_io_MatrixB_22_1;
    _zz_io_MatrixB_22_3 <= _zz_io_MatrixB_22_2;
    _zz_io_MatrixB_22_4 <= _zz_io_MatrixB_22_3;
    _zz_io_MatrixB_22_5 <= _zz_io_MatrixB_22_4;
    _zz_io_MatrixB_22_6 <= _zz_io_MatrixB_22_5;
    _zz_io_MatrixB_22_7 <= _zz_io_MatrixB_22_6;
    _zz_io_MatrixB_22_8 <= _zz_io_MatrixB_22_7;
    _zz_io_MatrixB_22_9 <= _zz_io_MatrixB_22_8;
    _zz_io_MatrixB_22_10 <= _zz_io_MatrixB_22_9;
    _zz_io_MatrixB_22_11 <= _zz_io_MatrixB_22_10;
    _zz_io_MatrixB_22_12 <= _zz_io_MatrixB_22_11;
    _zz_io_MatrixB_22_13 <= _zz_io_MatrixB_22_12;
    _zz_io_MatrixB_22_14 <= _zz_io_MatrixB_22_13;
    _zz_io_MatrixB_22_15 <= _zz_io_MatrixB_22_14;
    _zz_io_MatrixB_22_16 <= _zz_io_MatrixB_22_15;
    _zz_io_MatrixB_22_17 <= _zz_io_MatrixB_22_16;
    _zz_io_MatrixB_22_18 <= _zz_io_MatrixB_22_17;
    _zz_io_MatrixB_22_19 <= _zz_io_MatrixB_22_18;
    _zz_io_MatrixB_22_20 <= _zz_io_MatrixB_22_19;
    _zz_io_MatrixB_22_21 <= _zz_io_MatrixB_22_20;
    _zz_io_B_Valid_22 <= SubModule_WeightCache_MatrixCol_Switch[22];
    _zz_io_B_Valid_22_1 <= _zz_io_B_Valid_22;
    _zz_io_B_Valid_22_2 <= _zz_io_B_Valid_22_1;
    _zz_io_B_Valid_22_3 <= _zz_io_B_Valid_22_2;
    _zz_io_B_Valid_22_4 <= _zz_io_B_Valid_22_3;
    _zz_io_B_Valid_22_5 <= _zz_io_B_Valid_22_4;
    _zz_io_B_Valid_22_6 <= _zz_io_B_Valid_22_5;
    _zz_io_B_Valid_22_7 <= _zz_io_B_Valid_22_6;
    _zz_io_B_Valid_22_8 <= _zz_io_B_Valid_22_7;
    _zz_io_B_Valid_22_9 <= _zz_io_B_Valid_22_8;
    _zz_io_B_Valid_22_10 <= _zz_io_B_Valid_22_9;
    _zz_io_B_Valid_22_11 <= _zz_io_B_Valid_22_10;
    _zz_io_B_Valid_22_12 <= _zz_io_B_Valid_22_11;
    _zz_io_B_Valid_22_13 <= _zz_io_B_Valid_22_12;
    _zz_io_B_Valid_22_14 <= _zz_io_B_Valid_22_13;
    _zz_io_B_Valid_22_15 <= _zz_io_B_Valid_22_14;
    _zz_io_B_Valid_22_16 <= _zz_io_B_Valid_22_15;
    _zz_io_B_Valid_22_17 <= _zz_io_B_Valid_22_16;
    _zz_io_B_Valid_22_18 <= _zz_io_B_Valid_22_17;
    _zz_io_B_Valid_22_19 <= _zz_io_B_Valid_22_18;
    _zz_io_B_Valid_22_20 <= _zz_io_B_Valid_22_19;
    _zz_io_B_Valid_22_21 <= _zz_io_B_Valid_22_20;
    _zz_io_MatrixB_23 <= SubModule_WeightCache_mData_23;
    _zz_io_MatrixB_23_1 <= _zz_io_MatrixB_23;
    _zz_io_MatrixB_23_2 <= _zz_io_MatrixB_23_1;
    _zz_io_MatrixB_23_3 <= _zz_io_MatrixB_23_2;
    _zz_io_MatrixB_23_4 <= _zz_io_MatrixB_23_3;
    _zz_io_MatrixB_23_5 <= _zz_io_MatrixB_23_4;
    _zz_io_MatrixB_23_6 <= _zz_io_MatrixB_23_5;
    _zz_io_MatrixB_23_7 <= _zz_io_MatrixB_23_6;
    _zz_io_MatrixB_23_8 <= _zz_io_MatrixB_23_7;
    _zz_io_MatrixB_23_9 <= _zz_io_MatrixB_23_8;
    _zz_io_MatrixB_23_10 <= _zz_io_MatrixB_23_9;
    _zz_io_MatrixB_23_11 <= _zz_io_MatrixB_23_10;
    _zz_io_MatrixB_23_12 <= _zz_io_MatrixB_23_11;
    _zz_io_MatrixB_23_13 <= _zz_io_MatrixB_23_12;
    _zz_io_MatrixB_23_14 <= _zz_io_MatrixB_23_13;
    _zz_io_MatrixB_23_15 <= _zz_io_MatrixB_23_14;
    _zz_io_MatrixB_23_16 <= _zz_io_MatrixB_23_15;
    _zz_io_MatrixB_23_17 <= _zz_io_MatrixB_23_16;
    _zz_io_MatrixB_23_18 <= _zz_io_MatrixB_23_17;
    _zz_io_MatrixB_23_19 <= _zz_io_MatrixB_23_18;
    _zz_io_MatrixB_23_20 <= _zz_io_MatrixB_23_19;
    _zz_io_MatrixB_23_21 <= _zz_io_MatrixB_23_20;
    _zz_io_MatrixB_23_22 <= _zz_io_MatrixB_23_21;
    _zz_io_B_Valid_23 <= SubModule_WeightCache_MatrixCol_Switch[23];
    _zz_io_B_Valid_23_1 <= _zz_io_B_Valid_23;
    _zz_io_B_Valid_23_2 <= _zz_io_B_Valid_23_1;
    _zz_io_B_Valid_23_3 <= _zz_io_B_Valid_23_2;
    _zz_io_B_Valid_23_4 <= _zz_io_B_Valid_23_3;
    _zz_io_B_Valid_23_5 <= _zz_io_B_Valid_23_4;
    _zz_io_B_Valid_23_6 <= _zz_io_B_Valid_23_5;
    _zz_io_B_Valid_23_7 <= _zz_io_B_Valid_23_6;
    _zz_io_B_Valid_23_8 <= _zz_io_B_Valid_23_7;
    _zz_io_B_Valid_23_9 <= _zz_io_B_Valid_23_8;
    _zz_io_B_Valid_23_10 <= _zz_io_B_Valid_23_9;
    _zz_io_B_Valid_23_11 <= _zz_io_B_Valid_23_10;
    _zz_io_B_Valid_23_12 <= _zz_io_B_Valid_23_11;
    _zz_io_B_Valid_23_13 <= _zz_io_B_Valid_23_12;
    _zz_io_B_Valid_23_14 <= _zz_io_B_Valid_23_13;
    _zz_io_B_Valid_23_15 <= _zz_io_B_Valid_23_14;
    _zz_io_B_Valid_23_16 <= _zz_io_B_Valid_23_15;
    _zz_io_B_Valid_23_17 <= _zz_io_B_Valid_23_16;
    _zz_io_B_Valid_23_18 <= _zz_io_B_Valid_23_17;
    _zz_io_B_Valid_23_19 <= _zz_io_B_Valid_23_18;
    _zz_io_B_Valid_23_20 <= _zz_io_B_Valid_23_19;
    _zz_io_B_Valid_23_21 <= _zz_io_B_Valid_23_20;
    _zz_io_B_Valid_23_22 <= _zz_io_B_Valid_23_21;
    _zz_io_MatrixB_24 <= SubModule_WeightCache_mData_24;
    _zz_io_MatrixB_24_1 <= _zz_io_MatrixB_24;
    _zz_io_MatrixB_24_2 <= _zz_io_MatrixB_24_1;
    _zz_io_MatrixB_24_3 <= _zz_io_MatrixB_24_2;
    _zz_io_MatrixB_24_4 <= _zz_io_MatrixB_24_3;
    _zz_io_MatrixB_24_5 <= _zz_io_MatrixB_24_4;
    _zz_io_MatrixB_24_6 <= _zz_io_MatrixB_24_5;
    _zz_io_MatrixB_24_7 <= _zz_io_MatrixB_24_6;
    _zz_io_MatrixB_24_8 <= _zz_io_MatrixB_24_7;
    _zz_io_MatrixB_24_9 <= _zz_io_MatrixB_24_8;
    _zz_io_MatrixB_24_10 <= _zz_io_MatrixB_24_9;
    _zz_io_MatrixB_24_11 <= _zz_io_MatrixB_24_10;
    _zz_io_MatrixB_24_12 <= _zz_io_MatrixB_24_11;
    _zz_io_MatrixB_24_13 <= _zz_io_MatrixB_24_12;
    _zz_io_MatrixB_24_14 <= _zz_io_MatrixB_24_13;
    _zz_io_MatrixB_24_15 <= _zz_io_MatrixB_24_14;
    _zz_io_MatrixB_24_16 <= _zz_io_MatrixB_24_15;
    _zz_io_MatrixB_24_17 <= _zz_io_MatrixB_24_16;
    _zz_io_MatrixB_24_18 <= _zz_io_MatrixB_24_17;
    _zz_io_MatrixB_24_19 <= _zz_io_MatrixB_24_18;
    _zz_io_MatrixB_24_20 <= _zz_io_MatrixB_24_19;
    _zz_io_MatrixB_24_21 <= _zz_io_MatrixB_24_20;
    _zz_io_MatrixB_24_22 <= _zz_io_MatrixB_24_21;
    _zz_io_MatrixB_24_23 <= _zz_io_MatrixB_24_22;
    _zz_io_B_Valid_24 <= SubModule_WeightCache_MatrixCol_Switch[24];
    _zz_io_B_Valid_24_1 <= _zz_io_B_Valid_24;
    _zz_io_B_Valid_24_2 <= _zz_io_B_Valid_24_1;
    _zz_io_B_Valid_24_3 <= _zz_io_B_Valid_24_2;
    _zz_io_B_Valid_24_4 <= _zz_io_B_Valid_24_3;
    _zz_io_B_Valid_24_5 <= _zz_io_B_Valid_24_4;
    _zz_io_B_Valid_24_6 <= _zz_io_B_Valid_24_5;
    _zz_io_B_Valid_24_7 <= _zz_io_B_Valid_24_6;
    _zz_io_B_Valid_24_8 <= _zz_io_B_Valid_24_7;
    _zz_io_B_Valid_24_9 <= _zz_io_B_Valid_24_8;
    _zz_io_B_Valid_24_10 <= _zz_io_B_Valid_24_9;
    _zz_io_B_Valid_24_11 <= _zz_io_B_Valid_24_10;
    _zz_io_B_Valid_24_12 <= _zz_io_B_Valid_24_11;
    _zz_io_B_Valid_24_13 <= _zz_io_B_Valid_24_12;
    _zz_io_B_Valid_24_14 <= _zz_io_B_Valid_24_13;
    _zz_io_B_Valid_24_15 <= _zz_io_B_Valid_24_14;
    _zz_io_B_Valid_24_16 <= _zz_io_B_Valid_24_15;
    _zz_io_B_Valid_24_17 <= _zz_io_B_Valid_24_16;
    _zz_io_B_Valid_24_18 <= _zz_io_B_Valid_24_17;
    _zz_io_B_Valid_24_19 <= _zz_io_B_Valid_24_18;
    _zz_io_B_Valid_24_20 <= _zz_io_B_Valid_24_19;
    _zz_io_B_Valid_24_21 <= _zz_io_B_Valid_24_20;
    _zz_io_B_Valid_24_22 <= _zz_io_B_Valid_24_21;
    _zz_io_B_Valid_24_23 <= _zz_io_B_Valid_24_22;
    _zz_io_MatrixB_25 <= SubModule_WeightCache_mData_25;
    _zz_io_MatrixB_25_1 <= _zz_io_MatrixB_25;
    _zz_io_MatrixB_25_2 <= _zz_io_MatrixB_25_1;
    _zz_io_MatrixB_25_3 <= _zz_io_MatrixB_25_2;
    _zz_io_MatrixB_25_4 <= _zz_io_MatrixB_25_3;
    _zz_io_MatrixB_25_5 <= _zz_io_MatrixB_25_4;
    _zz_io_MatrixB_25_6 <= _zz_io_MatrixB_25_5;
    _zz_io_MatrixB_25_7 <= _zz_io_MatrixB_25_6;
    _zz_io_MatrixB_25_8 <= _zz_io_MatrixB_25_7;
    _zz_io_MatrixB_25_9 <= _zz_io_MatrixB_25_8;
    _zz_io_MatrixB_25_10 <= _zz_io_MatrixB_25_9;
    _zz_io_MatrixB_25_11 <= _zz_io_MatrixB_25_10;
    _zz_io_MatrixB_25_12 <= _zz_io_MatrixB_25_11;
    _zz_io_MatrixB_25_13 <= _zz_io_MatrixB_25_12;
    _zz_io_MatrixB_25_14 <= _zz_io_MatrixB_25_13;
    _zz_io_MatrixB_25_15 <= _zz_io_MatrixB_25_14;
    _zz_io_MatrixB_25_16 <= _zz_io_MatrixB_25_15;
    _zz_io_MatrixB_25_17 <= _zz_io_MatrixB_25_16;
    _zz_io_MatrixB_25_18 <= _zz_io_MatrixB_25_17;
    _zz_io_MatrixB_25_19 <= _zz_io_MatrixB_25_18;
    _zz_io_MatrixB_25_20 <= _zz_io_MatrixB_25_19;
    _zz_io_MatrixB_25_21 <= _zz_io_MatrixB_25_20;
    _zz_io_MatrixB_25_22 <= _zz_io_MatrixB_25_21;
    _zz_io_MatrixB_25_23 <= _zz_io_MatrixB_25_22;
    _zz_io_MatrixB_25_24 <= _zz_io_MatrixB_25_23;
    _zz_io_B_Valid_25 <= SubModule_WeightCache_MatrixCol_Switch[25];
    _zz_io_B_Valid_25_1 <= _zz_io_B_Valid_25;
    _zz_io_B_Valid_25_2 <= _zz_io_B_Valid_25_1;
    _zz_io_B_Valid_25_3 <= _zz_io_B_Valid_25_2;
    _zz_io_B_Valid_25_4 <= _zz_io_B_Valid_25_3;
    _zz_io_B_Valid_25_5 <= _zz_io_B_Valid_25_4;
    _zz_io_B_Valid_25_6 <= _zz_io_B_Valid_25_5;
    _zz_io_B_Valid_25_7 <= _zz_io_B_Valid_25_6;
    _zz_io_B_Valid_25_8 <= _zz_io_B_Valid_25_7;
    _zz_io_B_Valid_25_9 <= _zz_io_B_Valid_25_8;
    _zz_io_B_Valid_25_10 <= _zz_io_B_Valid_25_9;
    _zz_io_B_Valid_25_11 <= _zz_io_B_Valid_25_10;
    _zz_io_B_Valid_25_12 <= _zz_io_B_Valid_25_11;
    _zz_io_B_Valid_25_13 <= _zz_io_B_Valid_25_12;
    _zz_io_B_Valid_25_14 <= _zz_io_B_Valid_25_13;
    _zz_io_B_Valid_25_15 <= _zz_io_B_Valid_25_14;
    _zz_io_B_Valid_25_16 <= _zz_io_B_Valid_25_15;
    _zz_io_B_Valid_25_17 <= _zz_io_B_Valid_25_16;
    _zz_io_B_Valid_25_18 <= _zz_io_B_Valid_25_17;
    _zz_io_B_Valid_25_19 <= _zz_io_B_Valid_25_18;
    _zz_io_B_Valid_25_20 <= _zz_io_B_Valid_25_19;
    _zz_io_B_Valid_25_21 <= _zz_io_B_Valid_25_20;
    _zz_io_B_Valid_25_22 <= _zz_io_B_Valid_25_21;
    _zz_io_B_Valid_25_23 <= _zz_io_B_Valid_25_22;
    _zz_io_B_Valid_25_24 <= _zz_io_B_Valid_25_23;
    _zz_io_MatrixB_26 <= SubModule_WeightCache_mData_26;
    _zz_io_MatrixB_26_1 <= _zz_io_MatrixB_26;
    _zz_io_MatrixB_26_2 <= _zz_io_MatrixB_26_1;
    _zz_io_MatrixB_26_3 <= _zz_io_MatrixB_26_2;
    _zz_io_MatrixB_26_4 <= _zz_io_MatrixB_26_3;
    _zz_io_MatrixB_26_5 <= _zz_io_MatrixB_26_4;
    _zz_io_MatrixB_26_6 <= _zz_io_MatrixB_26_5;
    _zz_io_MatrixB_26_7 <= _zz_io_MatrixB_26_6;
    _zz_io_MatrixB_26_8 <= _zz_io_MatrixB_26_7;
    _zz_io_MatrixB_26_9 <= _zz_io_MatrixB_26_8;
    _zz_io_MatrixB_26_10 <= _zz_io_MatrixB_26_9;
    _zz_io_MatrixB_26_11 <= _zz_io_MatrixB_26_10;
    _zz_io_MatrixB_26_12 <= _zz_io_MatrixB_26_11;
    _zz_io_MatrixB_26_13 <= _zz_io_MatrixB_26_12;
    _zz_io_MatrixB_26_14 <= _zz_io_MatrixB_26_13;
    _zz_io_MatrixB_26_15 <= _zz_io_MatrixB_26_14;
    _zz_io_MatrixB_26_16 <= _zz_io_MatrixB_26_15;
    _zz_io_MatrixB_26_17 <= _zz_io_MatrixB_26_16;
    _zz_io_MatrixB_26_18 <= _zz_io_MatrixB_26_17;
    _zz_io_MatrixB_26_19 <= _zz_io_MatrixB_26_18;
    _zz_io_MatrixB_26_20 <= _zz_io_MatrixB_26_19;
    _zz_io_MatrixB_26_21 <= _zz_io_MatrixB_26_20;
    _zz_io_MatrixB_26_22 <= _zz_io_MatrixB_26_21;
    _zz_io_MatrixB_26_23 <= _zz_io_MatrixB_26_22;
    _zz_io_MatrixB_26_24 <= _zz_io_MatrixB_26_23;
    _zz_io_MatrixB_26_25 <= _zz_io_MatrixB_26_24;
    _zz_io_B_Valid_26 <= SubModule_WeightCache_MatrixCol_Switch[26];
    _zz_io_B_Valid_26_1 <= _zz_io_B_Valid_26;
    _zz_io_B_Valid_26_2 <= _zz_io_B_Valid_26_1;
    _zz_io_B_Valid_26_3 <= _zz_io_B_Valid_26_2;
    _zz_io_B_Valid_26_4 <= _zz_io_B_Valid_26_3;
    _zz_io_B_Valid_26_5 <= _zz_io_B_Valid_26_4;
    _zz_io_B_Valid_26_6 <= _zz_io_B_Valid_26_5;
    _zz_io_B_Valid_26_7 <= _zz_io_B_Valid_26_6;
    _zz_io_B_Valid_26_8 <= _zz_io_B_Valid_26_7;
    _zz_io_B_Valid_26_9 <= _zz_io_B_Valid_26_8;
    _zz_io_B_Valid_26_10 <= _zz_io_B_Valid_26_9;
    _zz_io_B_Valid_26_11 <= _zz_io_B_Valid_26_10;
    _zz_io_B_Valid_26_12 <= _zz_io_B_Valid_26_11;
    _zz_io_B_Valid_26_13 <= _zz_io_B_Valid_26_12;
    _zz_io_B_Valid_26_14 <= _zz_io_B_Valid_26_13;
    _zz_io_B_Valid_26_15 <= _zz_io_B_Valid_26_14;
    _zz_io_B_Valid_26_16 <= _zz_io_B_Valid_26_15;
    _zz_io_B_Valid_26_17 <= _zz_io_B_Valid_26_16;
    _zz_io_B_Valid_26_18 <= _zz_io_B_Valid_26_17;
    _zz_io_B_Valid_26_19 <= _zz_io_B_Valid_26_18;
    _zz_io_B_Valid_26_20 <= _zz_io_B_Valid_26_19;
    _zz_io_B_Valid_26_21 <= _zz_io_B_Valid_26_20;
    _zz_io_B_Valid_26_22 <= _zz_io_B_Valid_26_21;
    _zz_io_B_Valid_26_23 <= _zz_io_B_Valid_26_22;
    _zz_io_B_Valid_26_24 <= _zz_io_B_Valid_26_23;
    _zz_io_B_Valid_26_25 <= _zz_io_B_Valid_26_24;
    _zz_io_MatrixB_27 <= SubModule_WeightCache_mData_27;
    _zz_io_MatrixB_27_1 <= _zz_io_MatrixB_27;
    _zz_io_MatrixB_27_2 <= _zz_io_MatrixB_27_1;
    _zz_io_MatrixB_27_3 <= _zz_io_MatrixB_27_2;
    _zz_io_MatrixB_27_4 <= _zz_io_MatrixB_27_3;
    _zz_io_MatrixB_27_5 <= _zz_io_MatrixB_27_4;
    _zz_io_MatrixB_27_6 <= _zz_io_MatrixB_27_5;
    _zz_io_MatrixB_27_7 <= _zz_io_MatrixB_27_6;
    _zz_io_MatrixB_27_8 <= _zz_io_MatrixB_27_7;
    _zz_io_MatrixB_27_9 <= _zz_io_MatrixB_27_8;
    _zz_io_MatrixB_27_10 <= _zz_io_MatrixB_27_9;
    _zz_io_MatrixB_27_11 <= _zz_io_MatrixB_27_10;
    _zz_io_MatrixB_27_12 <= _zz_io_MatrixB_27_11;
    _zz_io_MatrixB_27_13 <= _zz_io_MatrixB_27_12;
    _zz_io_MatrixB_27_14 <= _zz_io_MatrixB_27_13;
    _zz_io_MatrixB_27_15 <= _zz_io_MatrixB_27_14;
    _zz_io_MatrixB_27_16 <= _zz_io_MatrixB_27_15;
    _zz_io_MatrixB_27_17 <= _zz_io_MatrixB_27_16;
    _zz_io_MatrixB_27_18 <= _zz_io_MatrixB_27_17;
    _zz_io_MatrixB_27_19 <= _zz_io_MatrixB_27_18;
    _zz_io_MatrixB_27_20 <= _zz_io_MatrixB_27_19;
    _zz_io_MatrixB_27_21 <= _zz_io_MatrixB_27_20;
    _zz_io_MatrixB_27_22 <= _zz_io_MatrixB_27_21;
    _zz_io_MatrixB_27_23 <= _zz_io_MatrixB_27_22;
    _zz_io_MatrixB_27_24 <= _zz_io_MatrixB_27_23;
    _zz_io_MatrixB_27_25 <= _zz_io_MatrixB_27_24;
    _zz_io_MatrixB_27_26 <= _zz_io_MatrixB_27_25;
    _zz_io_B_Valid_27 <= SubModule_WeightCache_MatrixCol_Switch[27];
    _zz_io_B_Valid_27_1 <= _zz_io_B_Valid_27;
    _zz_io_B_Valid_27_2 <= _zz_io_B_Valid_27_1;
    _zz_io_B_Valid_27_3 <= _zz_io_B_Valid_27_2;
    _zz_io_B_Valid_27_4 <= _zz_io_B_Valid_27_3;
    _zz_io_B_Valid_27_5 <= _zz_io_B_Valid_27_4;
    _zz_io_B_Valid_27_6 <= _zz_io_B_Valid_27_5;
    _zz_io_B_Valid_27_7 <= _zz_io_B_Valid_27_6;
    _zz_io_B_Valid_27_8 <= _zz_io_B_Valid_27_7;
    _zz_io_B_Valid_27_9 <= _zz_io_B_Valid_27_8;
    _zz_io_B_Valid_27_10 <= _zz_io_B_Valid_27_9;
    _zz_io_B_Valid_27_11 <= _zz_io_B_Valid_27_10;
    _zz_io_B_Valid_27_12 <= _zz_io_B_Valid_27_11;
    _zz_io_B_Valid_27_13 <= _zz_io_B_Valid_27_12;
    _zz_io_B_Valid_27_14 <= _zz_io_B_Valid_27_13;
    _zz_io_B_Valid_27_15 <= _zz_io_B_Valid_27_14;
    _zz_io_B_Valid_27_16 <= _zz_io_B_Valid_27_15;
    _zz_io_B_Valid_27_17 <= _zz_io_B_Valid_27_16;
    _zz_io_B_Valid_27_18 <= _zz_io_B_Valid_27_17;
    _zz_io_B_Valid_27_19 <= _zz_io_B_Valid_27_18;
    _zz_io_B_Valid_27_20 <= _zz_io_B_Valid_27_19;
    _zz_io_B_Valid_27_21 <= _zz_io_B_Valid_27_20;
    _zz_io_B_Valid_27_22 <= _zz_io_B_Valid_27_21;
    _zz_io_B_Valid_27_23 <= _zz_io_B_Valid_27_22;
    _zz_io_B_Valid_27_24 <= _zz_io_B_Valid_27_23;
    _zz_io_B_Valid_27_25 <= _zz_io_B_Valid_27_24;
    _zz_io_B_Valid_27_26 <= _zz_io_B_Valid_27_25;
    _zz_io_MatrixB_28 <= SubModule_WeightCache_mData_28;
    _zz_io_MatrixB_28_1 <= _zz_io_MatrixB_28;
    _zz_io_MatrixB_28_2 <= _zz_io_MatrixB_28_1;
    _zz_io_MatrixB_28_3 <= _zz_io_MatrixB_28_2;
    _zz_io_MatrixB_28_4 <= _zz_io_MatrixB_28_3;
    _zz_io_MatrixB_28_5 <= _zz_io_MatrixB_28_4;
    _zz_io_MatrixB_28_6 <= _zz_io_MatrixB_28_5;
    _zz_io_MatrixB_28_7 <= _zz_io_MatrixB_28_6;
    _zz_io_MatrixB_28_8 <= _zz_io_MatrixB_28_7;
    _zz_io_MatrixB_28_9 <= _zz_io_MatrixB_28_8;
    _zz_io_MatrixB_28_10 <= _zz_io_MatrixB_28_9;
    _zz_io_MatrixB_28_11 <= _zz_io_MatrixB_28_10;
    _zz_io_MatrixB_28_12 <= _zz_io_MatrixB_28_11;
    _zz_io_MatrixB_28_13 <= _zz_io_MatrixB_28_12;
    _zz_io_MatrixB_28_14 <= _zz_io_MatrixB_28_13;
    _zz_io_MatrixB_28_15 <= _zz_io_MatrixB_28_14;
    _zz_io_MatrixB_28_16 <= _zz_io_MatrixB_28_15;
    _zz_io_MatrixB_28_17 <= _zz_io_MatrixB_28_16;
    _zz_io_MatrixB_28_18 <= _zz_io_MatrixB_28_17;
    _zz_io_MatrixB_28_19 <= _zz_io_MatrixB_28_18;
    _zz_io_MatrixB_28_20 <= _zz_io_MatrixB_28_19;
    _zz_io_MatrixB_28_21 <= _zz_io_MatrixB_28_20;
    _zz_io_MatrixB_28_22 <= _zz_io_MatrixB_28_21;
    _zz_io_MatrixB_28_23 <= _zz_io_MatrixB_28_22;
    _zz_io_MatrixB_28_24 <= _zz_io_MatrixB_28_23;
    _zz_io_MatrixB_28_25 <= _zz_io_MatrixB_28_24;
    _zz_io_MatrixB_28_26 <= _zz_io_MatrixB_28_25;
    _zz_io_MatrixB_28_27 <= _zz_io_MatrixB_28_26;
    _zz_io_B_Valid_28 <= SubModule_WeightCache_MatrixCol_Switch[28];
    _zz_io_B_Valid_28_1 <= _zz_io_B_Valid_28;
    _zz_io_B_Valid_28_2 <= _zz_io_B_Valid_28_1;
    _zz_io_B_Valid_28_3 <= _zz_io_B_Valid_28_2;
    _zz_io_B_Valid_28_4 <= _zz_io_B_Valid_28_3;
    _zz_io_B_Valid_28_5 <= _zz_io_B_Valid_28_4;
    _zz_io_B_Valid_28_6 <= _zz_io_B_Valid_28_5;
    _zz_io_B_Valid_28_7 <= _zz_io_B_Valid_28_6;
    _zz_io_B_Valid_28_8 <= _zz_io_B_Valid_28_7;
    _zz_io_B_Valid_28_9 <= _zz_io_B_Valid_28_8;
    _zz_io_B_Valid_28_10 <= _zz_io_B_Valid_28_9;
    _zz_io_B_Valid_28_11 <= _zz_io_B_Valid_28_10;
    _zz_io_B_Valid_28_12 <= _zz_io_B_Valid_28_11;
    _zz_io_B_Valid_28_13 <= _zz_io_B_Valid_28_12;
    _zz_io_B_Valid_28_14 <= _zz_io_B_Valid_28_13;
    _zz_io_B_Valid_28_15 <= _zz_io_B_Valid_28_14;
    _zz_io_B_Valid_28_16 <= _zz_io_B_Valid_28_15;
    _zz_io_B_Valid_28_17 <= _zz_io_B_Valid_28_16;
    _zz_io_B_Valid_28_18 <= _zz_io_B_Valid_28_17;
    _zz_io_B_Valid_28_19 <= _zz_io_B_Valid_28_18;
    _zz_io_B_Valid_28_20 <= _zz_io_B_Valid_28_19;
    _zz_io_B_Valid_28_21 <= _zz_io_B_Valid_28_20;
    _zz_io_B_Valid_28_22 <= _zz_io_B_Valid_28_21;
    _zz_io_B_Valid_28_23 <= _zz_io_B_Valid_28_22;
    _zz_io_B_Valid_28_24 <= _zz_io_B_Valid_28_23;
    _zz_io_B_Valid_28_25 <= _zz_io_B_Valid_28_24;
    _zz_io_B_Valid_28_26 <= _zz_io_B_Valid_28_25;
    _zz_io_B_Valid_28_27 <= _zz_io_B_Valid_28_26;
    _zz_io_MatrixB_29 <= SubModule_WeightCache_mData_29;
    _zz_io_MatrixB_29_1 <= _zz_io_MatrixB_29;
    _zz_io_MatrixB_29_2 <= _zz_io_MatrixB_29_1;
    _zz_io_MatrixB_29_3 <= _zz_io_MatrixB_29_2;
    _zz_io_MatrixB_29_4 <= _zz_io_MatrixB_29_3;
    _zz_io_MatrixB_29_5 <= _zz_io_MatrixB_29_4;
    _zz_io_MatrixB_29_6 <= _zz_io_MatrixB_29_5;
    _zz_io_MatrixB_29_7 <= _zz_io_MatrixB_29_6;
    _zz_io_MatrixB_29_8 <= _zz_io_MatrixB_29_7;
    _zz_io_MatrixB_29_9 <= _zz_io_MatrixB_29_8;
    _zz_io_MatrixB_29_10 <= _zz_io_MatrixB_29_9;
    _zz_io_MatrixB_29_11 <= _zz_io_MatrixB_29_10;
    _zz_io_MatrixB_29_12 <= _zz_io_MatrixB_29_11;
    _zz_io_MatrixB_29_13 <= _zz_io_MatrixB_29_12;
    _zz_io_MatrixB_29_14 <= _zz_io_MatrixB_29_13;
    _zz_io_MatrixB_29_15 <= _zz_io_MatrixB_29_14;
    _zz_io_MatrixB_29_16 <= _zz_io_MatrixB_29_15;
    _zz_io_MatrixB_29_17 <= _zz_io_MatrixB_29_16;
    _zz_io_MatrixB_29_18 <= _zz_io_MatrixB_29_17;
    _zz_io_MatrixB_29_19 <= _zz_io_MatrixB_29_18;
    _zz_io_MatrixB_29_20 <= _zz_io_MatrixB_29_19;
    _zz_io_MatrixB_29_21 <= _zz_io_MatrixB_29_20;
    _zz_io_MatrixB_29_22 <= _zz_io_MatrixB_29_21;
    _zz_io_MatrixB_29_23 <= _zz_io_MatrixB_29_22;
    _zz_io_MatrixB_29_24 <= _zz_io_MatrixB_29_23;
    _zz_io_MatrixB_29_25 <= _zz_io_MatrixB_29_24;
    _zz_io_MatrixB_29_26 <= _zz_io_MatrixB_29_25;
    _zz_io_MatrixB_29_27 <= _zz_io_MatrixB_29_26;
    _zz_io_MatrixB_29_28 <= _zz_io_MatrixB_29_27;
    _zz_io_B_Valid_29 <= SubModule_WeightCache_MatrixCol_Switch[29];
    _zz_io_B_Valid_29_1 <= _zz_io_B_Valid_29;
    _zz_io_B_Valid_29_2 <= _zz_io_B_Valid_29_1;
    _zz_io_B_Valid_29_3 <= _zz_io_B_Valid_29_2;
    _zz_io_B_Valid_29_4 <= _zz_io_B_Valid_29_3;
    _zz_io_B_Valid_29_5 <= _zz_io_B_Valid_29_4;
    _zz_io_B_Valid_29_6 <= _zz_io_B_Valid_29_5;
    _zz_io_B_Valid_29_7 <= _zz_io_B_Valid_29_6;
    _zz_io_B_Valid_29_8 <= _zz_io_B_Valid_29_7;
    _zz_io_B_Valid_29_9 <= _zz_io_B_Valid_29_8;
    _zz_io_B_Valid_29_10 <= _zz_io_B_Valid_29_9;
    _zz_io_B_Valid_29_11 <= _zz_io_B_Valid_29_10;
    _zz_io_B_Valid_29_12 <= _zz_io_B_Valid_29_11;
    _zz_io_B_Valid_29_13 <= _zz_io_B_Valid_29_12;
    _zz_io_B_Valid_29_14 <= _zz_io_B_Valid_29_13;
    _zz_io_B_Valid_29_15 <= _zz_io_B_Valid_29_14;
    _zz_io_B_Valid_29_16 <= _zz_io_B_Valid_29_15;
    _zz_io_B_Valid_29_17 <= _zz_io_B_Valid_29_16;
    _zz_io_B_Valid_29_18 <= _zz_io_B_Valid_29_17;
    _zz_io_B_Valid_29_19 <= _zz_io_B_Valid_29_18;
    _zz_io_B_Valid_29_20 <= _zz_io_B_Valid_29_19;
    _zz_io_B_Valid_29_21 <= _zz_io_B_Valid_29_20;
    _zz_io_B_Valid_29_22 <= _zz_io_B_Valid_29_21;
    _zz_io_B_Valid_29_23 <= _zz_io_B_Valid_29_22;
    _zz_io_B_Valid_29_24 <= _zz_io_B_Valid_29_23;
    _zz_io_B_Valid_29_25 <= _zz_io_B_Valid_29_24;
    _zz_io_B_Valid_29_26 <= _zz_io_B_Valid_29_25;
    _zz_io_B_Valid_29_27 <= _zz_io_B_Valid_29_26;
    _zz_io_B_Valid_29_28 <= _zz_io_B_Valid_29_27;
    _zz_io_MatrixB_30 <= SubModule_WeightCache_mData_30;
    _zz_io_MatrixB_30_1 <= _zz_io_MatrixB_30;
    _zz_io_MatrixB_30_2 <= _zz_io_MatrixB_30_1;
    _zz_io_MatrixB_30_3 <= _zz_io_MatrixB_30_2;
    _zz_io_MatrixB_30_4 <= _zz_io_MatrixB_30_3;
    _zz_io_MatrixB_30_5 <= _zz_io_MatrixB_30_4;
    _zz_io_MatrixB_30_6 <= _zz_io_MatrixB_30_5;
    _zz_io_MatrixB_30_7 <= _zz_io_MatrixB_30_6;
    _zz_io_MatrixB_30_8 <= _zz_io_MatrixB_30_7;
    _zz_io_MatrixB_30_9 <= _zz_io_MatrixB_30_8;
    _zz_io_MatrixB_30_10 <= _zz_io_MatrixB_30_9;
    _zz_io_MatrixB_30_11 <= _zz_io_MatrixB_30_10;
    _zz_io_MatrixB_30_12 <= _zz_io_MatrixB_30_11;
    _zz_io_MatrixB_30_13 <= _zz_io_MatrixB_30_12;
    _zz_io_MatrixB_30_14 <= _zz_io_MatrixB_30_13;
    _zz_io_MatrixB_30_15 <= _zz_io_MatrixB_30_14;
    _zz_io_MatrixB_30_16 <= _zz_io_MatrixB_30_15;
    _zz_io_MatrixB_30_17 <= _zz_io_MatrixB_30_16;
    _zz_io_MatrixB_30_18 <= _zz_io_MatrixB_30_17;
    _zz_io_MatrixB_30_19 <= _zz_io_MatrixB_30_18;
    _zz_io_MatrixB_30_20 <= _zz_io_MatrixB_30_19;
    _zz_io_MatrixB_30_21 <= _zz_io_MatrixB_30_20;
    _zz_io_MatrixB_30_22 <= _zz_io_MatrixB_30_21;
    _zz_io_MatrixB_30_23 <= _zz_io_MatrixB_30_22;
    _zz_io_MatrixB_30_24 <= _zz_io_MatrixB_30_23;
    _zz_io_MatrixB_30_25 <= _zz_io_MatrixB_30_24;
    _zz_io_MatrixB_30_26 <= _zz_io_MatrixB_30_25;
    _zz_io_MatrixB_30_27 <= _zz_io_MatrixB_30_26;
    _zz_io_MatrixB_30_28 <= _zz_io_MatrixB_30_27;
    _zz_io_MatrixB_30_29 <= _zz_io_MatrixB_30_28;
    _zz_io_B_Valid_30 <= SubModule_WeightCache_MatrixCol_Switch[30];
    _zz_io_B_Valid_30_1 <= _zz_io_B_Valid_30;
    _zz_io_B_Valid_30_2 <= _zz_io_B_Valid_30_1;
    _zz_io_B_Valid_30_3 <= _zz_io_B_Valid_30_2;
    _zz_io_B_Valid_30_4 <= _zz_io_B_Valid_30_3;
    _zz_io_B_Valid_30_5 <= _zz_io_B_Valid_30_4;
    _zz_io_B_Valid_30_6 <= _zz_io_B_Valid_30_5;
    _zz_io_B_Valid_30_7 <= _zz_io_B_Valid_30_6;
    _zz_io_B_Valid_30_8 <= _zz_io_B_Valid_30_7;
    _zz_io_B_Valid_30_9 <= _zz_io_B_Valid_30_8;
    _zz_io_B_Valid_30_10 <= _zz_io_B_Valid_30_9;
    _zz_io_B_Valid_30_11 <= _zz_io_B_Valid_30_10;
    _zz_io_B_Valid_30_12 <= _zz_io_B_Valid_30_11;
    _zz_io_B_Valid_30_13 <= _zz_io_B_Valid_30_12;
    _zz_io_B_Valid_30_14 <= _zz_io_B_Valid_30_13;
    _zz_io_B_Valid_30_15 <= _zz_io_B_Valid_30_14;
    _zz_io_B_Valid_30_16 <= _zz_io_B_Valid_30_15;
    _zz_io_B_Valid_30_17 <= _zz_io_B_Valid_30_16;
    _zz_io_B_Valid_30_18 <= _zz_io_B_Valid_30_17;
    _zz_io_B_Valid_30_19 <= _zz_io_B_Valid_30_18;
    _zz_io_B_Valid_30_20 <= _zz_io_B_Valid_30_19;
    _zz_io_B_Valid_30_21 <= _zz_io_B_Valid_30_20;
    _zz_io_B_Valid_30_22 <= _zz_io_B_Valid_30_21;
    _zz_io_B_Valid_30_23 <= _zz_io_B_Valid_30_22;
    _zz_io_B_Valid_30_24 <= _zz_io_B_Valid_30_23;
    _zz_io_B_Valid_30_25 <= _zz_io_B_Valid_30_24;
    _zz_io_B_Valid_30_26 <= _zz_io_B_Valid_30_25;
    _zz_io_B_Valid_30_27 <= _zz_io_B_Valid_30_26;
    _zz_io_B_Valid_30_28 <= _zz_io_B_Valid_30_27;
    _zz_io_B_Valid_30_29 <= _zz_io_B_Valid_30_28;
    _zz_io_MatrixB_31 <= SubModule_WeightCache_mData_31;
    _zz_io_MatrixB_31_1 <= _zz_io_MatrixB_31;
    _zz_io_MatrixB_31_2 <= _zz_io_MatrixB_31_1;
    _zz_io_MatrixB_31_3 <= _zz_io_MatrixB_31_2;
    _zz_io_MatrixB_31_4 <= _zz_io_MatrixB_31_3;
    _zz_io_MatrixB_31_5 <= _zz_io_MatrixB_31_4;
    _zz_io_MatrixB_31_6 <= _zz_io_MatrixB_31_5;
    _zz_io_MatrixB_31_7 <= _zz_io_MatrixB_31_6;
    _zz_io_MatrixB_31_8 <= _zz_io_MatrixB_31_7;
    _zz_io_MatrixB_31_9 <= _zz_io_MatrixB_31_8;
    _zz_io_MatrixB_31_10 <= _zz_io_MatrixB_31_9;
    _zz_io_MatrixB_31_11 <= _zz_io_MatrixB_31_10;
    _zz_io_MatrixB_31_12 <= _zz_io_MatrixB_31_11;
    _zz_io_MatrixB_31_13 <= _zz_io_MatrixB_31_12;
    _zz_io_MatrixB_31_14 <= _zz_io_MatrixB_31_13;
    _zz_io_MatrixB_31_15 <= _zz_io_MatrixB_31_14;
    _zz_io_MatrixB_31_16 <= _zz_io_MatrixB_31_15;
    _zz_io_MatrixB_31_17 <= _zz_io_MatrixB_31_16;
    _zz_io_MatrixB_31_18 <= _zz_io_MatrixB_31_17;
    _zz_io_MatrixB_31_19 <= _zz_io_MatrixB_31_18;
    _zz_io_MatrixB_31_20 <= _zz_io_MatrixB_31_19;
    _zz_io_MatrixB_31_21 <= _zz_io_MatrixB_31_20;
    _zz_io_MatrixB_31_22 <= _zz_io_MatrixB_31_21;
    _zz_io_MatrixB_31_23 <= _zz_io_MatrixB_31_22;
    _zz_io_MatrixB_31_24 <= _zz_io_MatrixB_31_23;
    _zz_io_MatrixB_31_25 <= _zz_io_MatrixB_31_24;
    _zz_io_MatrixB_31_26 <= _zz_io_MatrixB_31_25;
    _zz_io_MatrixB_31_27 <= _zz_io_MatrixB_31_26;
    _zz_io_MatrixB_31_28 <= _zz_io_MatrixB_31_27;
    _zz_io_MatrixB_31_29 <= _zz_io_MatrixB_31_28;
    _zz_io_MatrixB_31_30 <= _zz_io_MatrixB_31_29;
    _zz_io_B_Valid_31 <= SubModule_WeightCache_MatrixCol_Switch[31];
    _zz_io_B_Valid_31_1 <= _zz_io_B_Valid_31;
    _zz_io_B_Valid_31_2 <= _zz_io_B_Valid_31_1;
    _zz_io_B_Valid_31_3 <= _zz_io_B_Valid_31_2;
    _zz_io_B_Valid_31_4 <= _zz_io_B_Valid_31_3;
    _zz_io_B_Valid_31_5 <= _zz_io_B_Valid_31_4;
    _zz_io_B_Valid_31_6 <= _zz_io_B_Valid_31_5;
    _zz_io_B_Valid_31_7 <= _zz_io_B_Valid_31_6;
    _zz_io_B_Valid_31_8 <= _zz_io_B_Valid_31_7;
    _zz_io_B_Valid_31_9 <= _zz_io_B_Valid_31_8;
    _zz_io_B_Valid_31_10 <= _zz_io_B_Valid_31_9;
    _zz_io_B_Valid_31_11 <= _zz_io_B_Valid_31_10;
    _zz_io_B_Valid_31_12 <= _zz_io_B_Valid_31_11;
    _zz_io_B_Valid_31_13 <= _zz_io_B_Valid_31_12;
    _zz_io_B_Valid_31_14 <= _zz_io_B_Valid_31_13;
    _zz_io_B_Valid_31_15 <= _zz_io_B_Valid_31_14;
    _zz_io_B_Valid_31_16 <= _zz_io_B_Valid_31_15;
    _zz_io_B_Valid_31_17 <= _zz_io_B_Valid_31_16;
    _zz_io_B_Valid_31_18 <= _zz_io_B_Valid_31_17;
    _zz_io_B_Valid_31_19 <= _zz_io_B_Valid_31_18;
    _zz_io_B_Valid_31_20 <= _zz_io_B_Valid_31_19;
    _zz_io_B_Valid_31_21 <= _zz_io_B_Valid_31_20;
    _zz_io_B_Valid_31_22 <= _zz_io_B_Valid_31_21;
    _zz_io_B_Valid_31_23 <= _zz_io_B_Valid_31_22;
    _zz_io_B_Valid_31_24 <= _zz_io_B_Valid_31_23;
    _zz_io_B_Valid_31_25 <= _zz_io_B_Valid_31_24;
    _zz_io_B_Valid_31_26 <= _zz_io_B_Valid_31_25;
    _zz_io_B_Valid_31_27 <= _zz_io_B_Valid_31_26;
    _zz_io_B_Valid_31_28 <= _zz_io_B_Valid_31_27;
    _zz_io_B_Valid_31_29 <= _zz_io_B_Valid_31_28;
    _zz_io_B_Valid_31_30 <= _zz_io_B_Valid_31_29;
    _zz_io_MatrixB_32 <= SubModule_WeightCache_mData_32;
    _zz_io_MatrixB_32_1 <= _zz_io_MatrixB_32;
    _zz_io_MatrixB_32_2 <= _zz_io_MatrixB_32_1;
    _zz_io_MatrixB_32_3 <= _zz_io_MatrixB_32_2;
    _zz_io_MatrixB_32_4 <= _zz_io_MatrixB_32_3;
    _zz_io_MatrixB_32_5 <= _zz_io_MatrixB_32_4;
    _zz_io_MatrixB_32_6 <= _zz_io_MatrixB_32_5;
    _zz_io_MatrixB_32_7 <= _zz_io_MatrixB_32_6;
    _zz_io_MatrixB_32_8 <= _zz_io_MatrixB_32_7;
    _zz_io_MatrixB_32_9 <= _zz_io_MatrixB_32_8;
    _zz_io_MatrixB_32_10 <= _zz_io_MatrixB_32_9;
    _zz_io_MatrixB_32_11 <= _zz_io_MatrixB_32_10;
    _zz_io_MatrixB_32_12 <= _zz_io_MatrixB_32_11;
    _zz_io_MatrixB_32_13 <= _zz_io_MatrixB_32_12;
    _zz_io_MatrixB_32_14 <= _zz_io_MatrixB_32_13;
    _zz_io_MatrixB_32_15 <= _zz_io_MatrixB_32_14;
    _zz_io_MatrixB_32_16 <= _zz_io_MatrixB_32_15;
    _zz_io_MatrixB_32_17 <= _zz_io_MatrixB_32_16;
    _zz_io_MatrixB_32_18 <= _zz_io_MatrixB_32_17;
    _zz_io_MatrixB_32_19 <= _zz_io_MatrixB_32_18;
    _zz_io_MatrixB_32_20 <= _zz_io_MatrixB_32_19;
    _zz_io_MatrixB_32_21 <= _zz_io_MatrixB_32_20;
    _zz_io_MatrixB_32_22 <= _zz_io_MatrixB_32_21;
    _zz_io_MatrixB_32_23 <= _zz_io_MatrixB_32_22;
    _zz_io_MatrixB_32_24 <= _zz_io_MatrixB_32_23;
    _zz_io_MatrixB_32_25 <= _zz_io_MatrixB_32_24;
    _zz_io_MatrixB_32_26 <= _zz_io_MatrixB_32_25;
    _zz_io_MatrixB_32_27 <= _zz_io_MatrixB_32_26;
    _zz_io_MatrixB_32_28 <= _zz_io_MatrixB_32_27;
    _zz_io_MatrixB_32_29 <= _zz_io_MatrixB_32_28;
    _zz_io_MatrixB_32_30 <= _zz_io_MatrixB_32_29;
    _zz_io_MatrixB_32_31 <= _zz_io_MatrixB_32_30;
    _zz_io_B_Valid_32 <= SubModule_WeightCache_MatrixCol_Switch[32];
    _zz_io_B_Valid_32_1 <= _zz_io_B_Valid_32;
    _zz_io_B_Valid_32_2 <= _zz_io_B_Valid_32_1;
    _zz_io_B_Valid_32_3 <= _zz_io_B_Valid_32_2;
    _zz_io_B_Valid_32_4 <= _zz_io_B_Valid_32_3;
    _zz_io_B_Valid_32_5 <= _zz_io_B_Valid_32_4;
    _zz_io_B_Valid_32_6 <= _zz_io_B_Valid_32_5;
    _zz_io_B_Valid_32_7 <= _zz_io_B_Valid_32_6;
    _zz_io_B_Valid_32_8 <= _zz_io_B_Valid_32_7;
    _zz_io_B_Valid_32_9 <= _zz_io_B_Valid_32_8;
    _zz_io_B_Valid_32_10 <= _zz_io_B_Valid_32_9;
    _zz_io_B_Valid_32_11 <= _zz_io_B_Valid_32_10;
    _zz_io_B_Valid_32_12 <= _zz_io_B_Valid_32_11;
    _zz_io_B_Valid_32_13 <= _zz_io_B_Valid_32_12;
    _zz_io_B_Valid_32_14 <= _zz_io_B_Valid_32_13;
    _zz_io_B_Valid_32_15 <= _zz_io_B_Valid_32_14;
    _zz_io_B_Valid_32_16 <= _zz_io_B_Valid_32_15;
    _zz_io_B_Valid_32_17 <= _zz_io_B_Valid_32_16;
    _zz_io_B_Valid_32_18 <= _zz_io_B_Valid_32_17;
    _zz_io_B_Valid_32_19 <= _zz_io_B_Valid_32_18;
    _zz_io_B_Valid_32_20 <= _zz_io_B_Valid_32_19;
    _zz_io_B_Valid_32_21 <= _zz_io_B_Valid_32_20;
    _zz_io_B_Valid_32_22 <= _zz_io_B_Valid_32_21;
    _zz_io_B_Valid_32_23 <= _zz_io_B_Valid_32_22;
    _zz_io_B_Valid_32_24 <= _zz_io_B_Valid_32_23;
    _zz_io_B_Valid_32_25 <= _zz_io_B_Valid_32_24;
    _zz_io_B_Valid_32_26 <= _zz_io_B_Valid_32_25;
    _zz_io_B_Valid_32_27 <= _zz_io_B_Valid_32_26;
    _zz_io_B_Valid_32_28 <= _zz_io_B_Valid_32_27;
    _zz_io_B_Valid_32_29 <= _zz_io_B_Valid_32_28;
    _zz_io_B_Valid_32_30 <= _zz_io_B_Valid_32_29;
    _zz_io_B_Valid_32_31 <= _zz_io_B_Valid_32_30;
    _zz_io_MatrixB_33 <= SubModule_WeightCache_mData_33;
    _zz_io_MatrixB_33_1 <= _zz_io_MatrixB_33;
    _zz_io_MatrixB_33_2 <= _zz_io_MatrixB_33_1;
    _zz_io_MatrixB_33_3 <= _zz_io_MatrixB_33_2;
    _zz_io_MatrixB_33_4 <= _zz_io_MatrixB_33_3;
    _zz_io_MatrixB_33_5 <= _zz_io_MatrixB_33_4;
    _zz_io_MatrixB_33_6 <= _zz_io_MatrixB_33_5;
    _zz_io_MatrixB_33_7 <= _zz_io_MatrixB_33_6;
    _zz_io_MatrixB_33_8 <= _zz_io_MatrixB_33_7;
    _zz_io_MatrixB_33_9 <= _zz_io_MatrixB_33_8;
    _zz_io_MatrixB_33_10 <= _zz_io_MatrixB_33_9;
    _zz_io_MatrixB_33_11 <= _zz_io_MatrixB_33_10;
    _zz_io_MatrixB_33_12 <= _zz_io_MatrixB_33_11;
    _zz_io_MatrixB_33_13 <= _zz_io_MatrixB_33_12;
    _zz_io_MatrixB_33_14 <= _zz_io_MatrixB_33_13;
    _zz_io_MatrixB_33_15 <= _zz_io_MatrixB_33_14;
    _zz_io_MatrixB_33_16 <= _zz_io_MatrixB_33_15;
    _zz_io_MatrixB_33_17 <= _zz_io_MatrixB_33_16;
    _zz_io_MatrixB_33_18 <= _zz_io_MatrixB_33_17;
    _zz_io_MatrixB_33_19 <= _zz_io_MatrixB_33_18;
    _zz_io_MatrixB_33_20 <= _zz_io_MatrixB_33_19;
    _zz_io_MatrixB_33_21 <= _zz_io_MatrixB_33_20;
    _zz_io_MatrixB_33_22 <= _zz_io_MatrixB_33_21;
    _zz_io_MatrixB_33_23 <= _zz_io_MatrixB_33_22;
    _zz_io_MatrixB_33_24 <= _zz_io_MatrixB_33_23;
    _zz_io_MatrixB_33_25 <= _zz_io_MatrixB_33_24;
    _zz_io_MatrixB_33_26 <= _zz_io_MatrixB_33_25;
    _zz_io_MatrixB_33_27 <= _zz_io_MatrixB_33_26;
    _zz_io_MatrixB_33_28 <= _zz_io_MatrixB_33_27;
    _zz_io_MatrixB_33_29 <= _zz_io_MatrixB_33_28;
    _zz_io_MatrixB_33_30 <= _zz_io_MatrixB_33_29;
    _zz_io_MatrixB_33_31 <= _zz_io_MatrixB_33_30;
    _zz_io_MatrixB_33_32 <= _zz_io_MatrixB_33_31;
    _zz_io_B_Valid_33 <= SubModule_WeightCache_MatrixCol_Switch[33];
    _zz_io_B_Valid_33_1 <= _zz_io_B_Valid_33;
    _zz_io_B_Valid_33_2 <= _zz_io_B_Valid_33_1;
    _zz_io_B_Valid_33_3 <= _zz_io_B_Valid_33_2;
    _zz_io_B_Valid_33_4 <= _zz_io_B_Valid_33_3;
    _zz_io_B_Valid_33_5 <= _zz_io_B_Valid_33_4;
    _zz_io_B_Valid_33_6 <= _zz_io_B_Valid_33_5;
    _zz_io_B_Valid_33_7 <= _zz_io_B_Valid_33_6;
    _zz_io_B_Valid_33_8 <= _zz_io_B_Valid_33_7;
    _zz_io_B_Valid_33_9 <= _zz_io_B_Valid_33_8;
    _zz_io_B_Valid_33_10 <= _zz_io_B_Valid_33_9;
    _zz_io_B_Valid_33_11 <= _zz_io_B_Valid_33_10;
    _zz_io_B_Valid_33_12 <= _zz_io_B_Valid_33_11;
    _zz_io_B_Valid_33_13 <= _zz_io_B_Valid_33_12;
    _zz_io_B_Valid_33_14 <= _zz_io_B_Valid_33_13;
    _zz_io_B_Valid_33_15 <= _zz_io_B_Valid_33_14;
    _zz_io_B_Valid_33_16 <= _zz_io_B_Valid_33_15;
    _zz_io_B_Valid_33_17 <= _zz_io_B_Valid_33_16;
    _zz_io_B_Valid_33_18 <= _zz_io_B_Valid_33_17;
    _zz_io_B_Valid_33_19 <= _zz_io_B_Valid_33_18;
    _zz_io_B_Valid_33_20 <= _zz_io_B_Valid_33_19;
    _zz_io_B_Valid_33_21 <= _zz_io_B_Valid_33_20;
    _zz_io_B_Valid_33_22 <= _zz_io_B_Valid_33_21;
    _zz_io_B_Valid_33_23 <= _zz_io_B_Valid_33_22;
    _zz_io_B_Valid_33_24 <= _zz_io_B_Valid_33_23;
    _zz_io_B_Valid_33_25 <= _zz_io_B_Valid_33_24;
    _zz_io_B_Valid_33_26 <= _zz_io_B_Valid_33_25;
    _zz_io_B_Valid_33_27 <= _zz_io_B_Valid_33_26;
    _zz_io_B_Valid_33_28 <= _zz_io_B_Valid_33_27;
    _zz_io_B_Valid_33_29 <= _zz_io_B_Valid_33_28;
    _zz_io_B_Valid_33_30 <= _zz_io_B_Valid_33_29;
    _zz_io_B_Valid_33_31 <= _zz_io_B_Valid_33_30;
    _zz_io_B_Valid_33_32 <= _zz_io_B_Valid_33_31;
    _zz_io_MatrixB_34 <= SubModule_WeightCache_mData_34;
    _zz_io_MatrixB_34_1 <= _zz_io_MatrixB_34;
    _zz_io_MatrixB_34_2 <= _zz_io_MatrixB_34_1;
    _zz_io_MatrixB_34_3 <= _zz_io_MatrixB_34_2;
    _zz_io_MatrixB_34_4 <= _zz_io_MatrixB_34_3;
    _zz_io_MatrixB_34_5 <= _zz_io_MatrixB_34_4;
    _zz_io_MatrixB_34_6 <= _zz_io_MatrixB_34_5;
    _zz_io_MatrixB_34_7 <= _zz_io_MatrixB_34_6;
    _zz_io_MatrixB_34_8 <= _zz_io_MatrixB_34_7;
    _zz_io_MatrixB_34_9 <= _zz_io_MatrixB_34_8;
    _zz_io_MatrixB_34_10 <= _zz_io_MatrixB_34_9;
    _zz_io_MatrixB_34_11 <= _zz_io_MatrixB_34_10;
    _zz_io_MatrixB_34_12 <= _zz_io_MatrixB_34_11;
    _zz_io_MatrixB_34_13 <= _zz_io_MatrixB_34_12;
    _zz_io_MatrixB_34_14 <= _zz_io_MatrixB_34_13;
    _zz_io_MatrixB_34_15 <= _zz_io_MatrixB_34_14;
    _zz_io_MatrixB_34_16 <= _zz_io_MatrixB_34_15;
    _zz_io_MatrixB_34_17 <= _zz_io_MatrixB_34_16;
    _zz_io_MatrixB_34_18 <= _zz_io_MatrixB_34_17;
    _zz_io_MatrixB_34_19 <= _zz_io_MatrixB_34_18;
    _zz_io_MatrixB_34_20 <= _zz_io_MatrixB_34_19;
    _zz_io_MatrixB_34_21 <= _zz_io_MatrixB_34_20;
    _zz_io_MatrixB_34_22 <= _zz_io_MatrixB_34_21;
    _zz_io_MatrixB_34_23 <= _zz_io_MatrixB_34_22;
    _zz_io_MatrixB_34_24 <= _zz_io_MatrixB_34_23;
    _zz_io_MatrixB_34_25 <= _zz_io_MatrixB_34_24;
    _zz_io_MatrixB_34_26 <= _zz_io_MatrixB_34_25;
    _zz_io_MatrixB_34_27 <= _zz_io_MatrixB_34_26;
    _zz_io_MatrixB_34_28 <= _zz_io_MatrixB_34_27;
    _zz_io_MatrixB_34_29 <= _zz_io_MatrixB_34_28;
    _zz_io_MatrixB_34_30 <= _zz_io_MatrixB_34_29;
    _zz_io_MatrixB_34_31 <= _zz_io_MatrixB_34_30;
    _zz_io_MatrixB_34_32 <= _zz_io_MatrixB_34_31;
    _zz_io_MatrixB_34_33 <= _zz_io_MatrixB_34_32;
    _zz_io_B_Valid_34 <= SubModule_WeightCache_MatrixCol_Switch[34];
    _zz_io_B_Valid_34_1 <= _zz_io_B_Valid_34;
    _zz_io_B_Valid_34_2 <= _zz_io_B_Valid_34_1;
    _zz_io_B_Valid_34_3 <= _zz_io_B_Valid_34_2;
    _zz_io_B_Valid_34_4 <= _zz_io_B_Valid_34_3;
    _zz_io_B_Valid_34_5 <= _zz_io_B_Valid_34_4;
    _zz_io_B_Valid_34_6 <= _zz_io_B_Valid_34_5;
    _zz_io_B_Valid_34_7 <= _zz_io_B_Valid_34_6;
    _zz_io_B_Valid_34_8 <= _zz_io_B_Valid_34_7;
    _zz_io_B_Valid_34_9 <= _zz_io_B_Valid_34_8;
    _zz_io_B_Valid_34_10 <= _zz_io_B_Valid_34_9;
    _zz_io_B_Valid_34_11 <= _zz_io_B_Valid_34_10;
    _zz_io_B_Valid_34_12 <= _zz_io_B_Valid_34_11;
    _zz_io_B_Valid_34_13 <= _zz_io_B_Valid_34_12;
    _zz_io_B_Valid_34_14 <= _zz_io_B_Valid_34_13;
    _zz_io_B_Valid_34_15 <= _zz_io_B_Valid_34_14;
    _zz_io_B_Valid_34_16 <= _zz_io_B_Valid_34_15;
    _zz_io_B_Valid_34_17 <= _zz_io_B_Valid_34_16;
    _zz_io_B_Valid_34_18 <= _zz_io_B_Valid_34_17;
    _zz_io_B_Valid_34_19 <= _zz_io_B_Valid_34_18;
    _zz_io_B_Valid_34_20 <= _zz_io_B_Valid_34_19;
    _zz_io_B_Valid_34_21 <= _zz_io_B_Valid_34_20;
    _zz_io_B_Valid_34_22 <= _zz_io_B_Valid_34_21;
    _zz_io_B_Valid_34_23 <= _zz_io_B_Valid_34_22;
    _zz_io_B_Valid_34_24 <= _zz_io_B_Valid_34_23;
    _zz_io_B_Valid_34_25 <= _zz_io_B_Valid_34_24;
    _zz_io_B_Valid_34_26 <= _zz_io_B_Valid_34_25;
    _zz_io_B_Valid_34_27 <= _zz_io_B_Valid_34_26;
    _zz_io_B_Valid_34_28 <= _zz_io_B_Valid_34_27;
    _zz_io_B_Valid_34_29 <= _zz_io_B_Valid_34_28;
    _zz_io_B_Valid_34_30 <= _zz_io_B_Valid_34_29;
    _zz_io_B_Valid_34_31 <= _zz_io_B_Valid_34_30;
    _zz_io_B_Valid_34_32 <= _zz_io_B_Valid_34_31;
    _zz_io_B_Valid_34_33 <= _zz_io_B_Valid_34_32;
    _zz_io_MatrixB_35 <= SubModule_WeightCache_mData_35;
    _zz_io_MatrixB_35_1 <= _zz_io_MatrixB_35;
    _zz_io_MatrixB_35_2 <= _zz_io_MatrixB_35_1;
    _zz_io_MatrixB_35_3 <= _zz_io_MatrixB_35_2;
    _zz_io_MatrixB_35_4 <= _zz_io_MatrixB_35_3;
    _zz_io_MatrixB_35_5 <= _zz_io_MatrixB_35_4;
    _zz_io_MatrixB_35_6 <= _zz_io_MatrixB_35_5;
    _zz_io_MatrixB_35_7 <= _zz_io_MatrixB_35_6;
    _zz_io_MatrixB_35_8 <= _zz_io_MatrixB_35_7;
    _zz_io_MatrixB_35_9 <= _zz_io_MatrixB_35_8;
    _zz_io_MatrixB_35_10 <= _zz_io_MatrixB_35_9;
    _zz_io_MatrixB_35_11 <= _zz_io_MatrixB_35_10;
    _zz_io_MatrixB_35_12 <= _zz_io_MatrixB_35_11;
    _zz_io_MatrixB_35_13 <= _zz_io_MatrixB_35_12;
    _zz_io_MatrixB_35_14 <= _zz_io_MatrixB_35_13;
    _zz_io_MatrixB_35_15 <= _zz_io_MatrixB_35_14;
    _zz_io_MatrixB_35_16 <= _zz_io_MatrixB_35_15;
    _zz_io_MatrixB_35_17 <= _zz_io_MatrixB_35_16;
    _zz_io_MatrixB_35_18 <= _zz_io_MatrixB_35_17;
    _zz_io_MatrixB_35_19 <= _zz_io_MatrixB_35_18;
    _zz_io_MatrixB_35_20 <= _zz_io_MatrixB_35_19;
    _zz_io_MatrixB_35_21 <= _zz_io_MatrixB_35_20;
    _zz_io_MatrixB_35_22 <= _zz_io_MatrixB_35_21;
    _zz_io_MatrixB_35_23 <= _zz_io_MatrixB_35_22;
    _zz_io_MatrixB_35_24 <= _zz_io_MatrixB_35_23;
    _zz_io_MatrixB_35_25 <= _zz_io_MatrixB_35_24;
    _zz_io_MatrixB_35_26 <= _zz_io_MatrixB_35_25;
    _zz_io_MatrixB_35_27 <= _zz_io_MatrixB_35_26;
    _zz_io_MatrixB_35_28 <= _zz_io_MatrixB_35_27;
    _zz_io_MatrixB_35_29 <= _zz_io_MatrixB_35_28;
    _zz_io_MatrixB_35_30 <= _zz_io_MatrixB_35_29;
    _zz_io_MatrixB_35_31 <= _zz_io_MatrixB_35_30;
    _zz_io_MatrixB_35_32 <= _zz_io_MatrixB_35_31;
    _zz_io_MatrixB_35_33 <= _zz_io_MatrixB_35_32;
    _zz_io_MatrixB_35_34 <= _zz_io_MatrixB_35_33;
    _zz_io_B_Valid_35 <= SubModule_WeightCache_MatrixCol_Switch[35];
    _zz_io_B_Valid_35_1 <= _zz_io_B_Valid_35;
    _zz_io_B_Valid_35_2 <= _zz_io_B_Valid_35_1;
    _zz_io_B_Valid_35_3 <= _zz_io_B_Valid_35_2;
    _zz_io_B_Valid_35_4 <= _zz_io_B_Valid_35_3;
    _zz_io_B_Valid_35_5 <= _zz_io_B_Valid_35_4;
    _zz_io_B_Valid_35_6 <= _zz_io_B_Valid_35_5;
    _zz_io_B_Valid_35_7 <= _zz_io_B_Valid_35_6;
    _zz_io_B_Valid_35_8 <= _zz_io_B_Valid_35_7;
    _zz_io_B_Valid_35_9 <= _zz_io_B_Valid_35_8;
    _zz_io_B_Valid_35_10 <= _zz_io_B_Valid_35_9;
    _zz_io_B_Valid_35_11 <= _zz_io_B_Valid_35_10;
    _zz_io_B_Valid_35_12 <= _zz_io_B_Valid_35_11;
    _zz_io_B_Valid_35_13 <= _zz_io_B_Valid_35_12;
    _zz_io_B_Valid_35_14 <= _zz_io_B_Valid_35_13;
    _zz_io_B_Valid_35_15 <= _zz_io_B_Valid_35_14;
    _zz_io_B_Valid_35_16 <= _zz_io_B_Valid_35_15;
    _zz_io_B_Valid_35_17 <= _zz_io_B_Valid_35_16;
    _zz_io_B_Valid_35_18 <= _zz_io_B_Valid_35_17;
    _zz_io_B_Valid_35_19 <= _zz_io_B_Valid_35_18;
    _zz_io_B_Valid_35_20 <= _zz_io_B_Valid_35_19;
    _zz_io_B_Valid_35_21 <= _zz_io_B_Valid_35_20;
    _zz_io_B_Valid_35_22 <= _zz_io_B_Valid_35_21;
    _zz_io_B_Valid_35_23 <= _zz_io_B_Valid_35_22;
    _zz_io_B_Valid_35_24 <= _zz_io_B_Valid_35_23;
    _zz_io_B_Valid_35_25 <= _zz_io_B_Valid_35_24;
    _zz_io_B_Valid_35_26 <= _zz_io_B_Valid_35_25;
    _zz_io_B_Valid_35_27 <= _zz_io_B_Valid_35_26;
    _zz_io_B_Valid_35_28 <= _zz_io_B_Valid_35_27;
    _zz_io_B_Valid_35_29 <= _zz_io_B_Valid_35_28;
    _zz_io_B_Valid_35_30 <= _zz_io_B_Valid_35_29;
    _zz_io_B_Valid_35_31 <= _zz_io_B_Valid_35_30;
    _zz_io_B_Valid_35_32 <= _zz_io_B_Valid_35_31;
    _zz_io_B_Valid_35_33 <= _zz_io_B_Valid_35_32;
    _zz_io_B_Valid_35_34 <= _zz_io_B_Valid_35_33;
    _zz_io_MatrixB_36 <= SubModule_WeightCache_mData_36;
    _zz_io_MatrixB_36_1 <= _zz_io_MatrixB_36;
    _zz_io_MatrixB_36_2 <= _zz_io_MatrixB_36_1;
    _zz_io_MatrixB_36_3 <= _zz_io_MatrixB_36_2;
    _zz_io_MatrixB_36_4 <= _zz_io_MatrixB_36_3;
    _zz_io_MatrixB_36_5 <= _zz_io_MatrixB_36_4;
    _zz_io_MatrixB_36_6 <= _zz_io_MatrixB_36_5;
    _zz_io_MatrixB_36_7 <= _zz_io_MatrixB_36_6;
    _zz_io_MatrixB_36_8 <= _zz_io_MatrixB_36_7;
    _zz_io_MatrixB_36_9 <= _zz_io_MatrixB_36_8;
    _zz_io_MatrixB_36_10 <= _zz_io_MatrixB_36_9;
    _zz_io_MatrixB_36_11 <= _zz_io_MatrixB_36_10;
    _zz_io_MatrixB_36_12 <= _zz_io_MatrixB_36_11;
    _zz_io_MatrixB_36_13 <= _zz_io_MatrixB_36_12;
    _zz_io_MatrixB_36_14 <= _zz_io_MatrixB_36_13;
    _zz_io_MatrixB_36_15 <= _zz_io_MatrixB_36_14;
    _zz_io_MatrixB_36_16 <= _zz_io_MatrixB_36_15;
    _zz_io_MatrixB_36_17 <= _zz_io_MatrixB_36_16;
    _zz_io_MatrixB_36_18 <= _zz_io_MatrixB_36_17;
    _zz_io_MatrixB_36_19 <= _zz_io_MatrixB_36_18;
    _zz_io_MatrixB_36_20 <= _zz_io_MatrixB_36_19;
    _zz_io_MatrixB_36_21 <= _zz_io_MatrixB_36_20;
    _zz_io_MatrixB_36_22 <= _zz_io_MatrixB_36_21;
    _zz_io_MatrixB_36_23 <= _zz_io_MatrixB_36_22;
    _zz_io_MatrixB_36_24 <= _zz_io_MatrixB_36_23;
    _zz_io_MatrixB_36_25 <= _zz_io_MatrixB_36_24;
    _zz_io_MatrixB_36_26 <= _zz_io_MatrixB_36_25;
    _zz_io_MatrixB_36_27 <= _zz_io_MatrixB_36_26;
    _zz_io_MatrixB_36_28 <= _zz_io_MatrixB_36_27;
    _zz_io_MatrixB_36_29 <= _zz_io_MatrixB_36_28;
    _zz_io_MatrixB_36_30 <= _zz_io_MatrixB_36_29;
    _zz_io_MatrixB_36_31 <= _zz_io_MatrixB_36_30;
    _zz_io_MatrixB_36_32 <= _zz_io_MatrixB_36_31;
    _zz_io_MatrixB_36_33 <= _zz_io_MatrixB_36_32;
    _zz_io_MatrixB_36_34 <= _zz_io_MatrixB_36_33;
    _zz_io_MatrixB_36_35 <= _zz_io_MatrixB_36_34;
    _zz_io_B_Valid_36 <= SubModule_WeightCache_MatrixCol_Switch[36];
    _zz_io_B_Valid_36_1 <= _zz_io_B_Valid_36;
    _zz_io_B_Valid_36_2 <= _zz_io_B_Valid_36_1;
    _zz_io_B_Valid_36_3 <= _zz_io_B_Valid_36_2;
    _zz_io_B_Valid_36_4 <= _zz_io_B_Valid_36_3;
    _zz_io_B_Valid_36_5 <= _zz_io_B_Valid_36_4;
    _zz_io_B_Valid_36_6 <= _zz_io_B_Valid_36_5;
    _zz_io_B_Valid_36_7 <= _zz_io_B_Valid_36_6;
    _zz_io_B_Valid_36_8 <= _zz_io_B_Valid_36_7;
    _zz_io_B_Valid_36_9 <= _zz_io_B_Valid_36_8;
    _zz_io_B_Valid_36_10 <= _zz_io_B_Valid_36_9;
    _zz_io_B_Valid_36_11 <= _zz_io_B_Valid_36_10;
    _zz_io_B_Valid_36_12 <= _zz_io_B_Valid_36_11;
    _zz_io_B_Valid_36_13 <= _zz_io_B_Valid_36_12;
    _zz_io_B_Valid_36_14 <= _zz_io_B_Valid_36_13;
    _zz_io_B_Valid_36_15 <= _zz_io_B_Valid_36_14;
    _zz_io_B_Valid_36_16 <= _zz_io_B_Valid_36_15;
    _zz_io_B_Valid_36_17 <= _zz_io_B_Valid_36_16;
    _zz_io_B_Valid_36_18 <= _zz_io_B_Valid_36_17;
    _zz_io_B_Valid_36_19 <= _zz_io_B_Valid_36_18;
    _zz_io_B_Valid_36_20 <= _zz_io_B_Valid_36_19;
    _zz_io_B_Valid_36_21 <= _zz_io_B_Valid_36_20;
    _zz_io_B_Valid_36_22 <= _zz_io_B_Valid_36_21;
    _zz_io_B_Valid_36_23 <= _zz_io_B_Valid_36_22;
    _zz_io_B_Valid_36_24 <= _zz_io_B_Valid_36_23;
    _zz_io_B_Valid_36_25 <= _zz_io_B_Valid_36_24;
    _zz_io_B_Valid_36_26 <= _zz_io_B_Valid_36_25;
    _zz_io_B_Valid_36_27 <= _zz_io_B_Valid_36_26;
    _zz_io_B_Valid_36_28 <= _zz_io_B_Valid_36_27;
    _zz_io_B_Valid_36_29 <= _zz_io_B_Valid_36_28;
    _zz_io_B_Valid_36_30 <= _zz_io_B_Valid_36_29;
    _zz_io_B_Valid_36_31 <= _zz_io_B_Valid_36_30;
    _zz_io_B_Valid_36_32 <= _zz_io_B_Valid_36_31;
    _zz_io_B_Valid_36_33 <= _zz_io_B_Valid_36_32;
    _zz_io_B_Valid_36_34 <= _zz_io_B_Valid_36_33;
    _zz_io_B_Valid_36_35 <= _zz_io_B_Valid_36_34;
    _zz_io_MatrixB_37 <= SubModule_WeightCache_mData_37;
    _zz_io_MatrixB_37_1 <= _zz_io_MatrixB_37;
    _zz_io_MatrixB_37_2 <= _zz_io_MatrixB_37_1;
    _zz_io_MatrixB_37_3 <= _zz_io_MatrixB_37_2;
    _zz_io_MatrixB_37_4 <= _zz_io_MatrixB_37_3;
    _zz_io_MatrixB_37_5 <= _zz_io_MatrixB_37_4;
    _zz_io_MatrixB_37_6 <= _zz_io_MatrixB_37_5;
    _zz_io_MatrixB_37_7 <= _zz_io_MatrixB_37_6;
    _zz_io_MatrixB_37_8 <= _zz_io_MatrixB_37_7;
    _zz_io_MatrixB_37_9 <= _zz_io_MatrixB_37_8;
    _zz_io_MatrixB_37_10 <= _zz_io_MatrixB_37_9;
    _zz_io_MatrixB_37_11 <= _zz_io_MatrixB_37_10;
    _zz_io_MatrixB_37_12 <= _zz_io_MatrixB_37_11;
    _zz_io_MatrixB_37_13 <= _zz_io_MatrixB_37_12;
    _zz_io_MatrixB_37_14 <= _zz_io_MatrixB_37_13;
    _zz_io_MatrixB_37_15 <= _zz_io_MatrixB_37_14;
    _zz_io_MatrixB_37_16 <= _zz_io_MatrixB_37_15;
    _zz_io_MatrixB_37_17 <= _zz_io_MatrixB_37_16;
    _zz_io_MatrixB_37_18 <= _zz_io_MatrixB_37_17;
    _zz_io_MatrixB_37_19 <= _zz_io_MatrixB_37_18;
    _zz_io_MatrixB_37_20 <= _zz_io_MatrixB_37_19;
    _zz_io_MatrixB_37_21 <= _zz_io_MatrixB_37_20;
    _zz_io_MatrixB_37_22 <= _zz_io_MatrixB_37_21;
    _zz_io_MatrixB_37_23 <= _zz_io_MatrixB_37_22;
    _zz_io_MatrixB_37_24 <= _zz_io_MatrixB_37_23;
    _zz_io_MatrixB_37_25 <= _zz_io_MatrixB_37_24;
    _zz_io_MatrixB_37_26 <= _zz_io_MatrixB_37_25;
    _zz_io_MatrixB_37_27 <= _zz_io_MatrixB_37_26;
    _zz_io_MatrixB_37_28 <= _zz_io_MatrixB_37_27;
    _zz_io_MatrixB_37_29 <= _zz_io_MatrixB_37_28;
    _zz_io_MatrixB_37_30 <= _zz_io_MatrixB_37_29;
    _zz_io_MatrixB_37_31 <= _zz_io_MatrixB_37_30;
    _zz_io_MatrixB_37_32 <= _zz_io_MatrixB_37_31;
    _zz_io_MatrixB_37_33 <= _zz_io_MatrixB_37_32;
    _zz_io_MatrixB_37_34 <= _zz_io_MatrixB_37_33;
    _zz_io_MatrixB_37_35 <= _zz_io_MatrixB_37_34;
    _zz_io_MatrixB_37_36 <= _zz_io_MatrixB_37_35;
    _zz_io_B_Valid_37 <= SubModule_WeightCache_MatrixCol_Switch[37];
    _zz_io_B_Valid_37_1 <= _zz_io_B_Valid_37;
    _zz_io_B_Valid_37_2 <= _zz_io_B_Valid_37_1;
    _zz_io_B_Valid_37_3 <= _zz_io_B_Valid_37_2;
    _zz_io_B_Valid_37_4 <= _zz_io_B_Valid_37_3;
    _zz_io_B_Valid_37_5 <= _zz_io_B_Valid_37_4;
    _zz_io_B_Valid_37_6 <= _zz_io_B_Valid_37_5;
    _zz_io_B_Valid_37_7 <= _zz_io_B_Valid_37_6;
    _zz_io_B_Valid_37_8 <= _zz_io_B_Valid_37_7;
    _zz_io_B_Valid_37_9 <= _zz_io_B_Valid_37_8;
    _zz_io_B_Valid_37_10 <= _zz_io_B_Valid_37_9;
    _zz_io_B_Valid_37_11 <= _zz_io_B_Valid_37_10;
    _zz_io_B_Valid_37_12 <= _zz_io_B_Valid_37_11;
    _zz_io_B_Valid_37_13 <= _zz_io_B_Valid_37_12;
    _zz_io_B_Valid_37_14 <= _zz_io_B_Valid_37_13;
    _zz_io_B_Valid_37_15 <= _zz_io_B_Valid_37_14;
    _zz_io_B_Valid_37_16 <= _zz_io_B_Valid_37_15;
    _zz_io_B_Valid_37_17 <= _zz_io_B_Valid_37_16;
    _zz_io_B_Valid_37_18 <= _zz_io_B_Valid_37_17;
    _zz_io_B_Valid_37_19 <= _zz_io_B_Valid_37_18;
    _zz_io_B_Valid_37_20 <= _zz_io_B_Valid_37_19;
    _zz_io_B_Valid_37_21 <= _zz_io_B_Valid_37_20;
    _zz_io_B_Valid_37_22 <= _zz_io_B_Valid_37_21;
    _zz_io_B_Valid_37_23 <= _zz_io_B_Valid_37_22;
    _zz_io_B_Valid_37_24 <= _zz_io_B_Valid_37_23;
    _zz_io_B_Valid_37_25 <= _zz_io_B_Valid_37_24;
    _zz_io_B_Valid_37_26 <= _zz_io_B_Valid_37_25;
    _zz_io_B_Valid_37_27 <= _zz_io_B_Valid_37_26;
    _zz_io_B_Valid_37_28 <= _zz_io_B_Valid_37_27;
    _zz_io_B_Valid_37_29 <= _zz_io_B_Valid_37_28;
    _zz_io_B_Valid_37_30 <= _zz_io_B_Valid_37_29;
    _zz_io_B_Valid_37_31 <= _zz_io_B_Valid_37_30;
    _zz_io_B_Valid_37_32 <= _zz_io_B_Valid_37_31;
    _zz_io_B_Valid_37_33 <= _zz_io_B_Valid_37_32;
    _zz_io_B_Valid_37_34 <= _zz_io_B_Valid_37_33;
    _zz_io_B_Valid_37_35 <= _zz_io_B_Valid_37_34;
    _zz_io_B_Valid_37_36 <= _zz_io_B_Valid_37_35;
    _zz_io_MatrixB_38 <= SubModule_WeightCache_mData_38;
    _zz_io_MatrixB_38_1 <= _zz_io_MatrixB_38;
    _zz_io_MatrixB_38_2 <= _zz_io_MatrixB_38_1;
    _zz_io_MatrixB_38_3 <= _zz_io_MatrixB_38_2;
    _zz_io_MatrixB_38_4 <= _zz_io_MatrixB_38_3;
    _zz_io_MatrixB_38_5 <= _zz_io_MatrixB_38_4;
    _zz_io_MatrixB_38_6 <= _zz_io_MatrixB_38_5;
    _zz_io_MatrixB_38_7 <= _zz_io_MatrixB_38_6;
    _zz_io_MatrixB_38_8 <= _zz_io_MatrixB_38_7;
    _zz_io_MatrixB_38_9 <= _zz_io_MatrixB_38_8;
    _zz_io_MatrixB_38_10 <= _zz_io_MatrixB_38_9;
    _zz_io_MatrixB_38_11 <= _zz_io_MatrixB_38_10;
    _zz_io_MatrixB_38_12 <= _zz_io_MatrixB_38_11;
    _zz_io_MatrixB_38_13 <= _zz_io_MatrixB_38_12;
    _zz_io_MatrixB_38_14 <= _zz_io_MatrixB_38_13;
    _zz_io_MatrixB_38_15 <= _zz_io_MatrixB_38_14;
    _zz_io_MatrixB_38_16 <= _zz_io_MatrixB_38_15;
    _zz_io_MatrixB_38_17 <= _zz_io_MatrixB_38_16;
    _zz_io_MatrixB_38_18 <= _zz_io_MatrixB_38_17;
    _zz_io_MatrixB_38_19 <= _zz_io_MatrixB_38_18;
    _zz_io_MatrixB_38_20 <= _zz_io_MatrixB_38_19;
    _zz_io_MatrixB_38_21 <= _zz_io_MatrixB_38_20;
    _zz_io_MatrixB_38_22 <= _zz_io_MatrixB_38_21;
    _zz_io_MatrixB_38_23 <= _zz_io_MatrixB_38_22;
    _zz_io_MatrixB_38_24 <= _zz_io_MatrixB_38_23;
    _zz_io_MatrixB_38_25 <= _zz_io_MatrixB_38_24;
    _zz_io_MatrixB_38_26 <= _zz_io_MatrixB_38_25;
    _zz_io_MatrixB_38_27 <= _zz_io_MatrixB_38_26;
    _zz_io_MatrixB_38_28 <= _zz_io_MatrixB_38_27;
    _zz_io_MatrixB_38_29 <= _zz_io_MatrixB_38_28;
    _zz_io_MatrixB_38_30 <= _zz_io_MatrixB_38_29;
    _zz_io_MatrixB_38_31 <= _zz_io_MatrixB_38_30;
    _zz_io_MatrixB_38_32 <= _zz_io_MatrixB_38_31;
    _zz_io_MatrixB_38_33 <= _zz_io_MatrixB_38_32;
    _zz_io_MatrixB_38_34 <= _zz_io_MatrixB_38_33;
    _zz_io_MatrixB_38_35 <= _zz_io_MatrixB_38_34;
    _zz_io_MatrixB_38_36 <= _zz_io_MatrixB_38_35;
    _zz_io_MatrixB_38_37 <= _zz_io_MatrixB_38_36;
    _zz_io_B_Valid_38 <= SubModule_WeightCache_MatrixCol_Switch[38];
    _zz_io_B_Valid_38_1 <= _zz_io_B_Valid_38;
    _zz_io_B_Valid_38_2 <= _zz_io_B_Valid_38_1;
    _zz_io_B_Valid_38_3 <= _zz_io_B_Valid_38_2;
    _zz_io_B_Valid_38_4 <= _zz_io_B_Valid_38_3;
    _zz_io_B_Valid_38_5 <= _zz_io_B_Valid_38_4;
    _zz_io_B_Valid_38_6 <= _zz_io_B_Valid_38_5;
    _zz_io_B_Valid_38_7 <= _zz_io_B_Valid_38_6;
    _zz_io_B_Valid_38_8 <= _zz_io_B_Valid_38_7;
    _zz_io_B_Valid_38_9 <= _zz_io_B_Valid_38_8;
    _zz_io_B_Valid_38_10 <= _zz_io_B_Valid_38_9;
    _zz_io_B_Valid_38_11 <= _zz_io_B_Valid_38_10;
    _zz_io_B_Valid_38_12 <= _zz_io_B_Valid_38_11;
    _zz_io_B_Valid_38_13 <= _zz_io_B_Valid_38_12;
    _zz_io_B_Valid_38_14 <= _zz_io_B_Valid_38_13;
    _zz_io_B_Valid_38_15 <= _zz_io_B_Valid_38_14;
    _zz_io_B_Valid_38_16 <= _zz_io_B_Valid_38_15;
    _zz_io_B_Valid_38_17 <= _zz_io_B_Valid_38_16;
    _zz_io_B_Valid_38_18 <= _zz_io_B_Valid_38_17;
    _zz_io_B_Valid_38_19 <= _zz_io_B_Valid_38_18;
    _zz_io_B_Valid_38_20 <= _zz_io_B_Valid_38_19;
    _zz_io_B_Valid_38_21 <= _zz_io_B_Valid_38_20;
    _zz_io_B_Valid_38_22 <= _zz_io_B_Valid_38_21;
    _zz_io_B_Valid_38_23 <= _zz_io_B_Valid_38_22;
    _zz_io_B_Valid_38_24 <= _zz_io_B_Valid_38_23;
    _zz_io_B_Valid_38_25 <= _zz_io_B_Valid_38_24;
    _zz_io_B_Valid_38_26 <= _zz_io_B_Valid_38_25;
    _zz_io_B_Valid_38_27 <= _zz_io_B_Valid_38_26;
    _zz_io_B_Valid_38_28 <= _zz_io_B_Valid_38_27;
    _zz_io_B_Valid_38_29 <= _zz_io_B_Valid_38_28;
    _zz_io_B_Valid_38_30 <= _zz_io_B_Valid_38_29;
    _zz_io_B_Valid_38_31 <= _zz_io_B_Valid_38_30;
    _zz_io_B_Valid_38_32 <= _zz_io_B_Valid_38_31;
    _zz_io_B_Valid_38_33 <= _zz_io_B_Valid_38_32;
    _zz_io_B_Valid_38_34 <= _zz_io_B_Valid_38_33;
    _zz_io_B_Valid_38_35 <= _zz_io_B_Valid_38_34;
    _zz_io_B_Valid_38_36 <= _zz_io_B_Valid_38_35;
    _zz_io_B_Valid_38_37 <= _zz_io_B_Valid_38_36;
    _zz_io_MatrixB_39 <= SubModule_WeightCache_mData_39;
    _zz_io_MatrixB_39_1 <= _zz_io_MatrixB_39;
    _zz_io_MatrixB_39_2 <= _zz_io_MatrixB_39_1;
    _zz_io_MatrixB_39_3 <= _zz_io_MatrixB_39_2;
    _zz_io_MatrixB_39_4 <= _zz_io_MatrixB_39_3;
    _zz_io_MatrixB_39_5 <= _zz_io_MatrixB_39_4;
    _zz_io_MatrixB_39_6 <= _zz_io_MatrixB_39_5;
    _zz_io_MatrixB_39_7 <= _zz_io_MatrixB_39_6;
    _zz_io_MatrixB_39_8 <= _zz_io_MatrixB_39_7;
    _zz_io_MatrixB_39_9 <= _zz_io_MatrixB_39_8;
    _zz_io_MatrixB_39_10 <= _zz_io_MatrixB_39_9;
    _zz_io_MatrixB_39_11 <= _zz_io_MatrixB_39_10;
    _zz_io_MatrixB_39_12 <= _zz_io_MatrixB_39_11;
    _zz_io_MatrixB_39_13 <= _zz_io_MatrixB_39_12;
    _zz_io_MatrixB_39_14 <= _zz_io_MatrixB_39_13;
    _zz_io_MatrixB_39_15 <= _zz_io_MatrixB_39_14;
    _zz_io_MatrixB_39_16 <= _zz_io_MatrixB_39_15;
    _zz_io_MatrixB_39_17 <= _zz_io_MatrixB_39_16;
    _zz_io_MatrixB_39_18 <= _zz_io_MatrixB_39_17;
    _zz_io_MatrixB_39_19 <= _zz_io_MatrixB_39_18;
    _zz_io_MatrixB_39_20 <= _zz_io_MatrixB_39_19;
    _zz_io_MatrixB_39_21 <= _zz_io_MatrixB_39_20;
    _zz_io_MatrixB_39_22 <= _zz_io_MatrixB_39_21;
    _zz_io_MatrixB_39_23 <= _zz_io_MatrixB_39_22;
    _zz_io_MatrixB_39_24 <= _zz_io_MatrixB_39_23;
    _zz_io_MatrixB_39_25 <= _zz_io_MatrixB_39_24;
    _zz_io_MatrixB_39_26 <= _zz_io_MatrixB_39_25;
    _zz_io_MatrixB_39_27 <= _zz_io_MatrixB_39_26;
    _zz_io_MatrixB_39_28 <= _zz_io_MatrixB_39_27;
    _zz_io_MatrixB_39_29 <= _zz_io_MatrixB_39_28;
    _zz_io_MatrixB_39_30 <= _zz_io_MatrixB_39_29;
    _zz_io_MatrixB_39_31 <= _zz_io_MatrixB_39_30;
    _zz_io_MatrixB_39_32 <= _zz_io_MatrixB_39_31;
    _zz_io_MatrixB_39_33 <= _zz_io_MatrixB_39_32;
    _zz_io_MatrixB_39_34 <= _zz_io_MatrixB_39_33;
    _zz_io_MatrixB_39_35 <= _zz_io_MatrixB_39_34;
    _zz_io_MatrixB_39_36 <= _zz_io_MatrixB_39_35;
    _zz_io_MatrixB_39_37 <= _zz_io_MatrixB_39_36;
    _zz_io_MatrixB_39_38 <= _zz_io_MatrixB_39_37;
    _zz_io_B_Valid_39 <= SubModule_WeightCache_MatrixCol_Switch[39];
    _zz_io_B_Valid_39_1 <= _zz_io_B_Valid_39;
    _zz_io_B_Valid_39_2 <= _zz_io_B_Valid_39_1;
    _zz_io_B_Valid_39_3 <= _zz_io_B_Valid_39_2;
    _zz_io_B_Valid_39_4 <= _zz_io_B_Valid_39_3;
    _zz_io_B_Valid_39_5 <= _zz_io_B_Valid_39_4;
    _zz_io_B_Valid_39_6 <= _zz_io_B_Valid_39_5;
    _zz_io_B_Valid_39_7 <= _zz_io_B_Valid_39_6;
    _zz_io_B_Valid_39_8 <= _zz_io_B_Valid_39_7;
    _zz_io_B_Valid_39_9 <= _zz_io_B_Valid_39_8;
    _zz_io_B_Valid_39_10 <= _zz_io_B_Valid_39_9;
    _zz_io_B_Valid_39_11 <= _zz_io_B_Valid_39_10;
    _zz_io_B_Valid_39_12 <= _zz_io_B_Valid_39_11;
    _zz_io_B_Valid_39_13 <= _zz_io_B_Valid_39_12;
    _zz_io_B_Valid_39_14 <= _zz_io_B_Valid_39_13;
    _zz_io_B_Valid_39_15 <= _zz_io_B_Valid_39_14;
    _zz_io_B_Valid_39_16 <= _zz_io_B_Valid_39_15;
    _zz_io_B_Valid_39_17 <= _zz_io_B_Valid_39_16;
    _zz_io_B_Valid_39_18 <= _zz_io_B_Valid_39_17;
    _zz_io_B_Valid_39_19 <= _zz_io_B_Valid_39_18;
    _zz_io_B_Valid_39_20 <= _zz_io_B_Valid_39_19;
    _zz_io_B_Valid_39_21 <= _zz_io_B_Valid_39_20;
    _zz_io_B_Valid_39_22 <= _zz_io_B_Valid_39_21;
    _zz_io_B_Valid_39_23 <= _zz_io_B_Valid_39_22;
    _zz_io_B_Valid_39_24 <= _zz_io_B_Valid_39_23;
    _zz_io_B_Valid_39_25 <= _zz_io_B_Valid_39_24;
    _zz_io_B_Valid_39_26 <= _zz_io_B_Valid_39_25;
    _zz_io_B_Valid_39_27 <= _zz_io_B_Valid_39_26;
    _zz_io_B_Valid_39_28 <= _zz_io_B_Valid_39_27;
    _zz_io_B_Valid_39_29 <= _zz_io_B_Valid_39_28;
    _zz_io_B_Valid_39_30 <= _zz_io_B_Valid_39_29;
    _zz_io_B_Valid_39_31 <= _zz_io_B_Valid_39_30;
    _zz_io_B_Valid_39_32 <= _zz_io_B_Valid_39_31;
    _zz_io_B_Valid_39_33 <= _zz_io_B_Valid_39_32;
    _zz_io_B_Valid_39_34 <= _zz_io_B_Valid_39_33;
    _zz_io_B_Valid_39_35 <= _zz_io_B_Valid_39_34;
    _zz_io_B_Valid_39_36 <= _zz_io_B_Valid_39_35;
    _zz_io_B_Valid_39_37 <= _zz_io_B_Valid_39_36;
    _zz_io_B_Valid_39_38 <= _zz_io_B_Valid_39_37;
    _zz_io_MatrixB_40 <= SubModule_WeightCache_mData_40;
    _zz_io_MatrixB_40_1 <= _zz_io_MatrixB_40;
    _zz_io_MatrixB_40_2 <= _zz_io_MatrixB_40_1;
    _zz_io_MatrixB_40_3 <= _zz_io_MatrixB_40_2;
    _zz_io_MatrixB_40_4 <= _zz_io_MatrixB_40_3;
    _zz_io_MatrixB_40_5 <= _zz_io_MatrixB_40_4;
    _zz_io_MatrixB_40_6 <= _zz_io_MatrixB_40_5;
    _zz_io_MatrixB_40_7 <= _zz_io_MatrixB_40_6;
    _zz_io_MatrixB_40_8 <= _zz_io_MatrixB_40_7;
    _zz_io_MatrixB_40_9 <= _zz_io_MatrixB_40_8;
    _zz_io_MatrixB_40_10 <= _zz_io_MatrixB_40_9;
    _zz_io_MatrixB_40_11 <= _zz_io_MatrixB_40_10;
    _zz_io_MatrixB_40_12 <= _zz_io_MatrixB_40_11;
    _zz_io_MatrixB_40_13 <= _zz_io_MatrixB_40_12;
    _zz_io_MatrixB_40_14 <= _zz_io_MatrixB_40_13;
    _zz_io_MatrixB_40_15 <= _zz_io_MatrixB_40_14;
    _zz_io_MatrixB_40_16 <= _zz_io_MatrixB_40_15;
    _zz_io_MatrixB_40_17 <= _zz_io_MatrixB_40_16;
    _zz_io_MatrixB_40_18 <= _zz_io_MatrixB_40_17;
    _zz_io_MatrixB_40_19 <= _zz_io_MatrixB_40_18;
    _zz_io_MatrixB_40_20 <= _zz_io_MatrixB_40_19;
    _zz_io_MatrixB_40_21 <= _zz_io_MatrixB_40_20;
    _zz_io_MatrixB_40_22 <= _zz_io_MatrixB_40_21;
    _zz_io_MatrixB_40_23 <= _zz_io_MatrixB_40_22;
    _zz_io_MatrixB_40_24 <= _zz_io_MatrixB_40_23;
    _zz_io_MatrixB_40_25 <= _zz_io_MatrixB_40_24;
    _zz_io_MatrixB_40_26 <= _zz_io_MatrixB_40_25;
    _zz_io_MatrixB_40_27 <= _zz_io_MatrixB_40_26;
    _zz_io_MatrixB_40_28 <= _zz_io_MatrixB_40_27;
    _zz_io_MatrixB_40_29 <= _zz_io_MatrixB_40_28;
    _zz_io_MatrixB_40_30 <= _zz_io_MatrixB_40_29;
    _zz_io_MatrixB_40_31 <= _zz_io_MatrixB_40_30;
    _zz_io_MatrixB_40_32 <= _zz_io_MatrixB_40_31;
    _zz_io_MatrixB_40_33 <= _zz_io_MatrixB_40_32;
    _zz_io_MatrixB_40_34 <= _zz_io_MatrixB_40_33;
    _zz_io_MatrixB_40_35 <= _zz_io_MatrixB_40_34;
    _zz_io_MatrixB_40_36 <= _zz_io_MatrixB_40_35;
    _zz_io_MatrixB_40_37 <= _zz_io_MatrixB_40_36;
    _zz_io_MatrixB_40_38 <= _zz_io_MatrixB_40_37;
    _zz_io_MatrixB_40_39 <= _zz_io_MatrixB_40_38;
    _zz_io_B_Valid_40 <= SubModule_WeightCache_MatrixCol_Switch[40];
    _zz_io_B_Valid_40_1 <= _zz_io_B_Valid_40;
    _zz_io_B_Valid_40_2 <= _zz_io_B_Valid_40_1;
    _zz_io_B_Valid_40_3 <= _zz_io_B_Valid_40_2;
    _zz_io_B_Valid_40_4 <= _zz_io_B_Valid_40_3;
    _zz_io_B_Valid_40_5 <= _zz_io_B_Valid_40_4;
    _zz_io_B_Valid_40_6 <= _zz_io_B_Valid_40_5;
    _zz_io_B_Valid_40_7 <= _zz_io_B_Valid_40_6;
    _zz_io_B_Valid_40_8 <= _zz_io_B_Valid_40_7;
    _zz_io_B_Valid_40_9 <= _zz_io_B_Valid_40_8;
    _zz_io_B_Valid_40_10 <= _zz_io_B_Valid_40_9;
    _zz_io_B_Valid_40_11 <= _zz_io_B_Valid_40_10;
    _zz_io_B_Valid_40_12 <= _zz_io_B_Valid_40_11;
    _zz_io_B_Valid_40_13 <= _zz_io_B_Valid_40_12;
    _zz_io_B_Valid_40_14 <= _zz_io_B_Valid_40_13;
    _zz_io_B_Valid_40_15 <= _zz_io_B_Valid_40_14;
    _zz_io_B_Valid_40_16 <= _zz_io_B_Valid_40_15;
    _zz_io_B_Valid_40_17 <= _zz_io_B_Valid_40_16;
    _zz_io_B_Valid_40_18 <= _zz_io_B_Valid_40_17;
    _zz_io_B_Valid_40_19 <= _zz_io_B_Valid_40_18;
    _zz_io_B_Valid_40_20 <= _zz_io_B_Valid_40_19;
    _zz_io_B_Valid_40_21 <= _zz_io_B_Valid_40_20;
    _zz_io_B_Valid_40_22 <= _zz_io_B_Valid_40_21;
    _zz_io_B_Valid_40_23 <= _zz_io_B_Valid_40_22;
    _zz_io_B_Valid_40_24 <= _zz_io_B_Valid_40_23;
    _zz_io_B_Valid_40_25 <= _zz_io_B_Valid_40_24;
    _zz_io_B_Valid_40_26 <= _zz_io_B_Valid_40_25;
    _zz_io_B_Valid_40_27 <= _zz_io_B_Valid_40_26;
    _zz_io_B_Valid_40_28 <= _zz_io_B_Valid_40_27;
    _zz_io_B_Valid_40_29 <= _zz_io_B_Valid_40_28;
    _zz_io_B_Valid_40_30 <= _zz_io_B_Valid_40_29;
    _zz_io_B_Valid_40_31 <= _zz_io_B_Valid_40_30;
    _zz_io_B_Valid_40_32 <= _zz_io_B_Valid_40_31;
    _zz_io_B_Valid_40_33 <= _zz_io_B_Valid_40_32;
    _zz_io_B_Valid_40_34 <= _zz_io_B_Valid_40_33;
    _zz_io_B_Valid_40_35 <= _zz_io_B_Valid_40_34;
    _zz_io_B_Valid_40_36 <= _zz_io_B_Valid_40_35;
    _zz_io_B_Valid_40_37 <= _zz_io_B_Valid_40_36;
    _zz_io_B_Valid_40_38 <= _zz_io_B_Valid_40_37;
    _zz_io_B_Valid_40_39 <= _zz_io_B_Valid_40_38;
    _zz_io_MatrixB_41 <= SubModule_WeightCache_mData_41;
    _zz_io_MatrixB_41_1 <= _zz_io_MatrixB_41;
    _zz_io_MatrixB_41_2 <= _zz_io_MatrixB_41_1;
    _zz_io_MatrixB_41_3 <= _zz_io_MatrixB_41_2;
    _zz_io_MatrixB_41_4 <= _zz_io_MatrixB_41_3;
    _zz_io_MatrixB_41_5 <= _zz_io_MatrixB_41_4;
    _zz_io_MatrixB_41_6 <= _zz_io_MatrixB_41_5;
    _zz_io_MatrixB_41_7 <= _zz_io_MatrixB_41_6;
    _zz_io_MatrixB_41_8 <= _zz_io_MatrixB_41_7;
    _zz_io_MatrixB_41_9 <= _zz_io_MatrixB_41_8;
    _zz_io_MatrixB_41_10 <= _zz_io_MatrixB_41_9;
    _zz_io_MatrixB_41_11 <= _zz_io_MatrixB_41_10;
    _zz_io_MatrixB_41_12 <= _zz_io_MatrixB_41_11;
    _zz_io_MatrixB_41_13 <= _zz_io_MatrixB_41_12;
    _zz_io_MatrixB_41_14 <= _zz_io_MatrixB_41_13;
    _zz_io_MatrixB_41_15 <= _zz_io_MatrixB_41_14;
    _zz_io_MatrixB_41_16 <= _zz_io_MatrixB_41_15;
    _zz_io_MatrixB_41_17 <= _zz_io_MatrixB_41_16;
    _zz_io_MatrixB_41_18 <= _zz_io_MatrixB_41_17;
    _zz_io_MatrixB_41_19 <= _zz_io_MatrixB_41_18;
    _zz_io_MatrixB_41_20 <= _zz_io_MatrixB_41_19;
    _zz_io_MatrixB_41_21 <= _zz_io_MatrixB_41_20;
    _zz_io_MatrixB_41_22 <= _zz_io_MatrixB_41_21;
    _zz_io_MatrixB_41_23 <= _zz_io_MatrixB_41_22;
    _zz_io_MatrixB_41_24 <= _zz_io_MatrixB_41_23;
    _zz_io_MatrixB_41_25 <= _zz_io_MatrixB_41_24;
    _zz_io_MatrixB_41_26 <= _zz_io_MatrixB_41_25;
    _zz_io_MatrixB_41_27 <= _zz_io_MatrixB_41_26;
    _zz_io_MatrixB_41_28 <= _zz_io_MatrixB_41_27;
    _zz_io_MatrixB_41_29 <= _zz_io_MatrixB_41_28;
    _zz_io_MatrixB_41_30 <= _zz_io_MatrixB_41_29;
    _zz_io_MatrixB_41_31 <= _zz_io_MatrixB_41_30;
    _zz_io_MatrixB_41_32 <= _zz_io_MatrixB_41_31;
    _zz_io_MatrixB_41_33 <= _zz_io_MatrixB_41_32;
    _zz_io_MatrixB_41_34 <= _zz_io_MatrixB_41_33;
    _zz_io_MatrixB_41_35 <= _zz_io_MatrixB_41_34;
    _zz_io_MatrixB_41_36 <= _zz_io_MatrixB_41_35;
    _zz_io_MatrixB_41_37 <= _zz_io_MatrixB_41_36;
    _zz_io_MatrixB_41_38 <= _zz_io_MatrixB_41_37;
    _zz_io_MatrixB_41_39 <= _zz_io_MatrixB_41_38;
    _zz_io_MatrixB_41_40 <= _zz_io_MatrixB_41_39;
    _zz_io_B_Valid_41 <= SubModule_WeightCache_MatrixCol_Switch[41];
    _zz_io_B_Valid_41_1 <= _zz_io_B_Valid_41;
    _zz_io_B_Valid_41_2 <= _zz_io_B_Valid_41_1;
    _zz_io_B_Valid_41_3 <= _zz_io_B_Valid_41_2;
    _zz_io_B_Valid_41_4 <= _zz_io_B_Valid_41_3;
    _zz_io_B_Valid_41_5 <= _zz_io_B_Valid_41_4;
    _zz_io_B_Valid_41_6 <= _zz_io_B_Valid_41_5;
    _zz_io_B_Valid_41_7 <= _zz_io_B_Valid_41_6;
    _zz_io_B_Valid_41_8 <= _zz_io_B_Valid_41_7;
    _zz_io_B_Valid_41_9 <= _zz_io_B_Valid_41_8;
    _zz_io_B_Valid_41_10 <= _zz_io_B_Valid_41_9;
    _zz_io_B_Valid_41_11 <= _zz_io_B_Valid_41_10;
    _zz_io_B_Valid_41_12 <= _zz_io_B_Valid_41_11;
    _zz_io_B_Valid_41_13 <= _zz_io_B_Valid_41_12;
    _zz_io_B_Valid_41_14 <= _zz_io_B_Valid_41_13;
    _zz_io_B_Valid_41_15 <= _zz_io_B_Valid_41_14;
    _zz_io_B_Valid_41_16 <= _zz_io_B_Valid_41_15;
    _zz_io_B_Valid_41_17 <= _zz_io_B_Valid_41_16;
    _zz_io_B_Valid_41_18 <= _zz_io_B_Valid_41_17;
    _zz_io_B_Valid_41_19 <= _zz_io_B_Valid_41_18;
    _zz_io_B_Valid_41_20 <= _zz_io_B_Valid_41_19;
    _zz_io_B_Valid_41_21 <= _zz_io_B_Valid_41_20;
    _zz_io_B_Valid_41_22 <= _zz_io_B_Valid_41_21;
    _zz_io_B_Valid_41_23 <= _zz_io_B_Valid_41_22;
    _zz_io_B_Valid_41_24 <= _zz_io_B_Valid_41_23;
    _zz_io_B_Valid_41_25 <= _zz_io_B_Valid_41_24;
    _zz_io_B_Valid_41_26 <= _zz_io_B_Valid_41_25;
    _zz_io_B_Valid_41_27 <= _zz_io_B_Valid_41_26;
    _zz_io_B_Valid_41_28 <= _zz_io_B_Valid_41_27;
    _zz_io_B_Valid_41_29 <= _zz_io_B_Valid_41_28;
    _zz_io_B_Valid_41_30 <= _zz_io_B_Valid_41_29;
    _zz_io_B_Valid_41_31 <= _zz_io_B_Valid_41_30;
    _zz_io_B_Valid_41_32 <= _zz_io_B_Valid_41_31;
    _zz_io_B_Valid_41_33 <= _zz_io_B_Valid_41_32;
    _zz_io_B_Valid_41_34 <= _zz_io_B_Valid_41_33;
    _zz_io_B_Valid_41_35 <= _zz_io_B_Valid_41_34;
    _zz_io_B_Valid_41_36 <= _zz_io_B_Valid_41_35;
    _zz_io_B_Valid_41_37 <= _zz_io_B_Valid_41_36;
    _zz_io_B_Valid_41_38 <= _zz_io_B_Valid_41_37;
    _zz_io_B_Valid_41_39 <= _zz_io_B_Valid_41_38;
    _zz_io_B_Valid_41_40 <= _zz_io_B_Valid_41_39;
    _zz_io_MatrixB_42 <= SubModule_WeightCache_mData_42;
    _zz_io_MatrixB_42_1 <= _zz_io_MatrixB_42;
    _zz_io_MatrixB_42_2 <= _zz_io_MatrixB_42_1;
    _zz_io_MatrixB_42_3 <= _zz_io_MatrixB_42_2;
    _zz_io_MatrixB_42_4 <= _zz_io_MatrixB_42_3;
    _zz_io_MatrixB_42_5 <= _zz_io_MatrixB_42_4;
    _zz_io_MatrixB_42_6 <= _zz_io_MatrixB_42_5;
    _zz_io_MatrixB_42_7 <= _zz_io_MatrixB_42_6;
    _zz_io_MatrixB_42_8 <= _zz_io_MatrixB_42_7;
    _zz_io_MatrixB_42_9 <= _zz_io_MatrixB_42_8;
    _zz_io_MatrixB_42_10 <= _zz_io_MatrixB_42_9;
    _zz_io_MatrixB_42_11 <= _zz_io_MatrixB_42_10;
    _zz_io_MatrixB_42_12 <= _zz_io_MatrixB_42_11;
    _zz_io_MatrixB_42_13 <= _zz_io_MatrixB_42_12;
    _zz_io_MatrixB_42_14 <= _zz_io_MatrixB_42_13;
    _zz_io_MatrixB_42_15 <= _zz_io_MatrixB_42_14;
    _zz_io_MatrixB_42_16 <= _zz_io_MatrixB_42_15;
    _zz_io_MatrixB_42_17 <= _zz_io_MatrixB_42_16;
    _zz_io_MatrixB_42_18 <= _zz_io_MatrixB_42_17;
    _zz_io_MatrixB_42_19 <= _zz_io_MatrixB_42_18;
    _zz_io_MatrixB_42_20 <= _zz_io_MatrixB_42_19;
    _zz_io_MatrixB_42_21 <= _zz_io_MatrixB_42_20;
    _zz_io_MatrixB_42_22 <= _zz_io_MatrixB_42_21;
    _zz_io_MatrixB_42_23 <= _zz_io_MatrixB_42_22;
    _zz_io_MatrixB_42_24 <= _zz_io_MatrixB_42_23;
    _zz_io_MatrixB_42_25 <= _zz_io_MatrixB_42_24;
    _zz_io_MatrixB_42_26 <= _zz_io_MatrixB_42_25;
    _zz_io_MatrixB_42_27 <= _zz_io_MatrixB_42_26;
    _zz_io_MatrixB_42_28 <= _zz_io_MatrixB_42_27;
    _zz_io_MatrixB_42_29 <= _zz_io_MatrixB_42_28;
    _zz_io_MatrixB_42_30 <= _zz_io_MatrixB_42_29;
    _zz_io_MatrixB_42_31 <= _zz_io_MatrixB_42_30;
    _zz_io_MatrixB_42_32 <= _zz_io_MatrixB_42_31;
    _zz_io_MatrixB_42_33 <= _zz_io_MatrixB_42_32;
    _zz_io_MatrixB_42_34 <= _zz_io_MatrixB_42_33;
    _zz_io_MatrixB_42_35 <= _zz_io_MatrixB_42_34;
    _zz_io_MatrixB_42_36 <= _zz_io_MatrixB_42_35;
    _zz_io_MatrixB_42_37 <= _zz_io_MatrixB_42_36;
    _zz_io_MatrixB_42_38 <= _zz_io_MatrixB_42_37;
    _zz_io_MatrixB_42_39 <= _zz_io_MatrixB_42_38;
    _zz_io_MatrixB_42_40 <= _zz_io_MatrixB_42_39;
    _zz_io_MatrixB_42_41 <= _zz_io_MatrixB_42_40;
    _zz_io_B_Valid_42 <= SubModule_WeightCache_MatrixCol_Switch[42];
    _zz_io_B_Valid_42_1 <= _zz_io_B_Valid_42;
    _zz_io_B_Valid_42_2 <= _zz_io_B_Valid_42_1;
    _zz_io_B_Valid_42_3 <= _zz_io_B_Valid_42_2;
    _zz_io_B_Valid_42_4 <= _zz_io_B_Valid_42_3;
    _zz_io_B_Valid_42_5 <= _zz_io_B_Valid_42_4;
    _zz_io_B_Valid_42_6 <= _zz_io_B_Valid_42_5;
    _zz_io_B_Valid_42_7 <= _zz_io_B_Valid_42_6;
    _zz_io_B_Valid_42_8 <= _zz_io_B_Valid_42_7;
    _zz_io_B_Valid_42_9 <= _zz_io_B_Valid_42_8;
    _zz_io_B_Valid_42_10 <= _zz_io_B_Valid_42_9;
    _zz_io_B_Valid_42_11 <= _zz_io_B_Valid_42_10;
    _zz_io_B_Valid_42_12 <= _zz_io_B_Valid_42_11;
    _zz_io_B_Valid_42_13 <= _zz_io_B_Valid_42_12;
    _zz_io_B_Valid_42_14 <= _zz_io_B_Valid_42_13;
    _zz_io_B_Valid_42_15 <= _zz_io_B_Valid_42_14;
    _zz_io_B_Valid_42_16 <= _zz_io_B_Valid_42_15;
    _zz_io_B_Valid_42_17 <= _zz_io_B_Valid_42_16;
    _zz_io_B_Valid_42_18 <= _zz_io_B_Valid_42_17;
    _zz_io_B_Valid_42_19 <= _zz_io_B_Valid_42_18;
    _zz_io_B_Valid_42_20 <= _zz_io_B_Valid_42_19;
    _zz_io_B_Valid_42_21 <= _zz_io_B_Valid_42_20;
    _zz_io_B_Valid_42_22 <= _zz_io_B_Valid_42_21;
    _zz_io_B_Valid_42_23 <= _zz_io_B_Valid_42_22;
    _zz_io_B_Valid_42_24 <= _zz_io_B_Valid_42_23;
    _zz_io_B_Valid_42_25 <= _zz_io_B_Valid_42_24;
    _zz_io_B_Valid_42_26 <= _zz_io_B_Valid_42_25;
    _zz_io_B_Valid_42_27 <= _zz_io_B_Valid_42_26;
    _zz_io_B_Valid_42_28 <= _zz_io_B_Valid_42_27;
    _zz_io_B_Valid_42_29 <= _zz_io_B_Valid_42_28;
    _zz_io_B_Valid_42_30 <= _zz_io_B_Valid_42_29;
    _zz_io_B_Valid_42_31 <= _zz_io_B_Valid_42_30;
    _zz_io_B_Valid_42_32 <= _zz_io_B_Valid_42_31;
    _zz_io_B_Valid_42_33 <= _zz_io_B_Valid_42_32;
    _zz_io_B_Valid_42_34 <= _zz_io_B_Valid_42_33;
    _zz_io_B_Valid_42_35 <= _zz_io_B_Valid_42_34;
    _zz_io_B_Valid_42_36 <= _zz_io_B_Valid_42_35;
    _zz_io_B_Valid_42_37 <= _zz_io_B_Valid_42_36;
    _zz_io_B_Valid_42_38 <= _zz_io_B_Valid_42_37;
    _zz_io_B_Valid_42_39 <= _zz_io_B_Valid_42_38;
    _zz_io_B_Valid_42_40 <= _zz_io_B_Valid_42_39;
    _zz_io_B_Valid_42_41 <= _zz_io_B_Valid_42_40;
    _zz_io_MatrixB_43 <= SubModule_WeightCache_mData_43;
    _zz_io_MatrixB_43_1 <= _zz_io_MatrixB_43;
    _zz_io_MatrixB_43_2 <= _zz_io_MatrixB_43_1;
    _zz_io_MatrixB_43_3 <= _zz_io_MatrixB_43_2;
    _zz_io_MatrixB_43_4 <= _zz_io_MatrixB_43_3;
    _zz_io_MatrixB_43_5 <= _zz_io_MatrixB_43_4;
    _zz_io_MatrixB_43_6 <= _zz_io_MatrixB_43_5;
    _zz_io_MatrixB_43_7 <= _zz_io_MatrixB_43_6;
    _zz_io_MatrixB_43_8 <= _zz_io_MatrixB_43_7;
    _zz_io_MatrixB_43_9 <= _zz_io_MatrixB_43_8;
    _zz_io_MatrixB_43_10 <= _zz_io_MatrixB_43_9;
    _zz_io_MatrixB_43_11 <= _zz_io_MatrixB_43_10;
    _zz_io_MatrixB_43_12 <= _zz_io_MatrixB_43_11;
    _zz_io_MatrixB_43_13 <= _zz_io_MatrixB_43_12;
    _zz_io_MatrixB_43_14 <= _zz_io_MatrixB_43_13;
    _zz_io_MatrixB_43_15 <= _zz_io_MatrixB_43_14;
    _zz_io_MatrixB_43_16 <= _zz_io_MatrixB_43_15;
    _zz_io_MatrixB_43_17 <= _zz_io_MatrixB_43_16;
    _zz_io_MatrixB_43_18 <= _zz_io_MatrixB_43_17;
    _zz_io_MatrixB_43_19 <= _zz_io_MatrixB_43_18;
    _zz_io_MatrixB_43_20 <= _zz_io_MatrixB_43_19;
    _zz_io_MatrixB_43_21 <= _zz_io_MatrixB_43_20;
    _zz_io_MatrixB_43_22 <= _zz_io_MatrixB_43_21;
    _zz_io_MatrixB_43_23 <= _zz_io_MatrixB_43_22;
    _zz_io_MatrixB_43_24 <= _zz_io_MatrixB_43_23;
    _zz_io_MatrixB_43_25 <= _zz_io_MatrixB_43_24;
    _zz_io_MatrixB_43_26 <= _zz_io_MatrixB_43_25;
    _zz_io_MatrixB_43_27 <= _zz_io_MatrixB_43_26;
    _zz_io_MatrixB_43_28 <= _zz_io_MatrixB_43_27;
    _zz_io_MatrixB_43_29 <= _zz_io_MatrixB_43_28;
    _zz_io_MatrixB_43_30 <= _zz_io_MatrixB_43_29;
    _zz_io_MatrixB_43_31 <= _zz_io_MatrixB_43_30;
    _zz_io_MatrixB_43_32 <= _zz_io_MatrixB_43_31;
    _zz_io_MatrixB_43_33 <= _zz_io_MatrixB_43_32;
    _zz_io_MatrixB_43_34 <= _zz_io_MatrixB_43_33;
    _zz_io_MatrixB_43_35 <= _zz_io_MatrixB_43_34;
    _zz_io_MatrixB_43_36 <= _zz_io_MatrixB_43_35;
    _zz_io_MatrixB_43_37 <= _zz_io_MatrixB_43_36;
    _zz_io_MatrixB_43_38 <= _zz_io_MatrixB_43_37;
    _zz_io_MatrixB_43_39 <= _zz_io_MatrixB_43_38;
    _zz_io_MatrixB_43_40 <= _zz_io_MatrixB_43_39;
    _zz_io_MatrixB_43_41 <= _zz_io_MatrixB_43_40;
    _zz_io_MatrixB_43_42 <= _zz_io_MatrixB_43_41;
    _zz_io_B_Valid_43 <= SubModule_WeightCache_MatrixCol_Switch[43];
    _zz_io_B_Valid_43_1 <= _zz_io_B_Valid_43;
    _zz_io_B_Valid_43_2 <= _zz_io_B_Valid_43_1;
    _zz_io_B_Valid_43_3 <= _zz_io_B_Valid_43_2;
    _zz_io_B_Valid_43_4 <= _zz_io_B_Valid_43_3;
    _zz_io_B_Valid_43_5 <= _zz_io_B_Valid_43_4;
    _zz_io_B_Valid_43_6 <= _zz_io_B_Valid_43_5;
    _zz_io_B_Valid_43_7 <= _zz_io_B_Valid_43_6;
    _zz_io_B_Valid_43_8 <= _zz_io_B_Valid_43_7;
    _zz_io_B_Valid_43_9 <= _zz_io_B_Valid_43_8;
    _zz_io_B_Valid_43_10 <= _zz_io_B_Valid_43_9;
    _zz_io_B_Valid_43_11 <= _zz_io_B_Valid_43_10;
    _zz_io_B_Valid_43_12 <= _zz_io_B_Valid_43_11;
    _zz_io_B_Valid_43_13 <= _zz_io_B_Valid_43_12;
    _zz_io_B_Valid_43_14 <= _zz_io_B_Valid_43_13;
    _zz_io_B_Valid_43_15 <= _zz_io_B_Valid_43_14;
    _zz_io_B_Valid_43_16 <= _zz_io_B_Valid_43_15;
    _zz_io_B_Valid_43_17 <= _zz_io_B_Valid_43_16;
    _zz_io_B_Valid_43_18 <= _zz_io_B_Valid_43_17;
    _zz_io_B_Valid_43_19 <= _zz_io_B_Valid_43_18;
    _zz_io_B_Valid_43_20 <= _zz_io_B_Valid_43_19;
    _zz_io_B_Valid_43_21 <= _zz_io_B_Valid_43_20;
    _zz_io_B_Valid_43_22 <= _zz_io_B_Valid_43_21;
    _zz_io_B_Valid_43_23 <= _zz_io_B_Valid_43_22;
    _zz_io_B_Valid_43_24 <= _zz_io_B_Valid_43_23;
    _zz_io_B_Valid_43_25 <= _zz_io_B_Valid_43_24;
    _zz_io_B_Valid_43_26 <= _zz_io_B_Valid_43_25;
    _zz_io_B_Valid_43_27 <= _zz_io_B_Valid_43_26;
    _zz_io_B_Valid_43_28 <= _zz_io_B_Valid_43_27;
    _zz_io_B_Valid_43_29 <= _zz_io_B_Valid_43_28;
    _zz_io_B_Valid_43_30 <= _zz_io_B_Valid_43_29;
    _zz_io_B_Valid_43_31 <= _zz_io_B_Valid_43_30;
    _zz_io_B_Valid_43_32 <= _zz_io_B_Valid_43_31;
    _zz_io_B_Valid_43_33 <= _zz_io_B_Valid_43_32;
    _zz_io_B_Valid_43_34 <= _zz_io_B_Valid_43_33;
    _zz_io_B_Valid_43_35 <= _zz_io_B_Valid_43_34;
    _zz_io_B_Valid_43_36 <= _zz_io_B_Valid_43_35;
    _zz_io_B_Valid_43_37 <= _zz_io_B_Valid_43_36;
    _zz_io_B_Valid_43_38 <= _zz_io_B_Valid_43_37;
    _zz_io_B_Valid_43_39 <= _zz_io_B_Valid_43_38;
    _zz_io_B_Valid_43_40 <= _zz_io_B_Valid_43_39;
    _zz_io_B_Valid_43_41 <= _zz_io_B_Valid_43_40;
    _zz_io_B_Valid_43_42 <= _zz_io_B_Valid_43_41;
    _zz_io_MatrixB_44 <= SubModule_WeightCache_mData_44;
    _zz_io_MatrixB_44_1 <= _zz_io_MatrixB_44;
    _zz_io_MatrixB_44_2 <= _zz_io_MatrixB_44_1;
    _zz_io_MatrixB_44_3 <= _zz_io_MatrixB_44_2;
    _zz_io_MatrixB_44_4 <= _zz_io_MatrixB_44_3;
    _zz_io_MatrixB_44_5 <= _zz_io_MatrixB_44_4;
    _zz_io_MatrixB_44_6 <= _zz_io_MatrixB_44_5;
    _zz_io_MatrixB_44_7 <= _zz_io_MatrixB_44_6;
    _zz_io_MatrixB_44_8 <= _zz_io_MatrixB_44_7;
    _zz_io_MatrixB_44_9 <= _zz_io_MatrixB_44_8;
    _zz_io_MatrixB_44_10 <= _zz_io_MatrixB_44_9;
    _zz_io_MatrixB_44_11 <= _zz_io_MatrixB_44_10;
    _zz_io_MatrixB_44_12 <= _zz_io_MatrixB_44_11;
    _zz_io_MatrixB_44_13 <= _zz_io_MatrixB_44_12;
    _zz_io_MatrixB_44_14 <= _zz_io_MatrixB_44_13;
    _zz_io_MatrixB_44_15 <= _zz_io_MatrixB_44_14;
    _zz_io_MatrixB_44_16 <= _zz_io_MatrixB_44_15;
    _zz_io_MatrixB_44_17 <= _zz_io_MatrixB_44_16;
    _zz_io_MatrixB_44_18 <= _zz_io_MatrixB_44_17;
    _zz_io_MatrixB_44_19 <= _zz_io_MatrixB_44_18;
    _zz_io_MatrixB_44_20 <= _zz_io_MatrixB_44_19;
    _zz_io_MatrixB_44_21 <= _zz_io_MatrixB_44_20;
    _zz_io_MatrixB_44_22 <= _zz_io_MatrixB_44_21;
    _zz_io_MatrixB_44_23 <= _zz_io_MatrixB_44_22;
    _zz_io_MatrixB_44_24 <= _zz_io_MatrixB_44_23;
    _zz_io_MatrixB_44_25 <= _zz_io_MatrixB_44_24;
    _zz_io_MatrixB_44_26 <= _zz_io_MatrixB_44_25;
    _zz_io_MatrixB_44_27 <= _zz_io_MatrixB_44_26;
    _zz_io_MatrixB_44_28 <= _zz_io_MatrixB_44_27;
    _zz_io_MatrixB_44_29 <= _zz_io_MatrixB_44_28;
    _zz_io_MatrixB_44_30 <= _zz_io_MatrixB_44_29;
    _zz_io_MatrixB_44_31 <= _zz_io_MatrixB_44_30;
    _zz_io_MatrixB_44_32 <= _zz_io_MatrixB_44_31;
    _zz_io_MatrixB_44_33 <= _zz_io_MatrixB_44_32;
    _zz_io_MatrixB_44_34 <= _zz_io_MatrixB_44_33;
    _zz_io_MatrixB_44_35 <= _zz_io_MatrixB_44_34;
    _zz_io_MatrixB_44_36 <= _zz_io_MatrixB_44_35;
    _zz_io_MatrixB_44_37 <= _zz_io_MatrixB_44_36;
    _zz_io_MatrixB_44_38 <= _zz_io_MatrixB_44_37;
    _zz_io_MatrixB_44_39 <= _zz_io_MatrixB_44_38;
    _zz_io_MatrixB_44_40 <= _zz_io_MatrixB_44_39;
    _zz_io_MatrixB_44_41 <= _zz_io_MatrixB_44_40;
    _zz_io_MatrixB_44_42 <= _zz_io_MatrixB_44_41;
    _zz_io_MatrixB_44_43 <= _zz_io_MatrixB_44_42;
    _zz_io_B_Valid_44 <= SubModule_WeightCache_MatrixCol_Switch[44];
    _zz_io_B_Valid_44_1 <= _zz_io_B_Valid_44;
    _zz_io_B_Valid_44_2 <= _zz_io_B_Valid_44_1;
    _zz_io_B_Valid_44_3 <= _zz_io_B_Valid_44_2;
    _zz_io_B_Valid_44_4 <= _zz_io_B_Valid_44_3;
    _zz_io_B_Valid_44_5 <= _zz_io_B_Valid_44_4;
    _zz_io_B_Valid_44_6 <= _zz_io_B_Valid_44_5;
    _zz_io_B_Valid_44_7 <= _zz_io_B_Valid_44_6;
    _zz_io_B_Valid_44_8 <= _zz_io_B_Valid_44_7;
    _zz_io_B_Valid_44_9 <= _zz_io_B_Valid_44_8;
    _zz_io_B_Valid_44_10 <= _zz_io_B_Valid_44_9;
    _zz_io_B_Valid_44_11 <= _zz_io_B_Valid_44_10;
    _zz_io_B_Valid_44_12 <= _zz_io_B_Valid_44_11;
    _zz_io_B_Valid_44_13 <= _zz_io_B_Valid_44_12;
    _zz_io_B_Valid_44_14 <= _zz_io_B_Valid_44_13;
    _zz_io_B_Valid_44_15 <= _zz_io_B_Valid_44_14;
    _zz_io_B_Valid_44_16 <= _zz_io_B_Valid_44_15;
    _zz_io_B_Valid_44_17 <= _zz_io_B_Valid_44_16;
    _zz_io_B_Valid_44_18 <= _zz_io_B_Valid_44_17;
    _zz_io_B_Valid_44_19 <= _zz_io_B_Valid_44_18;
    _zz_io_B_Valid_44_20 <= _zz_io_B_Valid_44_19;
    _zz_io_B_Valid_44_21 <= _zz_io_B_Valid_44_20;
    _zz_io_B_Valid_44_22 <= _zz_io_B_Valid_44_21;
    _zz_io_B_Valid_44_23 <= _zz_io_B_Valid_44_22;
    _zz_io_B_Valid_44_24 <= _zz_io_B_Valid_44_23;
    _zz_io_B_Valid_44_25 <= _zz_io_B_Valid_44_24;
    _zz_io_B_Valid_44_26 <= _zz_io_B_Valid_44_25;
    _zz_io_B_Valid_44_27 <= _zz_io_B_Valid_44_26;
    _zz_io_B_Valid_44_28 <= _zz_io_B_Valid_44_27;
    _zz_io_B_Valid_44_29 <= _zz_io_B_Valid_44_28;
    _zz_io_B_Valid_44_30 <= _zz_io_B_Valid_44_29;
    _zz_io_B_Valid_44_31 <= _zz_io_B_Valid_44_30;
    _zz_io_B_Valid_44_32 <= _zz_io_B_Valid_44_31;
    _zz_io_B_Valid_44_33 <= _zz_io_B_Valid_44_32;
    _zz_io_B_Valid_44_34 <= _zz_io_B_Valid_44_33;
    _zz_io_B_Valid_44_35 <= _zz_io_B_Valid_44_34;
    _zz_io_B_Valid_44_36 <= _zz_io_B_Valid_44_35;
    _zz_io_B_Valid_44_37 <= _zz_io_B_Valid_44_36;
    _zz_io_B_Valid_44_38 <= _zz_io_B_Valid_44_37;
    _zz_io_B_Valid_44_39 <= _zz_io_B_Valid_44_38;
    _zz_io_B_Valid_44_40 <= _zz_io_B_Valid_44_39;
    _zz_io_B_Valid_44_41 <= _zz_io_B_Valid_44_40;
    _zz_io_B_Valid_44_42 <= _zz_io_B_Valid_44_41;
    _zz_io_B_Valid_44_43 <= _zz_io_B_Valid_44_42;
    _zz_io_MatrixB_45 <= SubModule_WeightCache_mData_45;
    _zz_io_MatrixB_45_1 <= _zz_io_MatrixB_45;
    _zz_io_MatrixB_45_2 <= _zz_io_MatrixB_45_1;
    _zz_io_MatrixB_45_3 <= _zz_io_MatrixB_45_2;
    _zz_io_MatrixB_45_4 <= _zz_io_MatrixB_45_3;
    _zz_io_MatrixB_45_5 <= _zz_io_MatrixB_45_4;
    _zz_io_MatrixB_45_6 <= _zz_io_MatrixB_45_5;
    _zz_io_MatrixB_45_7 <= _zz_io_MatrixB_45_6;
    _zz_io_MatrixB_45_8 <= _zz_io_MatrixB_45_7;
    _zz_io_MatrixB_45_9 <= _zz_io_MatrixB_45_8;
    _zz_io_MatrixB_45_10 <= _zz_io_MatrixB_45_9;
    _zz_io_MatrixB_45_11 <= _zz_io_MatrixB_45_10;
    _zz_io_MatrixB_45_12 <= _zz_io_MatrixB_45_11;
    _zz_io_MatrixB_45_13 <= _zz_io_MatrixB_45_12;
    _zz_io_MatrixB_45_14 <= _zz_io_MatrixB_45_13;
    _zz_io_MatrixB_45_15 <= _zz_io_MatrixB_45_14;
    _zz_io_MatrixB_45_16 <= _zz_io_MatrixB_45_15;
    _zz_io_MatrixB_45_17 <= _zz_io_MatrixB_45_16;
    _zz_io_MatrixB_45_18 <= _zz_io_MatrixB_45_17;
    _zz_io_MatrixB_45_19 <= _zz_io_MatrixB_45_18;
    _zz_io_MatrixB_45_20 <= _zz_io_MatrixB_45_19;
    _zz_io_MatrixB_45_21 <= _zz_io_MatrixB_45_20;
    _zz_io_MatrixB_45_22 <= _zz_io_MatrixB_45_21;
    _zz_io_MatrixB_45_23 <= _zz_io_MatrixB_45_22;
    _zz_io_MatrixB_45_24 <= _zz_io_MatrixB_45_23;
    _zz_io_MatrixB_45_25 <= _zz_io_MatrixB_45_24;
    _zz_io_MatrixB_45_26 <= _zz_io_MatrixB_45_25;
    _zz_io_MatrixB_45_27 <= _zz_io_MatrixB_45_26;
    _zz_io_MatrixB_45_28 <= _zz_io_MatrixB_45_27;
    _zz_io_MatrixB_45_29 <= _zz_io_MatrixB_45_28;
    _zz_io_MatrixB_45_30 <= _zz_io_MatrixB_45_29;
    _zz_io_MatrixB_45_31 <= _zz_io_MatrixB_45_30;
    _zz_io_MatrixB_45_32 <= _zz_io_MatrixB_45_31;
    _zz_io_MatrixB_45_33 <= _zz_io_MatrixB_45_32;
    _zz_io_MatrixB_45_34 <= _zz_io_MatrixB_45_33;
    _zz_io_MatrixB_45_35 <= _zz_io_MatrixB_45_34;
    _zz_io_MatrixB_45_36 <= _zz_io_MatrixB_45_35;
    _zz_io_MatrixB_45_37 <= _zz_io_MatrixB_45_36;
    _zz_io_MatrixB_45_38 <= _zz_io_MatrixB_45_37;
    _zz_io_MatrixB_45_39 <= _zz_io_MatrixB_45_38;
    _zz_io_MatrixB_45_40 <= _zz_io_MatrixB_45_39;
    _zz_io_MatrixB_45_41 <= _zz_io_MatrixB_45_40;
    _zz_io_MatrixB_45_42 <= _zz_io_MatrixB_45_41;
    _zz_io_MatrixB_45_43 <= _zz_io_MatrixB_45_42;
    _zz_io_MatrixB_45_44 <= _zz_io_MatrixB_45_43;
    _zz_io_B_Valid_45 <= SubModule_WeightCache_MatrixCol_Switch[45];
    _zz_io_B_Valid_45_1 <= _zz_io_B_Valid_45;
    _zz_io_B_Valid_45_2 <= _zz_io_B_Valid_45_1;
    _zz_io_B_Valid_45_3 <= _zz_io_B_Valid_45_2;
    _zz_io_B_Valid_45_4 <= _zz_io_B_Valid_45_3;
    _zz_io_B_Valid_45_5 <= _zz_io_B_Valid_45_4;
    _zz_io_B_Valid_45_6 <= _zz_io_B_Valid_45_5;
    _zz_io_B_Valid_45_7 <= _zz_io_B_Valid_45_6;
    _zz_io_B_Valid_45_8 <= _zz_io_B_Valid_45_7;
    _zz_io_B_Valid_45_9 <= _zz_io_B_Valid_45_8;
    _zz_io_B_Valid_45_10 <= _zz_io_B_Valid_45_9;
    _zz_io_B_Valid_45_11 <= _zz_io_B_Valid_45_10;
    _zz_io_B_Valid_45_12 <= _zz_io_B_Valid_45_11;
    _zz_io_B_Valid_45_13 <= _zz_io_B_Valid_45_12;
    _zz_io_B_Valid_45_14 <= _zz_io_B_Valid_45_13;
    _zz_io_B_Valid_45_15 <= _zz_io_B_Valid_45_14;
    _zz_io_B_Valid_45_16 <= _zz_io_B_Valid_45_15;
    _zz_io_B_Valid_45_17 <= _zz_io_B_Valid_45_16;
    _zz_io_B_Valid_45_18 <= _zz_io_B_Valid_45_17;
    _zz_io_B_Valid_45_19 <= _zz_io_B_Valid_45_18;
    _zz_io_B_Valid_45_20 <= _zz_io_B_Valid_45_19;
    _zz_io_B_Valid_45_21 <= _zz_io_B_Valid_45_20;
    _zz_io_B_Valid_45_22 <= _zz_io_B_Valid_45_21;
    _zz_io_B_Valid_45_23 <= _zz_io_B_Valid_45_22;
    _zz_io_B_Valid_45_24 <= _zz_io_B_Valid_45_23;
    _zz_io_B_Valid_45_25 <= _zz_io_B_Valid_45_24;
    _zz_io_B_Valid_45_26 <= _zz_io_B_Valid_45_25;
    _zz_io_B_Valid_45_27 <= _zz_io_B_Valid_45_26;
    _zz_io_B_Valid_45_28 <= _zz_io_B_Valid_45_27;
    _zz_io_B_Valid_45_29 <= _zz_io_B_Valid_45_28;
    _zz_io_B_Valid_45_30 <= _zz_io_B_Valid_45_29;
    _zz_io_B_Valid_45_31 <= _zz_io_B_Valid_45_30;
    _zz_io_B_Valid_45_32 <= _zz_io_B_Valid_45_31;
    _zz_io_B_Valid_45_33 <= _zz_io_B_Valid_45_32;
    _zz_io_B_Valid_45_34 <= _zz_io_B_Valid_45_33;
    _zz_io_B_Valid_45_35 <= _zz_io_B_Valid_45_34;
    _zz_io_B_Valid_45_36 <= _zz_io_B_Valid_45_35;
    _zz_io_B_Valid_45_37 <= _zz_io_B_Valid_45_36;
    _zz_io_B_Valid_45_38 <= _zz_io_B_Valid_45_37;
    _zz_io_B_Valid_45_39 <= _zz_io_B_Valid_45_38;
    _zz_io_B_Valid_45_40 <= _zz_io_B_Valid_45_39;
    _zz_io_B_Valid_45_41 <= _zz_io_B_Valid_45_40;
    _zz_io_B_Valid_45_42 <= _zz_io_B_Valid_45_41;
    _zz_io_B_Valid_45_43 <= _zz_io_B_Valid_45_42;
    _zz_io_B_Valid_45_44 <= _zz_io_B_Valid_45_43;
    _zz_io_MatrixB_46 <= SubModule_WeightCache_mData_46;
    _zz_io_MatrixB_46_1 <= _zz_io_MatrixB_46;
    _zz_io_MatrixB_46_2 <= _zz_io_MatrixB_46_1;
    _zz_io_MatrixB_46_3 <= _zz_io_MatrixB_46_2;
    _zz_io_MatrixB_46_4 <= _zz_io_MatrixB_46_3;
    _zz_io_MatrixB_46_5 <= _zz_io_MatrixB_46_4;
    _zz_io_MatrixB_46_6 <= _zz_io_MatrixB_46_5;
    _zz_io_MatrixB_46_7 <= _zz_io_MatrixB_46_6;
    _zz_io_MatrixB_46_8 <= _zz_io_MatrixB_46_7;
    _zz_io_MatrixB_46_9 <= _zz_io_MatrixB_46_8;
    _zz_io_MatrixB_46_10 <= _zz_io_MatrixB_46_9;
    _zz_io_MatrixB_46_11 <= _zz_io_MatrixB_46_10;
    _zz_io_MatrixB_46_12 <= _zz_io_MatrixB_46_11;
    _zz_io_MatrixB_46_13 <= _zz_io_MatrixB_46_12;
    _zz_io_MatrixB_46_14 <= _zz_io_MatrixB_46_13;
    _zz_io_MatrixB_46_15 <= _zz_io_MatrixB_46_14;
    _zz_io_MatrixB_46_16 <= _zz_io_MatrixB_46_15;
    _zz_io_MatrixB_46_17 <= _zz_io_MatrixB_46_16;
    _zz_io_MatrixB_46_18 <= _zz_io_MatrixB_46_17;
    _zz_io_MatrixB_46_19 <= _zz_io_MatrixB_46_18;
    _zz_io_MatrixB_46_20 <= _zz_io_MatrixB_46_19;
    _zz_io_MatrixB_46_21 <= _zz_io_MatrixB_46_20;
    _zz_io_MatrixB_46_22 <= _zz_io_MatrixB_46_21;
    _zz_io_MatrixB_46_23 <= _zz_io_MatrixB_46_22;
    _zz_io_MatrixB_46_24 <= _zz_io_MatrixB_46_23;
    _zz_io_MatrixB_46_25 <= _zz_io_MatrixB_46_24;
    _zz_io_MatrixB_46_26 <= _zz_io_MatrixB_46_25;
    _zz_io_MatrixB_46_27 <= _zz_io_MatrixB_46_26;
    _zz_io_MatrixB_46_28 <= _zz_io_MatrixB_46_27;
    _zz_io_MatrixB_46_29 <= _zz_io_MatrixB_46_28;
    _zz_io_MatrixB_46_30 <= _zz_io_MatrixB_46_29;
    _zz_io_MatrixB_46_31 <= _zz_io_MatrixB_46_30;
    _zz_io_MatrixB_46_32 <= _zz_io_MatrixB_46_31;
    _zz_io_MatrixB_46_33 <= _zz_io_MatrixB_46_32;
    _zz_io_MatrixB_46_34 <= _zz_io_MatrixB_46_33;
    _zz_io_MatrixB_46_35 <= _zz_io_MatrixB_46_34;
    _zz_io_MatrixB_46_36 <= _zz_io_MatrixB_46_35;
    _zz_io_MatrixB_46_37 <= _zz_io_MatrixB_46_36;
    _zz_io_MatrixB_46_38 <= _zz_io_MatrixB_46_37;
    _zz_io_MatrixB_46_39 <= _zz_io_MatrixB_46_38;
    _zz_io_MatrixB_46_40 <= _zz_io_MatrixB_46_39;
    _zz_io_MatrixB_46_41 <= _zz_io_MatrixB_46_40;
    _zz_io_MatrixB_46_42 <= _zz_io_MatrixB_46_41;
    _zz_io_MatrixB_46_43 <= _zz_io_MatrixB_46_42;
    _zz_io_MatrixB_46_44 <= _zz_io_MatrixB_46_43;
    _zz_io_MatrixB_46_45 <= _zz_io_MatrixB_46_44;
    _zz_io_B_Valid_46 <= SubModule_WeightCache_MatrixCol_Switch[46];
    _zz_io_B_Valid_46_1 <= _zz_io_B_Valid_46;
    _zz_io_B_Valid_46_2 <= _zz_io_B_Valid_46_1;
    _zz_io_B_Valid_46_3 <= _zz_io_B_Valid_46_2;
    _zz_io_B_Valid_46_4 <= _zz_io_B_Valid_46_3;
    _zz_io_B_Valid_46_5 <= _zz_io_B_Valid_46_4;
    _zz_io_B_Valid_46_6 <= _zz_io_B_Valid_46_5;
    _zz_io_B_Valid_46_7 <= _zz_io_B_Valid_46_6;
    _zz_io_B_Valid_46_8 <= _zz_io_B_Valid_46_7;
    _zz_io_B_Valid_46_9 <= _zz_io_B_Valid_46_8;
    _zz_io_B_Valid_46_10 <= _zz_io_B_Valid_46_9;
    _zz_io_B_Valid_46_11 <= _zz_io_B_Valid_46_10;
    _zz_io_B_Valid_46_12 <= _zz_io_B_Valid_46_11;
    _zz_io_B_Valid_46_13 <= _zz_io_B_Valid_46_12;
    _zz_io_B_Valid_46_14 <= _zz_io_B_Valid_46_13;
    _zz_io_B_Valid_46_15 <= _zz_io_B_Valid_46_14;
    _zz_io_B_Valid_46_16 <= _zz_io_B_Valid_46_15;
    _zz_io_B_Valid_46_17 <= _zz_io_B_Valid_46_16;
    _zz_io_B_Valid_46_18 <= _zz_io_B_Valid_46_17;
    _zz_io_B_Valid_46_19 <= _zz_io_B_Valid_46_18;
    _zz_io_B_Valid_46_20 <= _zz_io_B_Valid_46_19;
    _zz_io_B_Valid_46_21 <= _zz_io_B_Valid_46_20;
    _zz_io_B_Valid_46_22 <= _zz_io_B_Valid_46_21;
    _zz_io_B_Valid_46_23 <= _zz_io_B_Valid_46_22;
    _zz_io_B_Valid_46_24 <= _zz_io_B_Valid_46_23;
    _zz_io_B_Valid_46_25 <= _zz_io_B_Valid_46_24;
    _zz_io_B_Valid_46_26 <= _zz_io_B_Valid_46_25;
    _zz_io_B_Valid_46_27 <= _zz_io_B_Valid_46_26;
    _zz_io_B_Valid_46_28 <= _zz_io_B_Valid_46_27;
    _zz_io_B_Valid_46_29 <= _zz_io_B_Valid_46_28;
    _zz_io_B_Valid_46_30 <= _zz_io_B_Valid_46_29;
    _zz_io_B_Valid_46_31 <= _zz_io_B_Valid_46_30;
    _zz_io_B_Valid_46_32 <= _zz_io_B_Valid_46_31;
    _zz_io_B_Valid_46_33 <= _zz_io_B_Valid_46_32;
    _zz_io_B_Valid_46_34 <= _zz_io_B_Valid_46_33;
    _zz_io_B_Valid_46_35 <= _zz_io_B_Valid_46_34;
    _zz_io_B_Valid_46_36 <= _zz_io_B_Valid_46_35;
    _zz_io_B_Valid_46_37 <= _zz_io_B_Valid_46_36;
    _zz_io_B_Valid_46_38 <= _zz_io_B_Valid_46_37;
    _zz_io_B_Valid_46_39 <= _zz_io_B_Valid_46_38;
    _zz_io_B_Valid_46_40 <= _zz_io_B_Valid_46_39;
    _zz_io_B_Valid_46_41 <= _zz_io_B_Valid_46_40;
    _zz_io_B_Valid_46_42 <= _zz_io_B_Valid_46_41;
    _zz_io_B_Valid_46_43 <= _zz_io_B_Valid_46_42;
    _zz_io_B_Valid_46_44 <= _zz_io_B_Valid_46_43;
    _zz_io_B_Valid_46_45 <= _zz_io_B_Valid_46_44;
    _zz_io_MatrixB_47 <= SubModule_WeightCache_mData_47;
    _zz_io_MatrixB_47_1 <= _zz_io_MatrixB_47;
    _zz_io_MatrixB_47_2 <= _zz_io_MatrixB_47_1;
    _zz_io_MatrixB_47_3 <= _zz_io_MatrixB_47_2;
    _zz_io_MatrixB_47_4 <= _zz_io_MatrixB_47_3;
    _zz_io_MatrixB_47_5 <= _zz_io_MatrixB_47_4;
    _zz_io_MatrixB_47_6 <= _zz_io_MatrixB_47_5;
    _zz_io_MatrixB_47_7 <= _zz_io_MatrixB_47_6;
    _zz_io_MatrixB_47_8 <= _zz_io_MatrixB_47_7;
    _zz_io_MatrixB_47_9 <= _zz_io_MatrixB_47_8;
    _zz_io_MatrixB_47_10 <= _zz_io_MatrixB_47_9;
    _zz_io_MatrixB_47_11 <= _zz_io_MatrixB_47_10;
    _zz_io_MatrixB_47_12 <= _zz_io_MatrixB_47_11;
    _zz_io_MatrixB_47_13 <= _zz_io_MatrixB_47_12;
    _zz_io_MatrixB_47_14 <= _zz_io_MatrixB_47_13;
    _zz_io_MatrixB_47_15 <= _zz_io_MatrixB_47_14;
    _zz_io_MatrixB_47_16 <= _zz_io_MatrixB_47_15;
    _zz_io_MatrixB_47_17 <= _zz_io_MatrixB_47_16;
    _zz_io_MatrixB_47_18 <= _zz_io_MatrixB_47_17;
    _zz_io_MatrixB_47_19 <= _zz_io_MatrixB_47_18;
    _zz_io_MatrixB_47_20 <= _zz_io_MatrixB_47_19;
    _zz_io_MatrixB_47_21 <= _zz_io_MatrixB_47_20;
    _zz_io_MatrixB_47_22 <= _zz_io_MatrixB_47_21;
    _zz_io_MatrixB_47_23 <= _zz_io_MatrixB_47_22;
    _zz_io_MatrixB_47_24 <= _zz_io_MatrixB_47_23;
    _zz_io_MatrixB_47_25 <= _zz_io_MatrixB_47_24;
    _zz_io_MatrixB_47_26 <= _zz_io_MatrixB_47_25;
    _zz_io_MatrixB_47_27 <= _zz_io_MatrixB_47_26;
    _zz_io_MatrixB_47_28 <= _zz_io_MatrixB_47_27;
    _zz_io_MatrixB_47_29 <= _zz_io_MatrixB_47_28;
    _zz_io_MatrixB_47_30 <= _zz_io_MatrixB_47_29;
    _zz_io_MatrixB_47_31 <= _zz_io_MatrixB_47_30;
    _zz_io_MatrixB_47_32 <= _zz_io_MatrixB_47_31;
    _zz_io_MatrixB_47_33 <= _zz_io_MatrixB_47_32;
    _zz_io_MatrixB_47_34 <= _zz_io_MatrixB_47_33;
    _zz_io_MatrixB_47_35 <= _zz_io_MatrixB_47_34;
    _zz_io_MatrixB_47_36 <= _zz_io_MatrixB_47_35;
    _zz_io_MatrixB_47_37 <= _zz_io_MatrixB_47_36;
    _zz_io_MatrixB_47_38 <= _zz_io_MatrixB_47_37;
    _zz_io_MatrixB_47_39 <= _zz_io_MatrixB_47_38;
    _zz_io_MatrixB_47_40 <= _zz_io_MatrixB_47_39;
    _zz_io_MatrixB_47_41 <= _zz_io_MatrixB_47_40;
    _zz_io_MatrixB_47_42 <= _zz_io_MatrixB_47_41;
    _zz_io_MatrixB_47_43 <= _zz_io_MatrixB_47_42;
    _zz_io_MatrixB_47_44 <= _zz_io_MatrixB_47_43;
    _zz_io_MatrixB_47_45 <= _zz_io_MatrixB_47_44;
    _zz_io_MatrixB_47_46 <= _zz_io_MatrixB_47_45;
    _zz_io_B_Valid_47 <= SubModule_WeightCache_MatrixCol_Switch[47];
    _zz_io_B_Valid_47_1 <= _zz_io_B_Valid_47;
    _zz_io_B_Valid_47_2 <= _zz_io_B_Valid_47_1;
    _zz_io_B_Valid_47_3 <= _zz_io_B_Valid_47_2;
    _zz_io_B_Valid_47_4 <= _zz_io_B_Valid_47_3;
    _zz_io_B_Valid_47_5 <= _zz_io_B_Valid_47_4;
    _zz_io_B_Valid_47_6 <= _zz_io_B_Valid_47_5;
    _zz_io_B_Valid_47_7 <= _zz_io_B_Valid_47_6;
    _zz_io_B_Valid_47_8 <= _zz_io_B_Valid_47_7;
    _zz_io_B_Valid_47_9 <= _zz_io_B_Valid_47_8;
    _zz_io_B_Valid_47_10 <= _zz_io_B_Valid_47_9;
    _zz_io_B_Valid_47_11 <= _zz_io_B_Valid_47_10;
    _zz_io_B_Valid_47_12 <= _zz_io_B_Valid_47_11;
    _zz_io_B_Valid_47_13 <= _zz_io_B_Valid_47_12;
    _zz_io_B_Valid_47_14 <= _zz_io_B_Valid_47_13;
    _zz_io_B_Valid_47_15 <= _zz_io_B_Valid_47_14;
    _zz_io_B_Valid_47_16 <= _zz_io_B_Valid_47_15;
    _zz_io_B_Valid_47_17 <= _zz_io_B_Valid_47_16;
    _zz_io_B_Valid_47_18 <= _zz_io_B_Valid_47_17;
    _zz_io_B_Valid_47_19 <= _zz_io_B_Valid_47_18;
    _zz_io_B_Valid_47_20 <= _zz_io_B_Valid_47_19;
    _zz_io_B_Valid_47_21 <= _zz_io_B_Valid_47_20;
    _zz_io_B_Valid_47_22 <= _zz_io_B_Valid_47_21;
    _zz_io_B_Valid_47_23 <= _zz_io_B_Valid_47_22;
    _zz_io_B_Valid_47_24 <= _zz_io_B_Valid_47_23;
    _zz_io_B_Valid_47_25 <= _zz_io_B_Valid_47_24;
    _zz_io_B_Valid_47_26 <= _zz_io_B_Valid_47_25;
    _zz_io_B_Valid_47_27 <= _zz_io_B_Valid_47_26;
    _zz_io_B_Valid_47_28 <= _zz_io_B_Valid_47_27;
    _zz_io_B_Valid_47_29 <= _zz_io_B_Valid_47_28;
    _zz_io_B_Valid_47_30 <= _zz_io_B_Valid_47_29;
    _zz_io_B_Valid_47_31 <= _zz_io_B_Valid_47_30;
    _zz_io_B_Valid_47_32 <= _zz_io_B_Valid_47_31;
    _zz_io_B_Valid_47_33 <= _zz_io_B_Valid_47_32;
    _zz_io_B_Valid_47_34 <= _zz_io_B_Valid_47_33;
    _zz_io_B_Valid_47_35 <= _zz_io_B_Valid_47_34;
    _zz_io_B_Valid_47_36 <= _zz_io_B_Valid_47_35;
    _zz_io_B_Valid_47_37 <= _zz_io_B_Valid_47_36;
    _zz_io_B_Valid_47_38 <= _zz_io_B_Valid_47_37;
    _zz_io_B_Valid_47_39 <= _zz_io_B_Valid_47_38;
    _zz_io_B_Valid_47_40 <= _zz_io_B_Valid_47_39;
    _zz_io_B_Valid_47_41 <= _zz_io_B_Valid_47_40;
    _zz_io_B_Valid_47_42 <= _zz_io_B_Valid_47_41;
    _zz_io_B_Valid_47_43 <= _zz_io_B_Valid_47_42;
    _zz_io_B_Valid_47_44 <= _zz_io_B_Valid_47_43;
    _zz_io_B_Valid_47_45 <= _zz_io_B_Valid_47_44;
    _zz_io_B_Valid_47_46 <= _zz_io_B_Valid_47_45;
    _zz_io_MatrixB_48 <= SubModule_WeightCache_mData_48;
    _zz_io_MatrixB_48_1 <= _zz_io_MatrixB_48;
    _zz_io_MatrixB_48_2 <= _zz_io_MatrixB_48_1;
    _zz_io_MatrixB_48_3 <= _zz_io_MatrixB_48_2;
    _zz_io_MatrixB_48_4 <= _zz_io_MatrixB_48_3;
    _zz_io_MatrixB_48_5 <= _zz_io_MatrixB_48_4;
    _zz_io_MatrixB_48_6 <= _zz_io_MatrixB_48_5;
    _zz_io_MatrixB_48_7 <= _zz_io_MatrixB_48_6;
    _zz_io_MatrixB_48_8 <= _zz_io_MatrixB_48_7;
    _zz_io_MatrixB_48_9 <= _zz_io_MatrixB_48_8;
    _zz_io_MatrixB_48_10 <= _zz_io_MatrixB_48_9;
    _zz_io_MatrixB_48_11 <= _zz_io_MatrixB_48_10;
    _zz_io_MatrixB_48_12 <= _zz_io_MatrixB_48_11;
    _zz_io_MatrixB_48_13 <= _zz_io_MatrixB_48_12;
    _zz_io_MatrixB_48_14 <= _zz_io_MatrixB_48_13;
    _zz_io_MatrixB_48_15 <= _zz_io_MatrixB_48_14;
    _zz_io_MatrixB_48_16 <= _zz_io_MatrixB_48_15;
    _zz_io_MatrixB_48_17 <= _zz_io_MatrixB_48_16;
    _zz_io_MatrixB_48_18 <= _zz_io_MatrixB_48_17;
    _zz_io_MatrixB_48_19 <= _zz_io_MatrixB_48_18;
    _zz_io_MatrixB_48_20 <= _zz_io_MatrixB_48_19;
    _zz_io_MatrixB_48_21 <= _zz_io_MatrixB_48_20;
    _zz_io_MatrixB_48_22 <= _zz_io_MatrixB_48_21;
    _zz_io_MatrixB_48_23 <= _zz_io_MatrixB_48_22;
    _zz_io_MatrixB_48_24 <= _zz_io_MatrixB_48_23;
    _zz_io_MatrixB_48_25 <= _zz_io_MatrixB_48_24;
    _zz_io_MatrixB_48_26 <= _zz_io_MatrixB_48_25;
    _zz_io_MatrixB_48_27 <= _zz_io_MatrixB_48_26;
    _zz_io_MatrixB_48_28 <= _zz_io_MatrixB_48_27;
    _zz_io_MatrixB_48_29 <= _zz_io_MatrixB_48_28;
    _zz_io_MatrixB_48_30 <= _zz_io_MatrixB_48_29;
    _zz_io_MatrixB_48_31 <= _zz_io_MatrixB_48_30;
    _zz_io_MatrixB_48_32 <= _zz_io_MatrixB_48_31;
    _zz_io_MatrixB_48_33 <= _zz_io_MatrixB_48_32;
    _zz_io_MatrixB_48_34 <= _zz_io_MatrixB_48_33;
    _zz_io_MatrixB_48_35 <= _zz_io_MatrixB_48_34;
    _zz_io_MatrixB_48_36 <= _zz_io_MatrixB_48_35;
    _zz_io_MatrixB_48_37 <= _zz_io_MatrixB_48_36;
    _zz_io_MatrixB_48_38 <= _zz_io_MatrixB_48_37;
    _zz_io_MatrixB_48_39 <= _zz_io_MatrixB_48_38;
    _zz_io_MatrixB_48_40 <= _zz_io_MatrixB_48_39;
    _zz_io_MatrixB_48_41 <= _zz_io_MatrixB_48_40;
    _zz_io_MatrixB_48_42 <= _zz_io_MatrixB_48_41;
    _zz_io_MatrixB_48_43 <= _zz_io_MatrixB_48_42;
    _zz_io_MatrixB_48_44 <= _zz_io_MatrixB_48_43;
    _zz_io_MatrixB_48_45 <= _zz_io_MatrixB_48_44;
    _zz_io_MatrixB_48_46 <= _zz_io_MatrixB_48_45;
    _zz_io_MatrixB_48_47 <= _zz_io_MatrixB_48_46;
    _zz_io_B_Valid_48 <= SubModule_WeightCache_MatrixCol_Switch[48];
    _zz_io_B_Valid_48_1 <= _zz_io_B_Valid_48;
    _zz_io_B_Valid_48_2 <= _zz_io_B_Valid_48_1;
    _zz_io_B_Valid_48_3 <= _zz_io_B_Valid_48_2;
    _zz_io_B_Valid_48_4 <= _zz_io_B_Valid_48_3;
    _zz_io_B_Valid_48_5 <= _zz_io_B_Valid_48_4;
    _zz_io_B_Valid_48_6 <= _zz_io_B_Valid_48_5;
    _zz_io_B_Valid_48_7 <= _zz_io_B_Valid_48_6;
    _zz_io_B_Valid_48_8 <= _zz_io_B_Valid_48_7;
    _zz_io_B_Valid_48_9 <= _zz_io_B_Valid_48_8;
    _zz_io_B_Valid_48_10 <= _zz_io_B_Valid_48_9;
    _zz_io_B_Valid_48_11 <= _zz_io_B_Valid_48_10;
    _zz_io_B_Valid_48_12 <= _zz_io_B_Valid_48_11;
    _zz_io_B_Valid_48_13 <= _zz_io_B_Valid_48_12;
    _zz_io_B_Valid_48_14 <= _zz_io_B_Valid_48_13;
    _zz_io_B_Valid_48_15 <= _zz_io_B_Valid_48_14;
    _zz_io_B_Valid_48_16 <= _zz_io_B_Valid_48_15;
    _zz_io_B_Valid_48_17 <= _zz_io_B_Valid_48_16;
    _zz_io_B_Valid_48_18 <= _zz_io_B_Valid_48_17;
    _zz_io_B_Valid_48_19 <= _zz_io_B_Valid_48_18;
    _zz_io_B_Valid_48_20 <= _zz_io_B_Valid_48_19;
    _zz_io_B_Valid_48_21 <= _zz_io_B_Valid_48_20;
    _zz_io_B_Valid_48_22 <= _zz_io_B_Valid_48_21;
    _zz_io_B_Valid_48_23 <= _zz_io_B_Valid_48_22;
    _zz_io_B_Valid_48_24 <= _zz_io_B_Valid_48_23;
    _zz_io_B_Valid_48_25 <= _zz_io_B_Valid_48_24;
    _zz_io_B_Valid_48_26 <= _zz_io_B_Valid_48_25;
    _zz_io_B_Valid_48_27 <= _zz_io_B_Valid_48_26;
    _zz_io_B_Valid_48_28 <= _zz_io_B_Valid_48_27;
    _zz_io_B_Valid_48_29 <= _zz_io_B_Valid_48_28;
    _zz_io_B_Valid_48_30 <= _zz_io_B_Valid_48_29;
    _zz_io_B_Valid_48_31 <= _zz_io_B_Valid_48_30;
    _zz_io_B_Valid_48_32 <= _zz_io_B_Valid_48_31;
    _zz_io_B_Valid_48_33 <= _zz_io_B_Valid_48_32;
    _zz_io_B_Valid_48_34 <= _zz_io_B_Valid_48_33;
    _zz_io_B_Valid_48_35 <= _zz_io_B_Valid_48_34;
    _zz_io_B_Valid_48_36 <= _zz_io_B_Valid_48_35;
    _zz_io_B_Valid_48_37 <= _zz_io_B_Valid_48_36;
    _zz_io_B_Valid_48_38 <= _zz_io_B_Valid_48_37;
    _zz_io_B_Valid_48_39 <= _zz_io_B_Valid_48_38;
    _zz_io_B_Valid_48_40 <= _zz_io_B_Valid_48_39;
    _zz_io_B_Valid_48_41 <= _zz_io_B_Valid_48_40;
    _zz_io_B_Valid_48_42 <= _zz_io_B_Valid_48_41;
    _zz_io_B_Valid_48_43 <= _zz_io_B_Valid_48_42;
    _zz_io_B_Valid_48_44 <= _zz_io_B_Valid_48_43;
    _zz_io_B_Valid_48_45 <= _zz_io_B_Valid_48_44;
    _zz_io_B_Valid_48_46 <= _zz_io_B_Valid_48_45;
    _zz_io_B_Valid_48_47 <= _zz_io_B_Valid_48_46;
    _zz_io_MatrixB_49 <= SubModule_WeightCache_mData_49;
    _zz_io_MatrixB_49_1 <= _zz_io_MatrixB_49;
    _zz_io_MatrixB_49_2 <= _zz_io_MatrixB_49_1;
    _zz_io_MatrixB_49_3 <= _zz_io_MatrixB_49_2;
    _zz_io_MatrixB_49_4 <= _zz_io_MatrixB_49_3;
    _zz_io_MatrixB_49_5 <= _zz_io_MatrixB_49_4;
    _zz_io_MatrixB_49_6 <= _zz_io_MatrixB_49_5;
    _zz_io_MatrixB_49_7 <= _zz_io_MatrixB_49_6;
    _zz_io_MatrixB_49_8 <= _zz_io_MatrixB_49_7;
    _zz_io_MatrixB_49_9 <= _zz_io_MatrixB_49_8;
    _zz_io_MatrixB_49_10 <= _zz_io_MatrixB_49_9;
    _zz_io_MatrixB_49_11 <= _zz_io_MatrixB_49_10;
    _zz_io_MatrixB_49_12 <= _zz_io_MatrixB_49_11;
    _zz_io_MatrixB_49_13 <= _zz_io_MatrixB_49_12;
    _zz_io_MatrixB_49_14 <= _zz_io_MatrixB_49_13;
    _zz_io_MatrixB_49_15 <= _zz_io_MatrixB_49_14;
    _zz_io_MatrixB_49_16 <= _zz_io_MatrixB_49_15;
    _zz_io_MatrixB_49_17 <= _zz_io_MatrixB_49_16;
    _zz_io_MatrixB_49_18 <= _zz_io_MatrixB_49_17;
    _zz_io_MatrixB_49_19 <= _zz_io_MatrixB_49_18;
    _zz_io_MatrixB_49_20 <= _zz_io_MatrixB_49_19;
    _zz_io_MatrixB_49_21 <= _zz_io_MatrixB_49_20;
    _zz_io_MatrixB_49_22 <= _zz_io_MatrixB_49_21;
    _zz_io_MatrixB_49_23 <= _zz_io_MatrixB_49_22;
    _zz_io_MatrixB_49_24 <= _zz_io_MatrixB_49_23;
    _zz_io_MatrixB_49_25 <= _zz_io_MatrixB_49_24;
    _zz_io_MatrixB_49_26 <= _zz_io_MatrixB_49_25;
    _zz_io_MatrixB_49_27 <= _zz_io_MatrixB_49_26;
    _zz_io_MatrixB_49_28 <= _zz_io_MatrixB_49_27;
    _zz_io_MatrixB_49_29 <= _zz_io_MatrixB_49_28;
    _zz_io_MatrixB_49_30 <= _zz_io_MatrixB_49_29;
    _zz_io_MatrixB_49_31 <= _zz_io_MatrixB_49_30;
    _zz_io_MatrixB_49_32 <= _zz_io_MatrixB_49_31;
    _zz_io_MatrixB_49_33 <= _zz_io_MatrixB_49_32;
    _zz_io_MatrixB_49_34 <= _zz_io_MatrixB_49_33;
    _zz_io_MatrixB_49_35 <= _zz_io_MatrixB_49_34;
    _zz_io_MatrixB_49_36 <= _zz_io_MatrixB_49_35;
    _zz_io_MatrixB_49_37 <= _zz_io_MatrixB_49_36;
    _zz_io_MatrixB_49_38 <= _zz_io_MatrixB_49_37;
    _zz_io_MatrixB_49_39 <= _zz_io_MatrixB_49_38;
    _zz_io_MatrixB_49_40 <= _zz_io_MatrixB_49_39;
    _zz_io_MatrixB_49_41 <= _zz_io_MatrixB_49_40;
    _zz_io_MatrixB_49_42 <= _zz_io_MatrixB_49_41;
    _zz_io_MatrixB_49_43 <= _zz_io_MatrixB_49_42;
    _zz_io_MatrixB_49_44 <= _zz_io_MatrixB_49_43;
    _zz_io_MatrixB_49_45 <= _zz_io_MatrixB_49_44;
    _zz_io_MatrixB_49_46 <= _zz_io_MatrixB_49_45;
    _zz_io_MatrixB_49_47 <= _zz_io_MatrixB_49_46;
    _zz_io_MatrixB_49_48 <= _zz_io_MatrixB_49_47;
    _zz_io_B_Valid_49 <= SubModule_WeightCache_MatrixCol_Switch[49];
    _zz_io_B_Valid_49_1 <= _zz_io_B_Valid_49;
    _zz_io_B_Valid_49_2 <= _zz_io_B_Valid_49_1;
    _zz_io_B_Valid_49_3 <= _zz_io_B_Valid_49_2;
    _zz_io_B_Valid_49_4 <= _zz_io_B_Valid_49_3;
    _zz_io_B_Valid_49_5 <= _zz_io_B_Valid_49_4;
    _zz_io_B_Valid_49_6 <= _zz_io_B_Valid_49_5;
    _zz_io_B_Valid_49_7 <= _zz_io_B_Valid_49_6;
    _zz_io_B_Valid_49_8 <= _zz_io_B_Valid_49_7;
    _zz_io_B_Valid_49_9 <= _zz_io_B_Valid_49_8;
    _zz_io_B_Valid_49_10 <= _zz_io_B_Valid_49_9;
    _zz_io_B_Valid_49_11 <= _zz_io_B_Valid_49_10;
    _zz_io_B_Valid_49_12 <= _zz_io_B_Valid_49_11;
    _zz_io_B_Valid_49_13 <= _zz_io_B_Valid_49_12;
    _zz_io_B_Valid_49_14 <= _zz_io_B_Valid_49_13;
    _zz_io_B_Valid_49_15 <= _zz_io_B_Valid_49_14;
    _zz_io_B_Valid_49_16 <= _zz_io_B_Valid_49_15;
    _zz_io_B_Valid_49_17 <= _zz_io_B_Valid_49_16;
    _zz_io_B_Valid_49_18 <= _zz_io_B_Valid_49_17;
    _zz_io_B_Valid_49_19 <= _zz_io_B_Valid_49_18;
    _zz_io_B_Valid_49_20 <= _zz_io_B_Valid_49_19;
    _zz_io_B_Valid_49_21 <= _zz_io_B_Valid_49_20;
    _zz_io_B_Valid_49_22 <= _zz_io_B_Valid_49_21;
    _zz_io_B_Valid_49_23 <= _zz_io_B_Valid_49_22;
    _zz_io_B_Valid_49_24 <= _zz_io_B_Valid_49_23;
    _zz_io_B_Valid_49_25 <= _zz_io_B_Valid_49_24;
    _zz_io_B_Valid_49_26 <= _zz_io_B_Valid_49_25;
    _zz_io_B_Valid_49_27 <= _zz_io_B_Valid_49_26;
    _zz_io_B_Valid_49_28 <= _zz_io_B_Valid_49_27;
    _zz_io_B_Valid_49_29 <= _zz_io_B_Valid_49_28;
    _zz_io_B_Valid_49_30 <= _zz_io_B_Valid_49_29;
    _zz_io_B_Valid_49_31 <= _zz_io_B_Valid_49_30;
    _zz_io_B_Valid_49_32 <= _zz_io_B_Valid_49_31;
    _zz_io_B_Valid_49_33 <= _zz_io_B_Valid_49_32;
    _zz_io_B_Valid_49_34 <= _zz_io_B_Valid_49_33;
    _zz_io_B_Valid_49_35 <= _zz_io_B_Valid_49_34;
    _zz_io_B_Valid_49_36 <= _zz_io_B_Valid_49_35;
    _zz_io_B_Valid_49_37 <= _zz_io_B_Valid_49_36;
    _zz_io_B_Valid_49_38 <= _zz_io_B_Valid_49_37;
    _zz_io_B_Valid_49_39 <= _zz_io_B_Valid_49_38;
    _zz_io_B_Valid_49_40 <= _zz_io_B_Valid_49_39;
    _zz_io_B_Valid_49_41 <= _zz_io_B_Valid_49_40;
    _zz_io_B_Valid_49_42 <= _zz_io_B_Valid_49_41;
    _zz_io_B_Valid_49_43 <= _zz_io_B_Valid_49_42;
    _zz_io_B_Valid_49_44 <= _zz_io_B_Valid_49_43;
    _zz_io_B_Valid_49_45 <= _zz_io_B_Valid_49_44;
    _zz_io_B_Valid_49_46 <= _zz_io_B_Valid_49_45;
    _zz_io_B_Valid_49_47 <= _zz_io_B_Valid_49_46;
    _zz_io_B_Valid_49_48 <= _zz_io_B_Valid_49_47;
    _zz_io_MatrixB_50 <= SubModule_WeightCache_mData_50;
    _zz_io_MatrixB_50_1 <= _zz_io_MatrixB_50;
    _zz_io_MatrixB_50_2 <= _zz_io_MatrixB_50_1;
    _zz_io_MatrixB_50_3 <= _zz_io_MatrixB_50_2;
    _zz_io_MatrixB_50_4 <= _zz_io_MatrixB_50_3;
    _zz_io_MatrixB_50_5 <= _zz_io_MatrixB_50_4;
    _zz_io_MatrixB_50_6 <= _zz_io_MatrixB_50_5;
    _zz_io_MatrixB_50_7 <= _zz_io_MatrixB_50_6;
    _zz_io_MatrixB_50_8 <= _zz_io_MatrixB_50_7;
    _zz_io_MatrixB_50_9 <= _zz_io_MatrixB_50_8;
    _zz_io_MatrixB_50_10 <= _zz_io_MatrixB_50_9;
    _zz_io_MatrixB_50_11 <= _zz_io_MatrixB_50_10;
    _zz_io_MatrixB_50_12 <= _zz_io_MatrixB_50_11;
    _zz_io_MatrixB_50_13 <= _zz_io_MatrixB_50_12;
    _zz_io_MatrixB_50_14 <= _zz_io_MatrixB_50_13;
    _zz_io_MatrixB_50_15 <= _zz_io_MatrixB_50_14;
    _zz_io_MatrixB_50_16 <= _zz_io_MatrixB_50_15;
    _zz_io_MatrixB_50_17 <= _zz_io_MatrixB_50_16;
    _zz_io_MatrixB_50_18 <= _zz_io_MatrixB_50_17;
    _zz_io_MatrixB_50_19 <= _zz_io_MatrixB_50_18;
    _zz_io_MatrixB_50_20 <= _zz_io_MatrixB_50_19;
    _zz_io_MatrixB_50_21 <= _zz_io_MatrixB_50_20;
    _zz_io_MatrixB_50_22 <= _zz_io_MatrixB_50_21;
    _zz_io_MatrixB_50_23 <= _zz_io_MatrixB_50_22;
    _zz_io_MatrixB_50_24 <= _zz_io_MatrixB_50_23;
    _zz_io_MatrixB_50_25 <= _zz_io_MatrixB_50_24;
    _zz_io_MatrixB_50_26 <= _zz_io_MatrixB_50_25;
    _zz_io_MatrixB_50_27 <= _zz_io_MatrixB_50_26;
    _zz_io_MatrixB_50_28 <= _zz_io_MatrixB_50_27;
    _zz_io_MatrixB_50_29 <= _zz_io_MatrixB_50_28;
    _zz_io_MatrixB_50_30 <= _zz_io_MatrixB_50_29;
    _zz_io_MatrixB_50_31 <= _zz_io_MatrixB_50_30;
    _zz_io_MatrixB_50_32 <= _zz_io_MatrixB_50_31;
    _zz_io_MatrixB_50_33 <= _zz_io_MatrixB_50_32;
    _zz_io_MatrixB_50_34 <= _zz_io_MatrixB_50_33;
    _zz_io_MatrixB_50_35 <= _zz_io_MatrixB_50_34;
    _zz_io_MatrixB_50_36 <= _zz_io_MatrixB_50_35;
    _zz_io_MatrixB_50_37 <= _zz_io_MatrixB_50_36;
    _zz_io_MatrixB_50_38 <= _zz_io_MatrixB_50_37;
    _zz_io_MatrixB_50_39 <= _zz_io_MatrixB_50_38;
    _zz_io_MatrixB_50_40 <= _zz_io_MatrixB_50_39;
    _zz_io_MatrixB_50_41 <= _zz_io_MatrixB_50_40;
    _zz_io_MatrixB_50_42 <= _zz_io_MatrixB_50_41;
    _zz_io_MatrixB_50_43 <= _zz_io_MatrixB_50_42;
    _zz_io_MatrixB_50_44 <= _zz_io_MatrixB_50_43;
    _zz_io_MatrixB_50_45 <= _zz_io_MatrixB_50_44;
    _zz_io_MatrixB_50_46 <= _zz_io_MatrixB_50_45;
    _zz_io_MatrixB_50_47 <= _zz_io_MatrixB_50_46;
    _zz_io_MatrixB_50_48 <= _zz_io_MatrixB_50_47;
    _zz_io_MatrixB_50_49 <= _zz_io_MatrixB_50_48;
    _zz_io_B_Valid_50 <= SubModule_WeightCache_MatrixCol_Switch[50];
    _zz_io_B_Valid_50_1 <= _zz_io_B_Valid_50;
    _zz_io_B_Valid_50_2 <= _zz_io_B_Valid_50_1;
    _zz_io_B_Valid_50_3 <= _zz_io_B_Valid_50_2;
    _zz_io_B_Valid_50_4 <= _zz_io_B_Valid_50_3;
    _zz_io_B_Valid_50_5 <= _zz_io_B_Valid_50_4;
    _zz_io_B_Valid_50_6 <= _zz_io_B_Valid_50_5;
    _zz_io_B_Valid_50_7 <= _zz_io_B_Valid_50_6;
    _zz_io_B_Valid_50_8 <= _zz_io_B_Valid_50_7;
    _zz_io_B_Valid_50_9 <= _zz_io_B_Valid_50_8;
    _zz_io_B_Valid_50_10 <= _zz_io_B_Valid_50_9;
    _zz_io_B_Valid_50_11 <= _zz_io_B_Valid_50_10;
    _zz_io_B_Valid_50_12 <= _zz_io_B_Valid_50_11;
    _zz_io_B_Valid_50_13 <= _zz_io_B_Valid_50_12;
    _zz_io_B_Valid_50_14 <= _zz_io_B_Valid_50_13;
    _zz_io_B_Valid_50_15 <= _zz_io_B_Valid_50_14;
    _zz_io_B_Valid_50_16 <= _zz_io_B_Valid_50_15;
    _zz_io_B_Valid_50_17 <= _zz_io_B_Valid_50_16;
    _zz_io_B_Valid_50_18 <= _zz_io_B_Valid_50_17;
    _zz_io_B_Valid_50_19 <= _zz_io_B_Valid_50_18;
    _zz_io_B_Valid_50_20 <= _zz_io_B_Valid_50_19;
    _zz_io_B_Valid_50_21 <= _zz_io_B_Valid_50_20;
    _zz_io_B_Valid_50_22 <= _zz_io_B_Valid_50_21;
    _zz_io_B_Valid_50_23 <= _zz_io_B_Valid_50_22;
    _zz_io_B_Valid_50_24 <= _zz_io_B_Valid_50_23;
    _zz_io_B_Valid_50_25 <= _zz_io_B_Valid_50_24;
    _zz_io_B_Valid_50_26 <= _zz_io_B_Valid_50_25;
    _zz_io_B_Valid_50_27 <= _zz_io_B_Valid_50_26;
    _zz_io_B_Valid_50_28 <= _zz_io_B_Valid_50_27;
    _zz_io_B_Valid_50_29 <= _zz_io_B_Valid_50_28;
    _zz_io_B_Valid_50_30 <= _zz_io_B_Valid_50_29;
    _zz_io_B_Valid_50_31 <= _zz_io_B_Valid_50_30;
    _zz_io_B_Valid_50_32 <= _zz_io_B_Valid_50_31;
    _zz_io_B_Valid_50_33 <= _zz_io_B_Valid_50_32;
    _zz_io_B_Valid_50_34 <= _zz_io_B_Valid_50_33;
    _zz_io_B_Valid_50_35 <= _zz_io_B_Valid_50_34;
    _zz_io_B_Valid_50_36 <= _zz_io_B_Valid_50_35;
    _zz_io_B_Valid_50_37 <= _zz_io_B_Valid_50_36;
    _zz_io_B_Valid_50_38 <= _zz_io_B_Valid_50_37;
    _zz_io_B_Valid_50_39 <= _zz_io_B_Valid_50_38;
    _zz_io_B_Valid_50_40 <= _zz_io_B_Valid_50_39;
    _zz_io_B_Valid_50_41 <= _zz_io_B_Valid_50_40;
    _zz_io_B_Valid_50_42 <= _zz_io_B_Valid_50_41;
    _zz_io_B_Valid_50_43 <= _zz_io_B_Valid_50_42;
    _zz_io_B_Valid_50_44 <= _zz_io_B_Valid_50_43;
    _zz_io_B_Valid_50_45 <= _zz_io_B_Valid_50_44;
    _zz_io_B_Valid_50_46 <= _zz_io_B_Valid_50_45;
    _zz_io_B_Valid_50_47 <= _zz_io_B_Valid_50_46;
    _zz_io_B_Valid_50_48 <= _zz_io_B_Valid_50_47;
    _zz_io_B_Valid_50_49 <= _zz_io_B_Valid_50_48;
    _zz_io_MatrixB_51 <= SubModule_WeightCache_mData_51;
    _zz_io_MatrixB_51_1 <= _zz_io_MatrixB_51;
    _zz_io_MatrixB_51_2 <= _zz_io_MatrixB_51_1;
    _zz_io_MatrixB_51_3 <= _zz_io_MatrixB_51_2;
    _zz_io_MatrixB_51_4 <= _zz_io_MatrixB_51_3;
    _zz_io_MatrixB_51_5 <= _zz_io_MatrixB_51_4;
    _zz_io_MatrixB_51_6 <= _zz_io_MatrixB_51_5;
    _zz_io_MatrixB_51_7 <= _zz_io_MatrixB_51_6;
    _zz_io_MatrixB_51_8 <= _zz_io_MatrixB_51_7;
    _zz_io_MatrixB_51_9 <= _zz_io_MatrixB_51_8;
    _zz_io_MatrixB_51_10 <= _zz_io_MatrixB_51_9;
    _zz_io_MatrixB_51_11 <= _zz_io_MatrixB_51_10;
    _zz_io_MatrixB_51_12 <= _zz_io_MatrixB_51_11;
    _zz_io_MatrixB_51_13 <= _zz_io_MatrixB_51_12;
    _zz_io_MatrixB_51_14 <= _zz_io_MatrixB_51_13;
    _zz_io_MatrixB_51_15 <= _zz_io_MatrixB_51_14;
    _zz_io_MatrixB_51_16 <= _zz_io_MatrixB_51_15;
    _zz_io_MatrixB_51_17 <= _zz_io_MatrixB_51_16;
    _zz_io_MatrixB_51_18 <= _zz_io_MatrixB_51_17;
    _zz_io_MatrixB_51_19 <= _zz_io_MatrixB_51_18;
    _zz_io_MatrixB_51_20 <= _zz_io_MatrixB_51_19;
    _zz_io_MatrixB_51_21 <= _zz_io_MatrixB_51_20;
    _zz_io_MatrixB_51_22 <= _zz_io_MatrixB_51_21;
    _zz_io_MatrixB_51_23 <= _zz_io_MatrixB_51_22;
    _zz_io_MatrixB_51_24 <= _zz_io_MatrixB_51_23;
    _zz_io_MatrixB_51_25 <= _zz_io_MatrixB_51_24;
    _zz_io_MatrixB_51_26 <= _zz_io_MatrixB_51_25;
    _zz_io_MatrixB_51_27 <= _zz_io_MatrixB_51_26;
    _zz_io_MatrixB_51_28 <= _zz_io_MatrixB_51_27;
    _zz_io_MatrixB_51_29 <= _zz_io_MatrixB_51_28;
    _zz_io_MatrixB_51_30 <= _zz_io_MatrixB_51_29;
    _zz_io_MatrixB_51_31 <= _zz_io_MatrixB_51_30;
    _zz_io_MatrixB_51_32 <= _zz_io_MatrixB_51_31;
    _zz_io_MatrixB_51_33 <= _zz_io_MatrixB_51_32;
    _zz_io_MatrixB_51_34 <= _zz_io_MatrixB_51_33;
    _zz_io_MatrixB_51_35 <= _zz_io_MatrixB_51_34;
    _zz_io_MatrixB_51_36 <= _zz_io_MatrixB_51_35;
    _zz_io_MatrixB_51_37 <= _zz_io_MatrixB_51_36;
    _zz_io_MatrixB_51_38 <= _zz_io_MatrixB_51_37;
    _zz_io_MatrixB_51_39 <= _zz_io_MatrixB_51_38;
    _zz_io_MatrixB_51_40 <= _zz_io_MatrixB_51_39;
    _zz_io_MatrixB_51_41 <= _zz_io_MatrixB_51_40;
    _zz_io_MatrixB_51_42 <= _zz_io_MatrixB_51_41;
    _zz_io_MatrixB_51_43 <= _zz_io_MatrixB_51_42;
    _zz_io_MatrixB_51_44 <= _zz_io_MatrixB_51_43;
    _zz_io_MatrixB_51_45 <= _zz_io_MatrixB_51_44;
    _zz_io_MatrixB_51_46 <= _zz_io_MatrixB_51_45;
    _zz_io_MatrixB_51_47 <= _zz_io_MatrixB_51_46;
    _zz_io_MatrixB_51_48 <= _zz_io_MatrixB_51_47;
    _zz_io_MatrixB_51_49 <= _zz_io_MatrixB_51_48;
    _zz_io_MatrixB_51_50 <= _zz_io_MatrixB_51_49;
    _zz_io_B_Valid_51 <= SubModule_WeightCache_MatrixCol_Switch[51];
    _zz_io_B_Valid_51_1 <= _zz_io_B_Valid_51;
    _zz_io_B_Valid_51_2 <= _zz_io_B_Valid_51_1;
    _zz_io_B_Valid_51_3 <= _zz_io_B_Valid_51_2;
    _zz_io_B_Valid_51_4 <= _zz_io_B_Valid_51_3;
    _zz_io_B_Valid_51_5 <= _zz_io_B_Valid_51_4;
    _zz_io_B_Valid_51_6 <= _zz_io_B_Valid_51_5;
    _zz_io_B_Valid_51_7 <= _zz_io_B_Valid_51_6;
    _zz_io_B_Valid_51_8 <= _zz_io_B_Valid_51_7;
    _zz_io_B_Valid_51_9 <= _zz_io_B_Valid_51_8;
    _zz_io_B_Valid_51_10 <= _zz_io_B_Valid_51_9;
    _zz_io_B_Valid_51_11 <= _zz_io_B_Valid_51_10;
    _zz_io_B_Valid_51_12 <= _zz_io_B_Valid_51_11;
    _zz_io_B_Valid_51_13 <= _zz_io_B_Valid_51_12;
    _zz_io_B_Valid_51_14 <= _zz_io_B_Valid_51_13;
    _zz_io_B_Valid_51_15 <= _zz_io_B_Valid_51_14;
    _zz_io_B_Valid_51_16 <= _zz_io_B_Valid_51_15;
    _zz_io_B_Valid_51_17 <= _zz_io_B_Valid_51_16;
    _zz_io_B_Valid_51_18 <= _zz_io_B_Valid_51_17;
    _zz_io_B_Valid_51_19 <= _zz_io_B_Valid_51_18;
    _zz_io_B_Valid_51_20 <= _zz_io_B_Valid_51_19;
    _zz_io_B_Valid_51_21 <= _zz_io_B_Valid_51_20;
    _zz_io_B_Valid_51_22 <= _zz_io_B_Valid_51_21;
    _zz_io_B_Valid_51_23 <= _zz_io_B_Valid_51_22;
    _zz_io_B_Valid_51_24 <= _zz_io_B_Valid_51_23;
    _zz_io_B_Valid_51_25 <= _zz_io_B_Valid_51_24;
    _zz_io_B_Valid_51_26 <= _zz_io_B_Valid_51_25;
    _zz_io_B_Valid_51_27 <= _zz_io_B_Valid_51_26;
    _zz_io_B_Valid_51_28 <= _zz_io_B_Valid_51_27;
    _zz_io_B_Valid_51_29 <= _zz_io_B_Valid_51_28;
    _zz_io_B_Valid_51_30 <= _zz_io_B_Valid_51_29;
    _zz_io_B_Valid_51_31 <= _zz_io_B_Valid_51_30;
    _zz_io_B_Valid_51_32 <= _zz_io_B_Valid_51_31;
    _zz_io_B_Valid_51_33 <= _zz_io_B_Valid_51_32;
    _zz_io_B_Valid_51_34 <= _zz_io_B_Valid_51_33;
    _zz_io_B_Valid_51_35 <= _zz_io_B_Valid_51_34;
    _zz_io_B_Valid_51_36 <= _zz_io_B_Valid_51_35;
    _zz_io_B_Valid_51_37 <= _zz_io_B_Valid_51_36;
    _zz_io_B_Valid_51_38 <= _zz_io_B_Valid_51_37;
    _zz_io_B_Valid_51_39 <= _zz_io_B_Valid_51_38;
    _zz_io_B_Valid_51_40 <= _zz_io_B_Valid_51_39;
    _zz_io_B_Valid_51_41 <= _zz_io_B_Valid_51_40;
    _zz_io_B_Valid_51_42 <= _zz_io_B_Valid_51_41;
    _zz_io_B_Valid_51_43 <= _zz_io_B_Valid_51_42;
    _zz_io_B_Valid_51_44 <= _zz_io_B_Valid_51_43;
    _zz_io_B_Valid_51_45 <= _zz_io_B_Valid_51_44;
    _zz_io_B_Valid_51_46 <= _zz_io_B_Valid_51_45;
    _zz_io_B_Valid_51_47 <= _zz_io_B_Valid_51_46;
    _zz_io_B_Valid_51_48 <= _zz_io_B_Valid_51_47;
    _zz_io_B_Valid_51_49 <= _zz_io_B_Valid_51_48;
    _zz_io_B_Valid_51_50 <= _zz_io_B_Valid_51_49;
    _zz_io_MatrixB_52 <= SubModule_WeightCache_mData_52;
    _zz_io_MatrixB_52_1 <= _zz_io_MatrixB_52;
    _zz_io_MatrixB_52_2 <= _zz_io_MatrixB_52_1;
    _zz_io_MatrixB_52_3 <= _zz_io_MatrixB_52_2;
    _zz_io_MatrixB_52_4 <= _zz_io_MatrixB_52_3;
    _zz_io_MatrixB_52_5 <= _zz_io_MatrixB_52_4;
    _zz_io_MatrixB_52_6 <= _zz_io_MatrixB_52_5;
    _zz_io_MatrixB_52_7 <= _zz_io_MatrixB_52_6;
    _zz_io_MatrixB_52_8 <= _zz_io_MatrixB_52_7;
    _zz_io_MatrixB_52_9 <= _zz_io_MatrixB_52_8;
    _zz_io_MatrixB_52_10 <= _zz_io_MatrixB_52_9;
    _zz_io_MatrixB_52_11 <= _zz_io_MatrixB_52_10;
    _zz_io_MatrixB_52_12 <= _zz_io_MatrixB_52_11;
    _zz_io_MatrixB_52_13 <= _zz_io_MatrixB_52_12;
    _zz_io_MatrixB_52_14 <= _zz_io_MatrixB_52_13;
    _zz_io_MatrixB_52_15 <= _zz_io_MatrixB_52_14;
    _zz_io_MatrixB_52_16 <= _zz_io_MatrixB_52_15;
    _zz_io_MatrixB_52_17 <= _zz_io_MatrixB_52_16;
    _zz_io_MatrixB_52_18 <= _zz_io_MatrixB_52_17;
    _zz_io_MatrixB_52_19 <= _zz_io_MatrixB_52_18;
    _zz_io_MatrixB_52_20 <= _zz_io_MatrixB_52_19;
    _zz_io_MatrixB_52_21 <= _zz_io_MatrixB_52_20;
    _zz_io_MatrixB_52_22 <= _zz_io_MatrixB_52_21;
    _zz_io_MatrixB_52_23 <= _zz_io_MatrixB_52_22;
    _zz_io_MatrixB_52_24 <= _zz_io_MatrixB_52_23;
    _zz_io_MatrixB_52_25 <= _zz_io_MatrixB_52_24;
    _zz_io_MatrixB_52_26 <= _zz_io_MatrixB_52_25;
    _zz_io_MatrixB_52_27 <= _zz_io_MatrixB_52_26;
    _zz_io_MatrixB_52_28 <= _zz_io_MatrixB_52_27;
    _zz_io_MatrixB_52_29 <= _zz_io_MatrixB_52_28;
    _zz_io_MatrixB_52_30 <= _zz_io_MatrixB_52_29;
    _zz_io_MatrixB_52_31 <= _zz_io_MatrixB_52_30;
    _zz_io_MatrixB_52_32 <= _zz_io_MatrixB_52_31;
    _zz_io_MatrixB_52_33 <= _zz_io_MatrixB_52_32;
    _zz_io_MatrixB_52_34 <= _zz_io_MatrixB_52_33;
    _zz_io_MatrixB_52_35 <= _zz_io_MatrixB_52_34;
    _zz_io_MatrixB_52_36 <= _zz_io_MatrixB_52_35;
    _zz_io_MatrixB_52_37 <= _zz_io_MatrixB_52_36;
    _zz_io_MatrixB_52_38 <= _zz_io_MatrixB_52_37;
    _zz_io_MatrixB_52_39 <= _zz_io_MatrixB_52_38;
    _zz_io_MatrixB_52_40 <= _zz_io_MatrixB_52_39;
    _zz_io_MatrixB_52_41 <= _zz_io_MatrixB_52_40;
    _zz_io_MatrixB_52_42 <= _zz_io_MatrixB_52_41;
    _zz_io_MatrixB_52_43 <= _zz_io_MatrixB_52_42;
    _zz_io_MatrixB_52_44 <= _zz_io_MatrixB_52_43;
    _zz_io_MatrixB_52_45 <= _zz_io_MatrixB_52_44;
    _zz_io_MatrixB_52_46 <= _zz_io_MatrixB_52_45;
    _zz_io_MatrixB_52_47 <= _zz_io_MatrixB_52_46;
    _zz_io_MatrixB_52_48 <= _zz_io_MatrixB_52_47;
    _zz_io_MatrixB_52_49 <= _zz_io_MatrixB_52_48;
    _zz_io_MatrixB_52_50 <= _zz_io_MatrixB_52_49;
    _zz_io_MatrixB_52_51 <= _zz_io_MatrixB_52_50;
    _zz_io_B_Valid_52 <= SubModule_WeightCache_MatrixCol_Switch[52];
    _zz_io_B_Valid_52_1 <= _zz_io_B_Valid_52;
    _zz_io_B_Valid_52_2 <= _zz_io_B_Valid_52_1;
    _zz_io_B_Valid_52_3 <= _zz_io_B_Valid_52_2;
    _zz_io_B_Valid_52_4 <= _zz_io_B_Valid_52_3;
    _zz_io_B_Valid_52_5 <= _zz_io_B_Valid_52_4;
    _zz_io_B_Valid_52_6 <= _zz_io_B_Valid_52_5;
    _zz_io_B_Valid_52_7 <= _zz_io_B_Valid_52_6;
    _zz_io_B_Valid_52_8 <= _zz_io_B_Valid_52_7;
    _zz_io_B_Valid_52_9 <= _zz_io_B_Valid_52_8;
    _zz_io_B_Valid_52_10 <= _zz_io_B_Valid_52_9;
    _zz_io_B_Valid_52_11 <= _zz_io_B_Valid_52_10;
    _zz_io_B_Valid_52_12 <= _zz_io_B_Valid_52_11;
    _zz_io_B_Valid_52_13 <= _zz_io_B_Valid_52_12;
    _zz_io_B_Valid_52_14 <= _zz_io_B_Valid_52_13;
    _zz_io_B_Valid_52_15 <= _zz_io_B_Valid_52_14;
    _zz_io_B_Valid_52_16 <= _zz_io_B_Valid_52_15;
    _zz_io_B_Valid_52_17 <= _zz_io_B_Valid_52_16;
    _zz_io_B_Valid_52_18 <= _zz_io_B_Valid_52_17;
    _zz_io_B_Valid_52_19 <= _zz_io_B_Valid_52_18;
    _zz_io_B_Valid_52_20 <= _zz_io_B_Valid_52_19;
    _zz_io_B_Valid_52_21 <= _zz_io_B_Valid_52_20;
    _zz_io_B_Valid_52_22 <= _zz_io_B_Valid_52_21;
    _zz_io_B_Valid_52_23 <= _zz_io_B_Valid_52_22;
    _zz_io_B_Valid_52_24 <= _zz_io_B_Valid_52_23;
    _zz_io_B_Valid_52_25 <= _zz_io_B_Valid_52_24;
    _zz_io_B_Valid_52_26 <= _zz_io_B_Valid_52_25;
    _zz_io_B_Valid_52_27 <= _zz_io_B_Valid_52_26;
    _zz_io_B_Valid_52_28 <= _zz_io_B_Valid_52_27;
    _zz_io_B_Valid_52_29 <= _zz_io_B_Valid_52_28;
    _zz_io_B_Valid_52_30 <= _zz_io_B_Valid_52_29;
    _zz_io_B_Valid_52_31 <= _zz_io_B_Valid_52_30;
    _zz_io_B_Valid_52_32 <= _zz_io_B_Valid_52_31;
    _zz_io_B_Valid_52_33 <= _zz_io_B_Valid_52_32;
    _zz_io_B_Valid_52_34 <= _zz_io_B_Valid_52_33;
    _zz_io_B_Valid_52_35 <= _zz_io_B_Valid_52_34;
    _zz_io_B_Valid_52_36 <= _zz_io_B_Valid_52_35;
    _zz_io_B_Valid_52_37 <= _zz_io_B_Valid_52_36;
    _zz_io_B_Valid_52_38 <= _zz_io_B_Valid_52_37;
    _zz_io_B_Valid_52_39 <= _zz_io_B_Valid_52_38;
    _zz_io_B_Valid_52_40 <= _zz_io_B_Valid_52_39;
    _zz_io_B_Valid_52_41 <= _zz_io_B_Valid_52_40;
    _zz_io_B_Valid_52_42 <= _zz_io_B_Valid_52_41;
    _zz_io_B_Valid_52_43 <= _zz_io_B_Valid_52_42;
    _zz_io_B_Valid_52_44 <= _zz_io_B_Valid_52_43;
    _zz_io_B_Valid_52_45 <= _zz_io_B_Valid_52_44;
    _zz_io_B_Valid_52_46 <= _zz_io_B_Valid_52_45;
    _zz_io_B_Valid_52_47 <= _zz_io_B_Valid_52_46;
    _zz_io_B_Valid_52_48 <= _zz_io_B_Valid_52_47;
    _zz_io_B_Valid_52_49 <= _zz_io_B_Valid_52_48;
    _zz_io_B_Valid_52_50 <= _zz_io_B_Valid_52_49;
    _zz_io_B_Valid_52_51 <= _zz_io_B_Valid_52_50;
    _zz_io_MatrixB_53 <= SubModule_WeightCache_mData_53;
    _zz_io_MatrixB_53_1 <= _zz_io_MatrixB_53;
    _zz_io_MatrixB_53_2 <= _zz_io_MatrixB_53_1;
    _zz_io_MatrixB_53_3 <= _zz_io_MatrixB_53_2;
    _zz_io_MatrixB_53_4 <= _zz_io_MatrixB_53_3;
    _zz_io_MatrixB_53_5 <= _zz_io_MatrixB_53_4;
    _zz_io_MatrixB_53_6 <= _zz_io_MatrixB_53_5;
    _zz_io_MatrixB_53_7 <= _zz_io_MatrixB_53_6;
    _zz_io_MatrixB_53_8 <= _zz_io_MatrixB_53_7;
    _zz_io_MatrixB_53_9 <= _zz_io_MatrixB_53_8;
    _zz_io_MatrixB_53_10 <= _zz_io_MatrixB_53_9;
    _zz_io_MatrixB_53_11 <= _zz_io_MatrixB_53_10;
    _zz_io_MatrixB_53_12 <= _zz_io_MatrixB_53_11;
    _zz_io_MatrixB_53_13 <= _zz_io_MatrixB_53_12;
    _zz_io_MatrixB_53_14 <= _zz_io_MatrixB_53_13;
    _zz_io_MatrixB_53_15 <= _zz_io_MatrixB_53_14;
    _zz_io_MatrixB_53_16 <= _zz_io_MatrixB_53_15;
    _zz_io_MatrixB_53_17 <= _zz_io_MatrixB_53_16;
    _zz_io_MatrixB_53_18 <= _zz_io_MatrixB_53_17;
    _zz_io_MatrixB_53_19 <= _zz_io_MatrixB_53_18;
    _zz_io_MatrixB_53_20 <= _zz_io_MatrixB_53_19;
    _zz_io_MatrixB_53_21 <= _zz_io_MatrixB_53_20;
    _zz_io_MatrixB_53_22 <= _zz_io_MatrixB_53_21;
    _zz_io_MatrixB_53_23 <= _zz_io_MatrixB_53_22;
    _zz_io_MatrixB_53_24 <= _zz_io_MatrixB_53_23;
    _zz_io_MatrixB_53_25 <= _zz_io_MatrixB_53_24;
    _zz_io_MatrixB_53_26 <= _zz_io_MatrixB_53_25;
    _zz_io_MatrixB_53_27 <= _zz_io_MatrixB_53_26;
    _zz_io_MatrixB_53_28 <= _zz_io_MatrixB_53_27;
    _zz_io_MatrixB_53_29 <= _zz_io_MatrixB_53_28;
    _zz_io_MatrixB_53_30 <= _zz_io_MatrixB_53_29;
    _zz_io_MatrixB_53_31 <= _zz_io_MatrixB_53_30;
    _zz_io_MatrixB_53_32 <= _zz_io_MatrixB_53_31;
    _zz_io_MatrixB_53_33 <= _zz_io_MatrixB_53_32;
    _zz_io_MatrixB_53_34 <= _zz_io_MatrixB_53_33;
    _zz_io_MatrixB_53_35 <= _zz_io_MatrixB_53_34;
    _zz_io_MatrixB_53_36 <= _zz_io_MatrixB_53_35;
    _zz_io_MatrixB_53_37 <= _zz_io_MatrixB_53_36;
    _zz_io_MatrixB_53_38 <= _zz_io_MatrixB_53_37;
    _zz_io_MatrixB_53_39 <= _zz_io_MatrixB_53_38;
    _zz_io_MatrixB_53_40 <= _zz_io_MatrixB_53_39;
    _zz_io_MatrixB_53_41 <= _zz_io_MatrixB_53_40;
    _zz_io_MatrixB_53_42 <= _zz_io_MatrixB_53_41;
    _zz_io_MatrixB_53_43 <= _zz_io_MatrixB_53_42;
    _zz_io_MatrixB_53_44 <= _zz_io_MatrixB_53_43;
    _zz_io_MatrixB_53_45 <= _zz_io_MatrixB_53_44;
    _zz_io_MatrixB_53_46 <= _zz_io_MatrixB_53_45;
    _zz_io_MatrixB_53_47 <= _zz_io_MatrixB_53_46;
    _zz_io_MatrixB_53_48 <= _zz_io_MatrixB_53_47;
    _zz_io_MatrixB_53_49 <= _zz_io_MatrixB_53_48;
    _zz_io_MatrixB_53_50 <= _zz_io_MatrixB_53_49;
    _zz_io_MatrixB_53_51 <= _zz_io_MatrixB_53_50;
    _zz_io_MatrixB_53_52 <= _zz_io_MatrixB_53_51;
    _zz_io_B_Valid_53 <= SubModule_WeightCache_MatrixCol_Switch[53];
    _zz_io_B_Valid_53_1 <= _zz_io_B_Valid_53;
    _zz_io_B_Valid_53_2 <= _zz_io_B_Valid_53_1;
    _zz_io_B_Valid_53_3 <= _zz_io_B_Valid_53_2;
    _zz_io_B_Valid_53_4 <= _zz_io_B_Valid_53_3;
    _zz_io_B_Valid_53_5 <= _zz_io_B_Valid_53_4;
    _zz_io_B_Valid_53_6 <= _zz_io_B_Valid_53_5;
    _zz_io_B_Valid_53_7 <= _zz_io_B_Valid_53_6;
    _zz_io_B_Valid_53_8 <= _zz_io_B_Valid_53_7;
    _zz_io_B_Valid_53_9 <= _zz_io_B_Valid_53_8;
    _zz_io_B_Valid_53_10 <= _zz_io_B_Valid_53_9;
    _zz_io_B_Valid_53_11 <= _zz_io_B_Valid_53_10;
    _zz_io_B_Valid_53_12 <= _zz_io_B_Valid_53_11;
    _zz_io_B_Valid_53_13 <= _zz_io_B_Valid_53_12;
    _zz_io_B_Valid_53_14 <= _zz_io_B_Valid_53_13;
    _zz_io_B_Valid_53_15 <= _zz_io_B_Valid_53_14;
    _zz_io_B_Valid_53_16 <= _zz_io_B_Valid_53_15;
    _zz_io_B_Valid_53_17 <= _zz_io_B_Valid_53_16;
    _zz_io_B_Valid_53_18 <= _zz_io_B_Valid_53_17;
    _zz_io_B_Valid_53_19 <= _zz_io_B_Valid_53_18;
    _zz_io_B_Valid_53_20 <= _zz_io_B_Valid_53_19;
    _zz_io_B_Valid_53_21 <= _zz_io_B_Valid_53_20;
    _zz_io_B_Valid_53_22 <= _zz_io_B_Valid_53_21;
    _zz_io_B_Valid_53_23 <= _zz_io_B_Valid_53_22;
    _zz_io_B_Valid_53_24 <= _zz_io_B_Valid_53_23;
    _zz_io_B_Valid_53_25 <= _zz_io_B_Valid_53_24;
    _zz_io_B_Valid_53_26 <= _zz_io_B_Valid_53_25;
    _zz_io_B_Valid_53_27 <= _zz_io_B_Valid_53_26;
    _zz_io_B_Valid_53_28 <= _zz_io_B_Valid_53_27;
    _zz_io_B_Valid_53_29 <= _zz_io_B_Valid_53_28;
    _zz_io_B_Valid_53_30 <= _zz_io_B_Valid_53_29;
    _zz_io_B_Valid_53_31 <= _zz_io_B_Valid_53_30;
    _zz_io_B_Valid_53_32 <= _zz_io_B_Valid_53_31;
    _zz_io_B_Valid_53_33 <= _zz_io_B_Valid_53_32;
    _zz_io_B_Valid_53_34 <= _zz_io_B_Valid_53_33;
    _zz_io_B_Valid_53_35 <= _zz_io_B_Valid_53_34;
    _zz_io_B_Valid_53_36 <= _zz_io_B_Valid_53_35;
    _zz_io_B_Valid_53_37 <= _zz_io_B_Valid_53_36;
    _zz_io_B_Valid_53_38 <= _zz_io_B_Valid_53_37;
    _zz_io_B_Valid_53_39 <= _zz_io_B_Valid_53_38;
    _zz_io_B_Valid_53_40 <= _zz_io_B_Valid_53_39;
    _zz_io_B_Valid_53_41 <= _zz_io_B_Valid_53_40;
    _zz_io_B_Valid_53_42 <= _zz_io_B_Valid_53_41;
    _zz_io_B_Valid_53_43 <= _zz_io_B_Valid_53_42;
    _zz_io_B_Valid_53_44 <= _zz_io_B_Valid_53_43;
    _zz_io_B_Valid_53_45 <= _zz_io_B_Valid_53_44;
    _zz_io_B_Valid_53_46 <= _zz_io_B_Valid_53_45;
    _zz_io_B_Valid_53_47 <= _zz_io_B_Valid_53_46;
    _zz_io_B_Valid_53_48 <= _zz_io_B_Valid_53_47;
    _zz_io_B_Valid_53_49 <= _zz_io_B_Valid_53_48;
    _zz_io_B_Valid_53_50 <= _zz_io_B_Valid_53_49;
    _zz_io_B_Valid_53_51 <= _zz_io_B_Valid_53_50;
    _zz_io_B_Valid_53_52 <= _zz_io_B_Valid_53_51;
    _zz_io_MatrixB_54 <= SubModule_WeightCache_mData_54;
    _zz_io_MatrixB_54_1 <= _zz_io_MatrixB_54;
    _zz_io_MatrixB_54_2 <= _zz_io_MatrixB_54_1;
    _zz_io_MatrixB_54_3 <= _zz_io_MatrixB_54_2;
    _zz_io_MatrixB_54_4 <= _zz_io_MatrixB_54_3;
    _zz_io_MatrixB_54_5 <= _zz_io_MatrixB_54_4;
    _zz_io_MatrixB_54_6 <= _zz_io_MatrixB_54_5;
    _zz_io_MatrixB_54_7 <= _zz_io_MatrixB_54_6;
    _zz_io_MatrixB_54_8 <= _zz_io_MatrixB_54_7;
    _zz_io_MatrixB_54_9 <= _zz_io_MatrixB_54_8;
    _zz_io_MatrixB_54_10 <= _zz_io_MatrixB_54_9;
    _zz_io_MatrixB_54_11 <= _zz_io_MatrixB_54_10;
    _zz_io_MatrixB_54_12 <= _zz_io_MatrixB_54_11;
    _zz_io_MatrixB_54_13 <= _zz_io_MatrixB_54_12;
    _zz_io_MatrixB_54_14 <= _zz_io_MatrixB_54_13;
    _zz_io_MatrixB_54_15 <= _zz_io_MatrixB_54_14;
    _zz_io_MatrixB_54_16 <= _zz_io_MatrixB_54_15;
    _zz_io_MatrixB_54_17 <= _zz_io_MatrixB_54_16;
    _zz_io_MatrixB_54_18 <= _zz_io_MatrixB_54_17;
    _zz_io_MatrixB_54_19 <= _zz_io_MatrixB_54_18;
    _zz_io_MatrixB_54_20 <= _zz_io_MatrixB_54_19;
    _zz_io_MatrixB_54_21 <= _zz_io_MatrixB_54_20;
    _zz_io_MatrixB_54_22 <= _zz_io_MatrixB_54_21;
    _zz_io_MatrixB_54_23 <= _zz_io_MatrixB_54_22;
    _zz_io_MatrixB_54_24 <= _zz_io_MatrixB_54_23;
    _zz_io_MatrixB_54_25 <= _zz_io_MatrixB_54_24;
    _zz_io_MatrixB_54_26 <= _zz_io_MatrixB_54_25;
    _zz_io_MatrixB_54_27 <= _zz_io_MatrixB_54_26;
    _zz_io_MatrixB_54_28 <= _zz_io_MatrixB_54_27;
    _zz_io_MatrixB_54_29 <= _zz_io_MatrixB_54_28;
    _zz_io_MatrixB_54_30 <= _zz_io_MatrixB_54_29;
    _zz_io_MatrixB_54_31 <= _zz_io_MatrixB_54_30;
    _zz_io_MatrixB_54_32 <= _zz_io_MatrixB_54_31;
    _zz_io_MatrixB_54_33 <= _zz_io_MatrixB_54_32;
    _zz_io_MatrixB_54_34 <= _zz_io_MatrixB_54_33;
    _zz_io_MatrixB_54_35 <= _zz_io_MatrixB_54_34;
    _zz_io_MatrixB_54_36 <= _zz_io_MatrixB_54_35;
    _zz_io_MatrixB_54_37 <= _zz_io_MatrixB_54_36;
    _zz_io_MatrixB_54_38 <= _zz_io_MatrixB_54_37;
    _zz_io_MatrixB_54_39 <= _zz_io_MatrixB_54_38;
    _zz_io_MatrixB_54_40 <= _zz_io_MatrixB_54_39;
    _zz_io_MatrixB_54_41 <= _zz_io_MatrixB_54_40;
    _zz_io_MatrixB_54_42 <= _zz_io_MatrixB_54_41;
    _zz_io_MatrixB_54_43 <= _zz_io_MatrixB_54_42;
    _zz_io_MatrixB_54_44 <= _zz_io_MatrixB_54_43;
    _zz_io_MatrixB_54_45 <= _zz_io_MatrixB_54_44;
    _zz_io_MatrixB_54_46 <= _zz_io_MatrixB_54_45;
    _zz_io_MatrixB_54_47 <= _zz_io_MatrixB_54_46;
    _zz_io_MatrixB_54_48 <= _zz_io_MatrixB_54_47;
    _zz_io_MatrixB_54_49 <= _zz_io_MatrixB_54_48;
    _zz_io_MatrixB_54_50 <= _zz_io_MatrixB_54_49;
    _zz_io_MatrixB_54_51 <= _zz_io_MatrixB_54_50;
    _zz_io_MatrixB_54_52 <= _zz_io_MatrixB_54_51;
    _zz_io_MatrixB_54_53 <= _zz_io_MatrixB_54_52;
    _zz_io_B_Valid_54 <= SubModule_WeightCache_MatrixCol_Switch[54];
    _zz_io_B_Valid_54_1 <= _zz_io_B_Valid_54;
    _zz_io_B_Valid_54_2 <= _zz_io_B_Valid_54_1;
    _zz_io_B_Valid_54_3 <= _zz_io_B_Valid_54_2;
    _zz_io_B_Valid_54_4 <= _zz_io_B_Valid_54_3;
    _zz_io_B_Valid_54_5 <= _zz_io_B_Valid_54_4;
    _zz_io_B_Valid_54_6 <= _zz_io_B_Valid_54_5;
    _zz_io_B_Valid_54_7 <= _zz_io_B_Valid_54_6;
    _zz_io_B_Valid_54_8 <= _zz_io_B_Valid_54_7;
    _zz_io_B_Valid_54_9 <= _zz_io_B_Valid_54_8;
    _zz_io_B_Valid_54_10 <= _zz_io_B_Valid_54_9;
    _zz_io_B_Valid_54_11 <= _zz_io_B_Valid_54_10;
    _zz_io_B_Valid_54_12 <= _zz_io_B_Valid_54_11;
    _zz_io_B_Valid_54_13 <= _zz_io_B_Valid_54_12;
    _zz_io_B_Valid_54_14 <= _zz_io_B_Valid_54_13;
    _zz_io_B_Valid_54_15 <= _zz_io_B_Valid_54_14;
    _zz_io_B_Valid_54_16 <= _zz_io_B_Valid_54_15;
    _zz_io_B_Valid_54_17 <= _zz_io_B_Valid_54_16;
    _zz_io_B_Valid_54_18 <= _zz_io_B_Valid_54_17;
    _zz_io_B_Valid_54_19 <= _zz_io_B_Valid_54_18;
    _zz_io_B_Valid_54_20 <= _zz_io_B_Valid_54_19;
    _zz_io_B_Valid_54_21 <= _zz_io_B_Valid_54_20;
    _zz_io_B_Valid_54_22 <= _zz_io_B_Valid_54_21;
    _zz_io_B_Valid_54_23 <= _zz_io_B_Valid_54_22;
    _zz_io_B_Valid_54_24 <= _zz_io_B_Valid_54_23;
    _zz_io_B_Valid_54_25 <= _zz_io_B_Valid_54_24;
    _zz_io_B_Valid_54_26 <= _zz_io_B_Valid_54_25;
    _zz_io_B_Valid_54_27 <= _zz_io_B_Valid_54_26;
    _zz_io_B_Valid_54_28 <= _zz_io_B_Valid_54_27;
    _zz_io_B_Valid_54_29 <= _zz_io_B_Valid_54_28;
    _zz_io_B_Valid_54_30 <= _zz_io_B_Valid_54_29;
    _zz_io_B_Valid_54_31 <= _zz_io_B_Valid_54_30;
    _zz_io_B_Valid_54_32 <= _zz_io_B_Valid_54_31;
    _zz_io_B_Valid_54_33 <= _zz_io_B_Valid_54_32;
    _zz_io_B_Valid_54_34 <= _zz_io_B_Valid_54_33;
    _zz_io_B_Valid_54_35 <= _zz_io_B_Valid_54_34;
    _zz_io_B_Valid_54_36 <= _zz_io_B_Valid_54_35;
    _zz_io_B_Valid_54_37 <= _zz_io_B_Valid_54_36;
    _zz_io_B_Valid_54_38 <= _zz_io_B_Valid_54_37;
    _zz_io_B_Valid_54_39 <= _zz_io_B_Valid_54_38;
    _zz_io_B_Valid_54_40 <= _zz_io_B_Valid_54_39;
    _zz_io_B_Valid_54_41 <= _zz_io_B_Valid_54_40;
    _zz_io_B_Valid_54_42 <= _zz_io_B_Valid_54_41;
    _zz_io_B_Valid_54_43 <= _zz_io_B_Valid_54_42;
    _zz_io_B_Valid_54_44 <= _zz_io_B_Valid_54_43;
    _zz_io_B_Valid_54_45 <= _zz_io_B_Valid_54_44;
    _zz_io_B_Valid_54_46 <= _zz_io_B_Valid_54_45;
    _zz_io_B_Valid_54_47 <= _zz_io_B_Valid_54_46;
    _zz_io_B_Valid_54_48 <= _zz_io_B_Valid_54_47;
    _zz_io_B_Valid_54_49 <= _zz_io_B_Valid_54_48;
    _zz_io_B_Valid_54_50 <= _zz_io_B_Valid_54_49;
    _zz_io_B_Valid_54_51 <= _zz_io_B_Valid_54_50;
    _zz_io_B_Valid_54_52 <= _zz_io_B_Valid_54_51;
    _zz_io_B_Valid_54_53 <= _zz_io_B_Valid_54_52;
    _zz_io_MatrixB_55 <= SubModule_WeightCache_mData_55;
    _zz_io_MatrixB_55_1 <= _zz_io_MatrixB_55;
    _zz_io_MatrixB_55_2 <= _zz_io_MatrixB_55_1;
    _zz_io_MatrixB_55_3 <= _zz_io_MatrixB_55_2;
    _zz_io_MatrixB_55_4 <= _zz_io_MatrixB_55_3;
    _zz_io_MatrixB_55_5 <= _zz_io_MatrixB_55_4;
    _zz_io_MatrixB_55_6 <= _zz_io_MatrixB_55_5;
    _zz_io_MatrixB_55_7 <= _zz_io_MatrixB_55_6;
    _zz_io_MatrixB_55_8 <= _zz_io_MatrixB_55_7;
    _zz_io_MatrixB_55_9 <= _zz_io_MatrixB_55_8;
    _zz_io_MatrixB_55_10 <= _zz_io_MatrixB_55_9;
    _zz_io_MatrixB_55_11 <= _zz_io_MatrixB_55_10;
    _zz_io_MatrixB_55_12 <= _zz_io_MatrixB_55_11;
    _zz_io_MatrixB_55_13 <= _zz_io_MatrixB_55_12;
    _zz_io_MatrixB_55_14 <= _zz_io_MatrixB_55_13;
    _zz_io_MatrixB_55_15 <= _zz_io_MatrixB_55_14;
    _zz_io_MatrixB_55_16 <= _zz_io_MatrixB_55_15;
    _zz_io_MatrixB_55_17 <= _zz_io_MatrixB_55_16;
    _zz_io_MatrixB_55_18 <= _zz_io_MatrixB_55_17;
    _zz_io_MatrixB_55_19 <= _zz_io_MatrixB_55_18;
    _zz_io_MatrixB_55_20 <= _zz_io_MatrixB_55_19;
    _zz_io_MatrixB_55_21 <= _zz_io_MatrixB_55_20;
    _zz_io_MatrixB_55_22 <= _zz_io_MatrixB_55_21;
    _zz_io_MatrixB_55_23 <= _zz_io_MatrixB_55_22;
    _zz_io_MatrixB_55_24 <= _zz_io_MatrixB_55_23;
    _zz_io_MatrixB_55_25 <= _zz_io_MatrixB_55_24;
    _zz_io_MatrixB_55_26 <= _zz_io_MatrixB_55_25;
    _zz_io_MatrixB_55_27 <= _zz_io_MatrixB_55_26;
    _zz_io_MatrixB_55_28 <= _zz_io_MatrixB_55_27;
    _zz_io_MatrixB_55_29 <= _zz_io_MatrixB_55_28;
    _zz_io_MatrixB_55_30 <= _zz_io_MatrixB_55_29;
    _zz_io_MatrixB_55_31 <= _zz_io_MatrixB_55_30;
    _zz_io_MatrixB_55_32 <= _zz_io_MatrixB_55_31;
    _zz_io_MatrixB_55_33 <= _zz_io_MatrixB_55_32;
    _zz_io_MatrixB_55_34 <= _zz_io_MatrixB_55_33;
    _zz_io_MatrixB_55_35 <= _zz_io_MatrixB_55_34;
    _zz_io_MatrixB_55_36 <= _zz_io_MatrixB_55_35;
    _zz_io_MatrixB_55_37 <= _zz_io_MatrixB_55_36;
    _zz_io_MatrixB_55_38 <= _zz_io_MatrixB_55_37;
    _zz_io_MatrixB_55_39 <= _zz_io_MatrixB_55_38;
    _zz_io_MatrixB_55_40 <= _zz_io_MatrixB_55_39;
    _zz_io_MatrixB_55_41 <= _zz_io_MatrixB_55_40;
    _zz_io_MatrixB_55_42 <= _zz_io_MatrixB_55_41;
    _zz_io_MatrixB_55_43 <= _zz_io_MatrixB_55_42;
    _zz_io_MatrixB_55_44 <= _zz_io_MatrixB_55_43;
    _zz_io_MatrixB_55_45 <= _zz_io_MatrixB_55_44;
    _zz_io_MatrixB_55_46 <= _zz_io_MatrixB_55_45;
    _zz_io_MatrixB_55_47 <= _zz_io_MatrixB_55_46;
    _zz_io_MatrixB_55_48 <= _zz_io_MatrixB_55_47;
    _zz_io_MatrixB_55_49 <= _zz_io_MatrixB_55_48;
    _zz_io_MatrixB_55_50 <= _zz_io_MatrixB_55_49;
    _zz_io_MatrixB_55_51 <= _zz_io_MatrixB_55_50;
    _zz_io_MatrixB_55_52 <= _zz_io_MatrixB_55_51;
    _zz_io_MatrixB_55_53 <= _zz_io_MatrixB_55_52;
    _zz_io_MatrixB_55_54 <= _zz_io_MatrixB_55_53;
    _zz_io_B_Valid_55 <= SubModule_WeightCache_MatrixCol_Switch[55];
    _zz_io_B_Valid_55_1 <= _zz_io_B_Valid_55;
    _zz_io_B_Valid_55_2 <= _zz_io_B_Valid_55_1;
    _zz_io_B_Valid_55_3 <= _zz_io_B_Valid_55_2;
    _zz_io_B_Valid_55_4 <= _zz_io_B_Valid_55_3;
    _zz_io_B_Valid_55_5 <= _zz_io_B_Valid_55_4;
    _zz_io_B_Valid_55_6 <= _zz_io_B_Valid_55_5;
    _zz_io_B_Valid_55_7 <= _zz_io_B_Valid_55_6;
    _zz_io_B_Valid_55_8 <= _zz_io_B_Valid_55_7;
    _zz_io_B_Valid_55_9 <= _zz_io_B_Valid_55_8;
    _zz_io_B_Valid_55_10 <= _zz_io_B_Valid_55_9;
    _zz_io_B_Valid_55_11 <= _zz_io_B_Valid_55_10;
    _zz_io_B_Valid_55_12 <= _zz_io_B_Valid_55_11;
    _zz_io_B_Valid_55_13 <= _zz_io_B_Valid_55_12;
    _zz_io_B_Valid_55_14 <= _zz_io_B_Valid_55_13;
    _zz_io_B_Valid_55_15 <= _zz_io_B_Valid_55_14;
    _zz_io_B_Valid_55_16 <= _zz_io_B_Valid_55_15;
    _zz_io_B_Valid_55_17 <= _zz_io_B_Valid_55_16;
    _zz_io_B_Valid_55_18 <= _zz_io_B_Valid_55_17;
    _zz_io_B_Valid_55_19 <= _zz_io_B_Valid_55_18;
    _zz_io_B_Valid_55_20 <= _zz_io_B_Valid_55_19;
    _zz_io_B_Valid_55_21 <= _zz_io_B_Valid_55_20;
    _zz_io_B_Valid_55_22 <= _zz_io_B_Valid_55_21;
    _zz_io_B_Valid_55_23 <= _zz_io_B_Valid_55_22;
    _zz_io_B_Valid_55_24 <= _zz_io_B_Valid_55_23;
    _zz_io_B_Valid_55_25 <= _zz_io_B_Valid_55_24;
    _zz_io_B_Valid_55_26 <= _zz_io_B_Valid_55_25;
    _zz_io_B_Valid_55_27 <= _zz_io_B_Valid_55_26;
    _zz_io_B_Valid_55_28 <= _zz_io_B_Valid_55_27;
    _zz_io_B_Valid_55_29 <= _zz_io_B_Valid_55_28;
    _zz_io_B_Valid_55_30 <= _zz_io_B_Valid_55_29;
    _zz_io_B_Valid_55_31 <= _zz_io_B_Valid_55_30;
    _zz_io_B_Valid_55_32 <= _zz_io_B_Valid_55_31;
    _zz_io_B_Valid_55_33 <= _zz_io_B_Valid_55_32;
    _zz_io_B_Valid_55_34 <= _zz_io_B_Valid_55_33;
    _zz_io_B_Valid_55_35 <= _zz_io_B_Valid_55_34;
    _zz_io_B_Valid_55_36 <= _zz_io_B_Valid_55_35;
    _zz_io_B_Valid_55_37 <= _zz_io_B_Valid_55_36;
    _zz_io_B_Valid_55_38 <= _zz_io_B_Valid_55_37;
    _zz_io_B_Valid_55_39 <= _zz_io_B_Valid_55_38;
    _zz_io_B_Valid_55_40 <= _zz_io_B_Valid_55_39;
    _zz_io_B_Valid_55_41 <= _zz_io_B_Valid_55_40;
    _zz_io_B_Valid_55_42 <= _zz_io_B_Valid_55_41;
    _zz_io_B_Valid_55_43 <= _zz_io_B_Valid_55_42;
    _zz_io_B_Valid_55_44 <= _zz_io_B_Valid_55_43;
    _zz_io_B_Valid_55_45 <= _zz_io_B_Valid_55_44;
    _zz_io_B_Valid_55_46 <= _zz_io_B_Valid_55_45;
    _zz_io_B_Valid_55_47 <= _zz_io_B_Valid_55_46;
    _zz_io_B_Valid_55_48 <= _zz_io_B_Valid_55_47;
    _zz_io_B_Valid_55_49 <= _zz_io_B_Valid_55_48;
    _zz_io_B_Valid_55_50 <= _zz_io_B_Valid_55_49;
    _zz_io_B_Valid_55_51 <= _zz_io_B_Valid_55_50;
    _zz_io_B_Valid_55_52 <= _zz_io_B_Valid_55_51;
    _zz_io_B_Valid_55_53 <= _zz_io_B_Valid_55_52;
    _zz_io_B_Valid_55_54 <= _zz_io_B_Valid_55_53;
    _zz_io_MatrixB_56 <= SubModule_WeightCache_mData_56;
    _zz_io_MatrixB_56_1 <= _zz_io_MatrixB_56;
    _zz_io_MatrixB_56_2 <= _zz_io_MatrixB_56_1;
    _zz_io_MatrixB_56_3 <= _zz_io_MatrixB_56_2;
    _zz_io_MatrixB_56_4 <= _zz_io_MatrixB_56_3;
    _zz_io_MatrixB_56_5 <= _zz_io_MatrixB_56_4;
    _zz_io_MatrixB_56_6 <= _zz_io_MatrixB_56_5;
    _zz_io_MatrixB_56_7 <= _zz_io_MatrixB_56_6;
    _zz_io_MatrixB_56_8 <= _zz_io_MatrixB_56_7;
    _zz_io_MatrixB_56_9 <= _zz_io_MatrixB_56_8;
    _zz_io_MatrixB_56_10 <= _zz_io_MatrixB_56_9;
    _zz_io_MatrixB_56_11 <= _zz_io_MatrixB_56_10;
    _zz_io_MatrixB_56_12 <= _zz_io_MatrixB_56_11;
    _zz_io_MatrixB_56_13 <= _zz_io_MatrixB_56_12;
    _zz_io_MatrixB_56_14 <= _zz_io_MatrixB_56_13;
    _zz_io_MatrixB_56_15 <= _zz_io_MatrixB_56_14;
    _zz_io_MatrixB_56_16 <= _zz_io_MatrixB_56_15;
    _zz_io_MatrixB_56_17 <= _zz_io_MatrixB_56_16;
    _zz_io_MatrixB_56_18 <= _zz_io_MatrixB_56_17;
    _zz_io_MatrixB_56_19 <= _zz_io_MatrixB_56_18;
    _zz_io_MatrixB_56_20 <= _zz_io_MatrixB_56_19;
    _zz_io_MatrixB_56_21 <= _zz_io_MatrixB_56_20;
    _zz_io_MatrixB_56_22 <= _zz_io_MatrixB_56_21;
    _zz_io_MatrixB_56_23 <= _zz_io_MatrixB_56_22;
    _zz_io_MatrixB_56_24 <= _zz_io_MatrixB_56_23;
    _zz_io_MatrixB_56_25 <= _zz_io_MatrixB_56_24;
    _zz_io_MatrixB_56_26 <= _zz_io_MatrixB_56_25;
    _zz_io_MatrixB_56_27 <= _zz_io_MatrixB_56_26;
    _zz_io_MatrixB_56_28 <= _zz_io_MatrixB_56_27;
    _zz_io_MatrixB_56_29 <= _zz_io_MatrixB_56_28;
    _zz_io_MatrixB_56_30 <= _zz_io_MatrixB_56_29;
    _zz_io_MatrixB_56_31 <= _zz_io_MatrixB_56_30;
    _zz_io_MatrixB_56_32 <= _zz_io_MatrixB_56_31;
    _zz_io_MatrixB_56_33 <= _zz_io_MatrixB_56_32;
    _zz_io_MatrixB_56_34 <= _zz_io_MatrixB_56_33;
    _zz_io_MatrixB_56_35 <= _zz_io_MatrixB_56_34;
    _zz_io_MatrixB_56_36 <= _zz_io_MatrixB_56_35;
    _zz_io_MatrixB_56_37 <= _zz_io_MatrixB_56_36;
    _zz_io_MatrixB_56_38 <= _zz_io_MatrixB_56_37;
    _zz_io_MatrixB_56_39 <= _zz_io_MatrixB_56_38;
    _zz_io_MatrixB_56_40 <= _zz_io_MatrixB_56_39;
    _zz_io_MatrixB_56_41 <= _zz_io_MatrixB_56_40;
    _zz_io_MatrixB_56_42 <= _zz_io_MatrixB_56_41;
    _zz_io_MatrixB_56_43 <= _zz_io_MatrixB_56_42;
    _zz_io_MatrixB_56_44 <= _zz_io_MatrixB_56_43;
    _zz_io_MatrixB_56_45 <= _zz_io_MatrixB_56_44;
    _zz_io_MatrixB_56_46 <= _zz_io_MatrixB_56_45;
    _zz_io_MatrixB_56_47 <= _zz_io_MatrixB_56_46;
    _zz_io_MatrixB_56_48 <= _zz_io_MatrixB_56_47;
    _zz_io_MatrixB_56_49 <= _zz_io_MatrixB_56_48;
    _zz_io_MatrixB_56_50 <= _zz_io_MatrixB_56_49;
    _zz_io_MatrixB_56_51 <= _zz_io_MatrixB_56_50;
    _zz_io_MatrixB_56_52 <= _zz_io_MatrixB_56_51;
    _zz_io_MatrixB_56_53 <= _zz_io_MatrixB_56_52;
    _zz_io_MatrixB_56_54 <= _zz_io_MatrixB_56_53;
    _zz_io_MatrixB_56_55 <= _zz_io_MatrixB_56_54;
    _zz_io_B_Valid_56 <= SubModule_WeightCache_MatrixCol_Switch[56];
    _zz_io_B_Valid_56_1 <= _zz_io_B_Valid_56;
    _zz_io_B_Valid_56_2 <= _zz_io_B_Valid_56_1;
    _zz_io_B_Valid_56_3 <= _zz_io_B_Valid_56_2;
    _zz_io_B_Valid_56_4 <= _zz_io_B_Valid_56_3;
    _zz_io_B_Valid_56_5 <= _zz_io_B_Valid_56_4;
    _zz_io_B_Valid_56_6 <= _zz_io_B_Valid_56_5;
    _zz_io_B_Valid_56_7 <= _zz_io_B_Valid_56_6;
    _zz_io_B_Valid_56_8 <= _zz_io_B_Valid_56_7;
    _zz_io_B_Valid_56_9 <= _zz_io_B_Valid_56_8;
    _zz_io_B_Valid_56_10 <= _zz_io_B_Valid_56_9;
    _zz_io_B_Valid_56_11 <= _zz_io_B_Valid_56_10;
    _zz_io_B_Valid_56_12 <= _zz_io_B_Valid_56_11;
    _zz_io_B_Valid_56_13 <= _zz_io_B_Valid_56_12;
    _zz_io_B_Valid_56_14 <= _zz_io_B_Valid_56_13;
    _zz_io_B_Valid_56_15 <= _zz_io_B_Valid_56_14;
    _zz_io_B_Valid_56_16 <= _zz_io_B_Valid_56_15;
    _zz_io_B_Valid_56_17 <= _zz_io_B_Valid_56_16;
    _zz_io_B_Valid_56_18 <= _zz_io_B_Valid_56_17;
    _zz_io_B_Valid_56_19 <= _zz_io_B_Valid_56_18;
    _zz_io_B_Valid_56_20 <= _zz_io_B_Valid_56_19;
    _zz_io_B_Valid_56_21 <= _zz_io_B_Valid_56_20;
    _zz_io_B_Valid_56_22 <= _zz_io_B_Valid_56_21;
    _zz_io_B_Valid_56_23 <= _zz_io_B_Valid_56_22;
    _zz_io_B_Valid_56_24 <= _zz_io_B_Valid_56_23;
    _zz_io_B_Valid_56_25 <= _zz_io_B_Valid_56_24;
    _zz_io_B_Valid_56_26 <= _zz_io_B_Valid_56_25;
    _zz_io_B_Valid_56_27 <= _zz_io_B_Valid_56_26;
    _zz_io_B_Valid_56_28 <= _zz_io_B_Valid_56_27;
    _zz_io_B_Valid_56_29 <= _zz_io_B_Valid_56_28;
    _zz_io_B_Valid_56_30 <= _zz_io_B_Valid_56_29;
    _zz_io_B_Valid_56_31 <= _zz_io_B_Valid_56_30;
    _zz_io_B_Valid_56_32 <= _zz_io_B_Valid_56_31;
    _zz_io_B_Valid_56_33 <= _zz_io_B_Valid_56_32;
    _zz_io_B_Valid_56_34 <= _zz_io_B_Valid_56_33;
    _zz_io_B_Valid_56_35 <= _zz_io_B_Valid_56_34;
    _zz_io_B_Valid_56_36 <= _zz_io_B_Valid_56_35;
    _zz_io_B_Valid_56_37 <= _zz_io_B_Valid_56_36;
    _zz_io_B_Valid_56_38 <= _zz_io_B_Valid_56_37;
    _zz_io_B_Valid_56_39 <= _zz_io_B_Valid_56_38;
    _zz_io_B_Valid_56_40 <= _zz_io_B_Valid_56_39;
    _zz_io_B_Valid_56_41 <= _zz_io_B_Valid_56_40;
    _zz_io_B_Valid_56_42 <= _zz_io_B_Valid_56_41;
    _zz_io_B_Valid_56_43 <= _zz_io_B_Valid_56_42;
    _zz_io_B_Valid_56_44 <= _zz_io_B_Valid_56_43;
    _zz_io_B_Valid_56_45 <= _zz_io_B_Valid_56_44;
    _zz_io_B_Valid_56_46 <= _zz_io_B_Valid_56_45;
    _zz_io_B_Valid_56_47 <= _zz_io_B_Valid_56_46;
    _zz_io_B_Valid_56_48 <= _zz_io_B_Valid_56_47;
    _zz_io_B_Valid_56_49 <= _zz_io_B_Valid_56_48;
    _zz_io_B_Valid_56_50 <= _zz_io_B_Valid_56_49;
    _zz_io_B_Valid_56_51 <= _zz_io_B_Valid_56_50;
    _zz_io_B_Valid_56_52 <= _zz_io_B_Valid_56_51;
    _zz_io_B_Valid_56_53 <= _zz_io_B_Valid_56_52;
    _zz_io_B_Valid_56_54 <= _zz_io_B_Valid_56_53;
    _zz_io_B_Valid_56_55 <= _zz_io_B_Valid_56_54;
    _zz_io_MatrixB_57 <= SubModule_WeightCache_mData_57;
    _zz_io_MatrixB_57_1 <= _zz_io_MatrixB_57;
    _zz_io_MatrixB_57_2 <= _zz_io_MatrixB_57_1;
    _zz_io_MatrixB_57_3 <= _zz_io_MatrixB_57_2;
    _zz_io_MatrixB_57_4 <= _zz_io_MatrixB_57_3;
    _zz_io_MatrixB_57_5 <= _zz_io_MatrixB_57_4;
    _zz_io_MatrixB_57_6 <= _zz_io_MatrixB_57_5;
    _zz_io_MatrixB_57_7 <= _zz_io_MatrixB_57_6;
    _zz_io_MatrixB_57_8 <= _zz_io_MatrixB_57_7;
    _zz_io_MatrixB_57_9 <= _zz_io_MatrixB_57_8;
    _zz_io_MatrixB_57_10 <= _zz_io_MatrixB_57_9;
    _zz_io_MatrixB_57_11 <= _zz_io_MatrixB_57_10;
    _zz_io_MatrixB_57_12 <= _zz_io_MatrixB_57_11;
    _zz_io_MatrixB_57_13 <= _zz_io_MatrixB_57_12;
    _zz_io_MatrixB_57_14 <= _zz_io_MatrixB_57_13;
    _zz_io_MatrixB_57_15 <= _zz_io_MatrixB_57_14;
    _zz_io_MatrixB_57_16 <= _zz_io_MatrixB_57_15;
    _zz_io_MatrixB_57_17 <= _zz_io_MatrixB_57_16;
    _zz_io_MatrixB_57_18 <= _zz_io_MatrixB_57_17;
    _zz_io_MatrixB_57_19 <= _zz_io_MatrixB_57_18;
    _zz_io_MatrixB_57_20 <= _zz_io_MatrixB_57_19;
    _zz_io_MatrixB_57_21 <= _zz_io_MatrixB_57_20;
    _zz_io_MatrixB_57_22 <= _zz_io_MatrixB_57_21;
    _zz_io_MatrixB_57_23 <= _zz_io_MatrixB_57_22;
    _zz_io_MatrixB_57_24 <= _zz_io_MatrixB_57_23;
    _zz_io_MatrixB_57_25 <= _zz_io_MatrixB_57_24;
    _zz_io_MatrixB_57_26 <= _zz_io_MatrixB_57_25;
    _zz_io_MatrixB_57_27 <= _zz_io_MatrixB_57_26;
    _zz_io_MatrixB_57_28 <= _zz_io_MatrixB_57_27;
    _zz_io_MatrixB_57_29 <= _zz_io_MatrixB_57_28;
    _zz_io_MatrixB_57_30 <= _zz_io_MatrixB_57_29;
    _zz_io_MatrixB_57_31 <= _zz_io_MatrixB_57_30;
    _zz_io_MatrixB_57_32 <= _zz_io_MatrixB_57_31;
    _zz_io_MatrixB_57_33 <= _zz_io_MatrixB_57_32;
    _zz_io_MatrixB_57_34 <= _zz_io_MatrixB_57_33;
    _zz_io_MatrixB_57_35 <= _zz_io_MatrixB_57_34;
    _zz_io_MatrixB_57_36 <= _zz_io_MatrixB_57_35;
    _zz_io_MatrixB_57_37 <= _zz_io_MatrixB_57_36;
    _zz_io_MatrixB_57_38 <= _zz_io_MatrixB_57_37;
    _zz_io_MatrixB_57_39 <= _zz_io_MatrixB_57_38;
    _zz_io_MatrixB_57_40 <= _zz_io_MatrixB_57_39;
    _zz_io_MatrixB_57_41 <= _zz_io_MatrixB_57_40;
    _zz_io_MatrixB_57_42 <= _zz_io_MatrixB_57_41;
    _zz_io_MatrixB_57_43 <= _zz_io_MatrixB_57_42;
    _zz_io_MatrixB_57_44 <= _zz_io_MatrixB_57_43;
    _zz_io_MatrixB_57_45 <= _zz_io_MatrixB_57_44;
    _zz_io_MatrixB_57_46 <= _zz_io_MatrixB_57_45;
    _zz_io_MatrixB_57_47 <= _zz_io_MatrixB_57_46;
    _zz_io_MatrixB_57_48 <= _zz_io_MatrixB_57_47;
    _zz_io_MatrixB_57_49 <= _zz_io_MatrixB_57_48;
    _zz_io_MatrixB_57_50 <= _zz_io_MatrixB_57_49;
    _zz_io_MatrixB_57_51 <= _zz_io_MatrixB_57_50;
    _zz_io_MatrixB_57_52 <= _zz_io_MatrixB_57_51;
    _zz_io_MatrixB_57_53 <= _zz_io_MatrixB_57_52;
    _zz_io_MatrixB_57_54 <= _zz_io_MatrixB_57_53;
    _zz_io_MatrixB_57_55 <= _zz_io_MatrixB_57_54;
    _zz_io_MatrixB_57_56 <= _zz_io_MatrixB_57_55;
    _zz_io_B_Valid_57 <= SubModule_WeightCache_MatrixCol_Switch[57];
    _zz_io_B_Valid_57_1 <= _zz_io_B_Valid_57;
    _zz_io_B_Valid_57_2 <= _zz_io_B_Valid_57_1;
    _zz_io_B_Valid_57_3 <= _zz_io_B_Valid_57_2;
    _zz_io_B_Valid_57_4 <= _zz_io_B_Valid_57_3;
    _zz_io_B_Valid_57_5 <= _zz_io_B_Valid_57_4;
    _zz_io_B_Valid_57_6 <= _zz_io_B_Valid_57_5;
    _zz_io_B_Valid_57_7 <= _zz_io_B_Valid_57_6;
    _zz_io_B_Valid_57_8 <= _zz_io_B_Valid_57_7;
    _zz_io_B_Valid_57_9 <= _zz_io_B_Valid_57_8;
    _zz_io_B_Valid_57_10 <= _zz_io_B_Valid_57_9;
    _zz_io_B_Valid_57_11 <= _zz_io_B_Valid_57_10;
    _zz_io_B_Valid_57_12 <= _zz_io_B_Valid_57_11;
    _zz_io_B_Valid_57_13 <= _zz_io_B_Valid_57_12;
    _zz_io_B_Valid_57_14 <= _zz_io_B_Valid_57_13;
    _zz_io_B_Valid_57_15 <= _zz_io_B_Valid_57_14;
    _zz_io_B_Valid_57_16 <= _zz_io_B_Valid_57_15;
    _zz_io_B_Valid_57_17 <= _zz_io_B_Valid_57_16;
    _zz_io_B_Valid_57_18 <= _zz_io_B_Valid_57_17;
    _zz_io_B_Valid_57_19 <= _zz_io_B_Valid_57_18;
    _zz_io_B_Valid_57_20 <= _zz_io_B_Valid_57_19;
    _zz_io_B_Valid_57_21 <= _zz_io_B_Valid_57_20;
    _zz_io_B_Valid_57_22 <= _zz_io_B_Valid_57_21;
    _zz_io_B_Valid_57_23 <= _zz_io_B_Valid_57_22;
    _zz_io_B_Valid_57_24 <= _zz_io_B_Valid_57_23;
    _zz_io_B_Valid_57_25 <= _zz_io_B_Valid_57_24;
    _zz_io_B_Valid_57_26 <= _zz_io_B_Valid_57_25;
    _zz_io_B_Valid_57_27 <= _zz_io_B_Valid_57_26;
    _zz_io_B_Valid_57_28 <= _zz_io_B_Valid_57_27;
    _zz_io_B_Valid_57_29 <= _zz_io_B_Valid_57_28;
    _zz_io_B_Valid_57_30 <= _zz_io_B_Valid_57_29;
    _zz_io_B_Valid_57_31 <= _zz_io_B_Valid_57_30;
    _zz_io_B_Valid_57_32 <= _zz_io_B_Valid_57_31;
    _zz_io_B_Valid_57_33 <= _zz_io_B_Valid_57_32;
    _zz_io_B_Valid_57_34 <= _zz_io_B_Valid_57_33;
    _zz_io_B_Valid_57_35 <= _zz_io_B_Valid_57_34;
    _zz_io_B_Valid_57_36 <= _zz_io_B_Valid_57_35;
    _zz_io_B_Valid_57_37 <= _zz_io_B_Valid_57_36;
    _zz_io_B_Valid_57_38 <= _zz_io_B_Valid_57_37;
    _zz_io_B_Valid_57_39 <= _zz_io_B_Valid_57_38;
    _zz_io_B_Valid_57_40 <= _zz_io_B_Valid_57_39;
    _zz_io_B_Valid_57_41 <= _zz_io_B_Valid_57_40;
    _zz_io_B_Valid_57_42 <= _zz_io_B_Valid_57_41;
    _zz_io_B_Valid_57_43 <= _zz_io_B_Valid_57_42;
    _zz_io_B_Valid_57_44 <= _zz_io_B_Valid_57_43;
    _zz_io_B_Valid_57_45 <= _zz_io_B_Valid_57_44;
    _zz_io_B_Valid_57_46 <= _zz_io_B_Valid_57_45;
    _zz_io_B_Valid_57_47 <= _zz_io_B_Valid_57_46;
    _zz_io_B_Valid_57_48 <= _zz_io_B_Valid_57_47;
    _zz_io_B_Valid_57_49 <= _zz_io_B_Valid_57_48;
    _zz_io_B_Valid_57_50 <= _zz_io_B_Valid_57_49;
    _zz_io_B_Valid_57_51 <= _zz_io_B_Valid_57_50;
    _zz_io_B_Valid_57_52 <= _zz_io_B_Valid_57_51;
    _zz_io_B_Valid_57_53 <= _zz_io_B_Valid_57_52;
    _zz_io_B_Valid_57_54 <= _zz_io_B_Valid_57_53;
    _zz_io_B_Valid_57_55 <= _zz_io_B_Valid_57_54;
    _zz_io_B_Valid_57_56 <= _zz_io_B_Valid_57_55;
    _zz_io_MatrixB_58 <= SubModule_WeightCache_mData_58;
    _zz_io_MatrixB_58_1 <= _zz_io_MatrixB_58;
    _zz_io_MatrixB_58_2 <= _zz_io_MatrixB_58_1;
    _zz_io_MatrixB_58_3 <= _zz_io_MatrixB_58_2;
    _zz_io_MatrixB_58_4 <= _zz_io_MatrixB_58_3;
    _zz_io_MatrixB_58_5 <= _zz_io_MatrixB_58_4;
    _zz_io_MatrixB_58_6 <= _zz_io_MatrixB_58_5;
    _zz_io_MatrixB_58_7 <= _zz_io_MatrixB_58_6;
    _zz_io_MatrixB_58_8 <= _zz_io_MatrixB_58_7;
    _zz_io_MatrixB_58_9 <= _zz_io_MatrixB_58_8;
    _zz_io_MatrixB_58_10 <= _zz_io_MatrixB_58_9;
    _zz_io_MatrixB_58_11 <= _zz_io_MatrixB_58_10;
    _zz_io_MatrixB_58_12 <= _zz_io_MatrixB_58_11;
    _zz_io_MatrixB_58_13 <= _zz_io_MatrixB_58_12;
    _zz_io_MatrixB_58_14 <= _zz_io_MatrixB_58_13;
    _zz_io_MatrixB_58_15 <= _zz_io_MatrixB_58_14;
    _zz_io_MatrixB_58_16 <= _zz_io_MatrixB_58_15;
    _zz_io_MatrixB_58_17 <= _zz_io_MatrixB_58_16;
    _zz_io_MatrixB_58_18 <= _zz_io_MatrixB_58_17;
    _zz_io_MatrixB_58_19 <= _zz_io_MatrixB_58_18;
    _zz_io_MatrixB_58_20 <= _zz_io_MatrixB_58_19;
    _zz_io_MatrixB_58_21 <= _zz_io_MatrixB_58_20;
    _zz_io_MatrixB_58_22 <= _zz_io_MatrixB_58_21;
    _zz_io_MatrixB_58_23 <= _zz_io_MatrixB_58_22;
    _zz_io_MatrixB_58_24 <= _zz_io_MatrixB_58_23;
    _zz_io_MatrixB_58_25 <= _zz_io_MatrixB_58_24;
    _zz_io_MatrixB_58_26 <= _zz_io_MatrixB_58_25;
    _zz_io_MatrixB_58_27 <= _zz_io_MatrixB_58_26;
    _zz_io_MatrixB_58_28 <= _zz_io_MatrixB_58_27;
    _zz_io_MatrixB_58_29 <= _zz_io_MatrixB_58_28;
    _zz_io_MatrixB_58_30 <= _zz_io_MatrixB_58_29;
    _zz_io_MatrixB_58_31 <= _zz_io_MatrixB_58_30;
    _zz_io_MatrixB_58_32 <= _zz_io_MatrixB_58_31;
    _zz_io_MatrixB_58_33 <= _zz_io_MatrixB_58_32;
    _zz_io_MatrixB_58_34 <= _zz_io_MatrixB_58_33;
    _zz_io_MatrixB_58_35 <= _zz_io_MatrixB_58_34;
    _zz_io_MatrixB_58_36 <= _zz_io_MatrixB_58_35;
    _zz_io_MatrixB_58_37 <= _zz_io_MatrixB_58_36;
    _zz_io_MatrixB_58_38 <= _zz_io_MatrixB_58_37;
    _zz_io_MatrixB_58_39 <= _zz_io_MatrixB_58_38;
    _zz_io_MatrixB_58_40 <= _zz_io_MatrixB_58_39;
    _zz_io_MatrixB_58_41 <= _zz_io_MatrixB_58_40;
    _zz_io_MatrixB_58_42 <= _zz_io_MatrixB_58_41;
    _zz_io_MatrixB_58_43 <= _zz_io_MatrixB_58_42;
    _zz_io_MatrixB_58_44 <= _zz_io_MatrixB_58_43;
    _zz_io_MatrixB_58_45 <= _zz_io_MatrixB_58_44;
    _zz_io_MatrixB_58_46 <= _zz_io_MatrixB_58_45;
    _zz_io_MatrixB_58_47 <= _zz_io_MatrixB_58_46;
    _zz_io_MatrixB_58_48 <= _zz_io_MatrixB_58_47;
    _zz_io_MatrixB_58_49 <= _zz_io_MatrixB_58_48;
    _zz_io_MatrixB_58_50 <= _zz_io_MatrixB_58_49;
    _zz_io_MatrixB_58_51 <= _zz_io_MatrixB_58_50;
    _zz_io_MatrixB_58_52 <= _zz_io_MatrixB_58_51;
    _zz_io_MatrixB_58_53 <= _zz_io_MatrixB_58_52;
    _zz_io_MatrixB_58_54 <= _zz_io_MatrixB_58_53;
    _zz_io_MatrixB_58_55 <= _zz_io_MatrixB_58_54;
    _zz_io_MatrixB_58_56 <= _zz_io_MatrixB_58_55;
    _zz_io_MatrixB_58_57 <= _zz_io_MatrixB_58_56;
    _zz_io_B_Valid_58 <= SubModule_WeightCache_MatrixCol_Switch[58];
    _zz_io_B_Valid_58_1 <= _zz_io_B_Valid_58;
    _zz_io_B_Valid_58_2 <= _zz_io_B_Valid_58_1;
    _zz_io_B_Valid_58_3 <= _zz_io_B_Valid_58_2;
    _zz_io_B_Valid_58_4 <= _zz_io_B_Valid_58_3;
    _zz_io_B_Valid_58_5 <= _zz_io_B_Valid_58_4;
    _zz_io_B_Valid_58_6 <= _zz_io_B_Valid_58_5;
    _zz_io_B_Valid_58_7 <= _zz_io_B_Valid_58_6;
    _zz_io_B_Valid_58_8 <= _zz_io_B_Valid_58_7;
    _zz_io_B_Valid_58_9 <= _zz_io_B_Valid_58_8;
    _zz_io_B_Valid_58_10 <= _zz_io_B_Valid_58_9;
    _zz_io_B_Valid_58_11 <= _zz_io_B_Valid_58_10;
    _zz_io_B_Valid_58_12 <= _zz_io_B_Valid_58_11;
    _zz_io_B_Valid_58_13 <= _zz_io_B_Valid_58_12;
    _zz_io_B_Valid_58_14 <= _zz_io_B_Valid_58_13;
    _zz_io_B_Valid_58_15 <= _zz_io_B_Valid_58_14;
    _zz_io_B_Valid_58_16 <= _zz_io_B_Valid_58_15;
    _zz_io_B_Valid_58_17 <= _zz_io_B_Valid_58_16;
    _zz_io_B_Valid_58_18 <= _zz_io_B_Valid_58_17;
    _zz_io_B_Valid_58_19 <= _zz_io_B_Valid_58_18;
    _zz_io_B_Valid_58_20 <= _zz_io_B_Valid_58_19;
    _zz_io_B_Valid_58_21 <= _zz_io_B_Valid_58_20;
    _zz_io_B_Valid_58_22 <= _zz_io_B_Valid_58_21;
    _zz_io_B_Valid_58_23 <= _zz_io_B_Valid_58_22;
    _zz_io_B_Valid_58_24 <= _zz_io_B_Valid_58_23;
    _zz_io_B_Valid_58_25 <= _zz_io_B_Valid_58_24;
    _zz_io_B_Valid_58_26 <= _zz_io_B_Valid_58_25;
    _zz_io_B_Valid_58_27 <= _zz_io_B_Valid_58_26;
    _zz_io_B_Valid_58_28 <= _zz_io_B_Valid_58_27;
    _zz_io_B_Valid_58_29 <= _zz_io_B_Valid_58_28;
    _zz_io_B_Valid_58_30 <= _zz_io_B_Valid_58_29;
    _zz_io_B_Valid_58_31 <= _zz_io_B_Valid_58_30;
    _zz_io_B_Valid_58_32 <= _zz_io_B_Valid_58_31;
    _zz_io_B_Valid_58_33 <= _zz_io_B_Valid_58_32;
    _zz_io_B_Valid_58_34 <= _zz_io_B_Valid_58_33;
    _zz_io_B_Valid_58_35 <= _zz_io_B_Valid_58_34;
    _zz_io_B_Valid_58_36 <= _zz_io_B_Valid_58_35;
    _zz_io_B_Valid_58_37 <= _zz_io_B_Valid_58_36;
    _zz_io_B_Valid_58_38 <= _zz_io_B_Valid_58_37;
    _zz_io_B_Valid_58_39 <= _zz_io_B_Valid_58_38;
    _zz_io_B_Valid_58_40 <= _zz_io_B_Valid_58_39;
    _zz_io_B_Valid_58_41 <= _zz_io_B_Valid_58_40;
    _zz_io_B_Valid_58_42 <= _zz_io_B_Valid_58_41;
    _zz_io_B_Valid_58_43 <= _zz_io_B_Valid_58_42;
    _zz_io_B_Valid_58_44 <= _zz_io_B_Valid_58_43;
    _zz_io_B_Valid_58_45 <= _zz_io_B_Valid_58_44;
    _zz_io_B_Valid_58_46 <= _zz_io_B_Valid_58_45;
    _zz_io_B_Valid_58_47 <= _zz_io_B_Valid_58_46;
    _zz_io_B_Valid_58_48 <= _zz_io_B_Valid_58_47;
    _zz_io_B_Valid_58_49 <= _zz_io_B_Valid_58_48;
    _zz_io_B_Valid_58_50 <= _zz_io_B_Valid_58_49;
    _zz_io_B_Valid_58_51 <= _zz_io_B_Valid_58_50;
    _zz_io_B_Valid_58_52 <= _zz_io_B_Valid_58_51;
    _zz_io_B_Valid_58_53 <= _zz_io_B_Valid_58_52;
    _zz_io_B_Valid_58_54 <= _zz_io_B_Valid_58_53;
    _zz_io_B_Valid_58_55 <= _zz_io_B_Valid_58_54;
    _zz_io_B_Valid_58_56 <= _zz_io_B_Valid_58_55;
    _zz_io_B_Valid_58_57 <= _zz_io_B_Valid_58_56;
    _zz_io_MatrixB_59 <= SubModule_WeightCache_mData_59;
    _zz_io_MatrixB_59_1 <= _zz_io_MatrixB_59;
    _zz_io_MatrixB_59_2 <= _zz_io_MatrixB_59_1;
    _zz_io_MatrixB_59_3 <= _zz_io_MatrixB_59_2;
    _zz_io_MatrixB_59_4 <= _zz_io_MatrixB_59_3;
    _zz_io_MatrixB_59_5 <= _zz_io_MatrixB_59_4;
    _zz_io_MatrixB_59_6 <= _zz_io_MatrixB_59_5;
    _zz_io_MatrixB_59_7 <= _zz_io_MatrixB_59_6;
    _zz_io_MatrixB_59_8 <= _zz_io_MatrixB_59_7;
    _zz_io_MatrixB_59_9 <= _zz_io_MatrixB_59_8;
    _zz_io_MatrixB_59_10 <= _zz_io_MatrixB_59_9;
    _zz_io_MatrixB_59_11 <= _zz_io_MatrixB_59_10;
    _zz_io_MatrixB_59_12 <= _zz_io_MatrixB_59_11;
    _zz_io_MatrixB_59_13 <= _zz_io_MatrixB_59_12;
    _zz_io_MatrixB_59_14 <= _zz_io_MatrixB_59_13;
    _zz_io_MatrixB_59_15 <= _zz_io_MatrixB_59_14;
    _zz_io_MatrixB_59_16 <= _zz_io_MatrixB_59_15;
    _zz_io_MatrixB_59_17 <= _zz_io_MatrixB_59_16;
    _zz_io_MatrixB_59_18 <= _zz_io_MatrixB_59_17;
    _zz_io_MatrixB_59_19 <= _zz_io_MatrixB_59_18;
    _zz_io_MatrixB_59_20 <= _zz_io_MatrixB_59_19;
    _zz_io_MatrixB_59_21 <= _zz_io_MatrixB_59_20;
    _zz_io_MatrixB_59_22 <= _zz_io_MatrixB_59_21;
    _zz_io_MatrixB_59_23 <= _zz_io_MatrixB_59_22;
    _zz_io_MatrixB_59_24 <= _zz_io_MatrixB_59_23;
    _zz_io_MatrixB_59_25 <= _zz_io_MatrixB_59_24;
    _zz_io_MatrixB_59_26 <= _zz_io_MatrixB_59_25;
    _zz_io_MatrixB_59_27 <= _zz_io_MatrixB_59_26;
    _zz_io_MatrixB_59_28 <= _zz_io_MatrixB_59_27;
    _zz_io_MatrixB_59_29 <= _zz_io_MatrixB_59_28;
    _zz_io_MatrixB_59_30 <= _zz_io_MatrixB_59_29;
    _zz_io_MatrixB_59_31 <= _zz_io_MatrixB_59_30;
    _zz_io_MatrixB_59_32 <= _zz_io_MatrixB_59_31;
    _zz_io_MatrixB_59_33 <= _zz_io_MatrixB_59_32;
    _zz_io_MatrixB_59_34 <= _zz_io_MatrixB_59_33;
    _zz_io_MatrixB_59_35 <= _zz_io_MatrixB_59_34;
    _zz_io_MatrixB_59_36 <= _zz_io_MatrixB_59_35;
    _zz_io_MatrixB_59_37 <= _zz_io_MatrixB_59_36;
    _zz_io_MatrixB_59_38 <= _zz_io_MatrixB_59_37;
    _zz_io_MatrixB_59_39 <= _zz_io_MatrixB_59_38;
    _zz_io_MatrixB_59_40 <= _zz_io_MatrixB_59_39;
    _zz_io_MatrixB_59_41 <= _zz_io_MatrixB_59_40;
    _zz_io_MatrixB_59_42 <= _zz_io_MatrixB_59_41;
    _zz_io_MatrixB_59_43 <= _zz_io_MatrixB_59_42;
    _zz_io_MatrixB_59_44 <= _zz_io_MatrixB_59_43;
    _zz_io_MatrixB_59_45 <= _zz_io_MatrixB_59_44;
    _zz_io_MatrixB_59_46 <= _zz_io_MatrixB_59_45;
    _zz_io_MatrixB_59_47 <= _zz_io_MatrixB_59_46;
    _zz_io_MatrixB_59_48 <= _zz_io_MatrixB_59_47;
    _zz_io_MatrixB_59_49 <= _zz_io_MatrixB_59_48;
    _zz_io_MatrixB_59_50 <= _zz_io_MatrixB_59_49;
    _zz_io_MatrixB_59_51 <= _zz_io_MatrixB_59_50;
    _zz_io_MatrixB_59_52 <= _zz_io_MatrixB_59_51;
    _zz_io_MatrixB_59_53 <= _zz_io_MatrixB_59_52;
    _zz_io_MatrixB_59_54 <= _zz_io_MatrixB_59_53;
    _zz_io_MatrixB_59_55 <= _zz_io_MatrixB_59_54;
    _zz_io_MatrixB_59_56 <= _zz_io_MatrixB_59_55;
    _zz_io_MatrixB_59_57 <= _zz_io_MatrixB_59_56;
    _zz_io_MatrixB_59_58 <= _zz_io_MatrixB_59_57;
    _zz_io_B_Valid_59 <= SubModule_WeightCache_MatrixCol_Switch[59];
    _zz_io_B_Valid_59_1 <= _zz_io_B_Valid_59;
    _zz_io_B_Valid_59_2 <= _zz_io_B_Valid_59_1;
    _zz_io_B_Valid_59_3 <= _zz_io_B_Valid_59_2;
    _zz_io_B_Valid_59_4 <= _zz_io_B_Valid_59_3;
    _zz_io_B_Valid_59_5 <= _zz_io_B_Valid_59_4;
    _zz_io_B_Valid_59_6 <= _zz_io_B_Valid_59_5;
    _zz_io_B_Valid_59_7 <= _zz_io_B_Valid_59_6;
    _zz_io_B_Valid_59_8 <= _zz_io_B_Valid_59_7;
    _zz_io_B_Valid_59_9 <= _zz_io_B_Valid_59_8;
    _zz_io_B_Valid_59_10 <= _zz_io_B_Valid_59_9;
    _zz_io_B_Valid_59_11 <= _zz_io_B_Valid_59_10;
    _zz_io_B_Valid_59_12 <= _zz_io_B_Valid_59_11;
    _zz_io_B_Valid_59_13 <= _zz_io_B_Valid_59_12;
    _zz_io_B_Valid_59_14 <= _zz_io_B_Valid_59_13;
    _zz_io_B_Valid_59_15 <= _zz_io_B_Valid_59_14;
    _zz_io_B_Valid_59_16 <= _zz_io_B_Valid_59_15;
    _zz_io_B_Valid_59_17 <= _zz_io_B_Valid_59_16;
    _zz_io_B_Valid_59_18 <= _zz_io_B_Valid_59_17;
    _zz_io_B_Valid_59_19 <= _zz_io_B_Valid_59_18;
    _zz_io_B_Valid_59_20 <= _zz_io_B_Valid_59_19;
    _zz_io_B_Valid_59_21 <= _zz_io_B_Valid_59_20;
    _zz_io_B_Valid_59_22 <= _zz_io_B_Valid_59_21;
    _zz_io_B_Valid_59_23 <= _zz_io_B_Valid_59_22;
    _zz_io_B_Valid_59_24 <= _zz_io_B_Valid_59_23;
    _zz_io_B_Valid_59_25 <= _zz_io_B_Valid_59_24;
    _zz_io_B_Valid_59_26 <= _zz_io_B_Valid_59_25;
    _zz_io_B_Valid_59_27 <= _zz_io_B_Valid_59_26;
    _zz_io_B_Valid_59_28 <= _zz_io_B_Valid_59_27;
    _zz_io_B_Valid_59_29 <= _zz_io_B_Valid_59_28;
    _zz_io_B_Valid_59_30 <= _zz_io_B_Valid_59_29;
    _zz_io_B_Valid_59_31 <= _zz_io_B_Valid_59_30;
    _zz_io_B_Valid_59_32 <= _zz_io_B_Valid_59_31;
    _zz_io_B_Valid_59_33 <= _zz_io_B_Valid_59_32;
    _zz_io_B_Valid_59_34 <= _zz_io_B_Valid_59_33;
    _zz_io_B_Valid_59_35 <= _zz_io_B_Valid_59_34;
    _zz_io_B_Valid_59_36 <= _zz_io_B_Valid_59_35;
    _zz_io_B_Valid_59_37 <= _zz_io_B_Valid_59_36;
    _zz_io_B_Valid_59_38 <= _zz_io_B_Valid_59_37;
    _zz_io_B_Valid_59_39 <= _zz_io_B_Valid_59_38;
    _zz_io_B_Valid_59_40 <= _zz_io_B_Valid_59_39;
    _zz_io_B_Valid_59_41 <= _zz_io_B_Valid_59_40;
    _zz_io_B_Valid_59_42 <= _zz_io_B_Valid_59_41;
    _zz_io_B_Valid_59_43 <= _zz_io_B_Valid_59_42;
    _zz_io_B_Valid_59_44 <= _zz_io_B_Valid_59_43;
    _zz_io_B_Valid_59_45 <= _zz_io_B_Valid_59_44;
    _zz_io_B_Valid_59_46 <= _zz_io_B_Valid_59_45;
    _zz_io_B_Valid_59_47 <= _zz_io_B_Valid_59_46;
    _zz_io_B_Valid_59_48 <= _zz_io_B_Valid_59_47;
    _zz_io_B_Valid_59_49 <= _zz_io_B_Valid_59_48;
    _zz_io_B_Valid_59_50 <= _zz_io_B_Valid_59_49;
    _zz_io_B_Valid_59_51 <= _zz_io_B_Valid_59_50;
    _zz_io_B_Valid_59_52 <= _zz_io_B_Valid_59_51;
    _zz_io_B_Valid_59_53 <= _zz_io_B_Valid_59_52;
    _zz_io_B_Valid_59_54 <= _zz_io_B_Valid_59_53;
    _zz_io_B_Valid_59_55 <= _zz_io_B_Valid_59_54;
    _zz_io_B_Valid_59_56 <= _zz_io_B_Valid_59_55;
    _zz_io_B_Valid_59_57 <= _zz_io_B_Valid_59_56;
    _zz_io_B_Valid_59_58 <= _zz_io_B_Valid_59_57;
    _zz_io_MatrixB_60 <= SubModule_WeightCache_mData_60;
    _zz_io_MatrixB_60_1 <= _zz_io_MatrixB_60;
    _zz_io_MatrixB_60_2 <= _zz_io_MatrixB_60_1;
    _zz_io_MatrixB_60_3 <= _zz_io_MatrixB_60_2;
    _zz_io_MatrixB_60_4 <= _zz_io_MatrixB_60_3;
    _zz_io_MatrixB_60_5 <= _zz_io_MatrixB_60_4;
    _zz_io_MatrixB_60_6 <= _zz_io_MatrixB_60_5;
    _zz_io_MatrixB_60_7 <= _zz_io_MatrixB_60_6;
    _zz_io_MatrixB_60_8 <= _zz_io_MatrixB_60_7;
    _zz_io_MatrixB_60_9 <= _zz_io_MatrixB_60_8;
    _zz_io_MatrixB_60_10 <= _zz_io_MatrixB_60_9;
    _zz_io_MatrixB_60_11 <= _zz_io_MatrixB_60_10;
    _zz_io_MatrixB_60_12 <= _zz_io_MatrixB_60_11;
    _zz_io_MatrixB_60_13 <= _zz_io_MatrixB_60_12;
    _zz_io_MatrixB_60_14 <= _zz_io_MatrixB_60_13;
    _zz_io_MatrixB_60_15 <= _zz_io_MatrixB_60_14;
    _zz_io_MatrixB_60_16 <= _zz_io_MatrixB_60_15;
    _zz_io_MatrixB_60_17 <= _zz_io_MatrixB_60_16;
    _zz_io_MatrixB_60_18 <= _zz_io_MatrixB_60_17;
    _zz_io_MatrixB_60_19 <= _zz_io_MatrixB_60_18;
    _zz_io_MatrixB_60_20 <= _zz_io_MatrixB_60_19;
    _zz_io_MatrixB_60_21 <= _zz_io_MatrixB_60_20;
    _zz_io_MatrixB_60_22 <= _zz_io_MatrixB_60_21;
    _zz_io_MatrixB_60_23 <= _zz_io_MatrixB_60_22;
    _zz_io_MatrixB_60_24 <= _zz_io_MatrixB_60_23;
    _zz_io_MatrixB_60_25 <= _zz_io_MatrixB_60_24;
    _zz_io_MatrixB_60_26 <= _zz_io_MatrixB_60_25;
    _zz_io_MatrixB_60_27 <= _zz_io_MatrixB_60_26;
    _zz_io_MatrixB_60_28 <= _zz_io_MatrixB_60_27;
    _zz_io_MatrixB_60_29 <= _zz_io_MatrixB_60_28;
    _zz_io_MatrixB_60_30 <= _zz_io_MatrixB_60_29;
    _zz_io_MatrixB_60_31 <= _zz_io_MatrixB_60_30;
    _zz_io_MatrixB_60_32 <= _zz_io_MatrixB_60_31;
    _zz_io_MatrixB_60_33 <= _zz_io_MatrixB_60_32;
    _zz_io_MatrixB_60_34 <= _zz_io_MatrixB_60_33;
    _zz_io_MatrixB_60_35 <= _zz_io_MatrixB_60_34;
    _zz_io_MatrixB_60_36 <= _zz_io_MatrixB_60_35;
    _zz_io_MatrixB_60_37 <= _zz_io_MatrixB_60_36;
    _zz_io_MatrixB_60_38 <= _zz_io_MatrixB_60_37;
    _zz_io_MatrixB_60_39 <= _zz_io_MatrixB_60_38;
    _zz_io_MatrixB_60_40 <= _zz_io_MatrixB_60_39;
    _zz_io_MatrixB_60_41 <= _zz_io_MatrixB_60_40;
    _zz_io_MatrixB_60_42 <= _zz_io_MatrixB_60_41;
    _zz_io_MatrixB_60_43 <= _zz_io_MatrixB_60_42;
    _zz_io_MatrixB_60_44 <= _zz_io_MatrixB_60_43;
    _zz_io_MatrixB_60_45 <= _zz_io_MatrixB_60_44;
    _zz_io_MatrixB_60_46 <= _zz_io_MatrixB_60_45;
    _zz_io_MatrixB_60_47 <= _zz_io_MatrixB_60_46;
    _zz_io_MatrixB_60_48 <= _zz_io_MatrixB_60_47;
    _zz_io_MatrixB_60_49 <= _zz_io_MatrixB_60_48;
    _zz_io_MatrixB_60_50 <= _zz_io_MatrixB_60_49;
    _zz_io_MatrixB_60_51 <= _zz_io_MatrixB_60_50;
    _zz_io_MatrixB_60_52 <= _zz_io_MatrixB_60_51;
    _zz_io_MatrixB_60_53 <= _zz_io_MatrixB_60_52;
    _zz_io_MatrixB_60_54 <= _zz_io_MatrixB_60_53;
    _zz_io_MatrixB_60_55 <= _zz_io_MatrixB_60_54;
    _zz_io_MatrixB_60_56 <= _zz_io_MatrixB_60_55;
    _zz_io_MatrixB_60_57 <= _zz_io_MatrixB_60_56;
    _zz_io_MatrixB_60_58 <= _zz_io_MatrixB_60_57;
    _zz_io_MatrixB_60_59 <= _zz_io_MatrixB_60_58;
    _zz_io_B_Valid_60 <= SubModule_WeightCache_MatrixCol_Switch[60];
    _zz_io_B_Valid_60_1 <= _zz_io_B_Valid_60;
    _zz_io_B_Valid_60_2 <= _zz_io_B_Valid_60_1;
    _zz_io_B_Valid_60_3 <= _zz_io_B_Valid_60_2;
    _zz_io_B_Valid_60_4 <= _zz_io_B_Valid_60_3;
    _zz_io_B_Valid_60_5 <= _zz_io_B_Valid_60_4;
    _zz_io_B_Valid_60_6 <= _zz_io_B_Valid_60_5;
    _zz_io_B_Valid_60_7 <= _zz_io_B_Valid_60_6;
    _zz_io_B_Valid_60_8 <= _zz_io_B_Valid_60_7;
    _zz_io_B_Valid_60_9 <= _zz_io_B_Valid_60_8;
    _zz_io_B_Valid_60_10 <= _zz_io_B_Valid_60_9;
    _zz_io_B_Valid_60_11 <= _zz_io_B_Valid_60_10;
    _zz_io_B_Valid_60_12 <= _zz_io_B_Valid_60_11;
    _zz_io_B_Valid_60_13 <= _zz_io_B_Valid_60_12;
    _zz_io_B_Valid_60_14 <= _zz_io_B_Valid_60_13;
    _zz_io_B_Valid_60_15 <= _zz_io_B_Valid_60_14;
    _zz_io_B_Valid_60_16 <= _zz_io_B_Valid_60_15;
    _zz_io_B_Valid_60_17 <= _zz_io_B_Valid_60_16;
    _zz_io_B_Valid_60_18 <= _zz_io_B_Valid_60_17;
    _zz_io_B_Valid_60_19 <= _zz_io_B_Valid_60_18;
    _zz_io_B_Valid_60_20 <= _zz_io_B_Valid_60_19;
    _zz_io_B_Valid_60_21 <= _zz_io_B_Valid_60_20;
    _zz_io_B_Valid_60_22 <= _zz_io_B_Valid_60_21;
    _zz_io_B_Valid_60_23 <= _zz_io_B_Valid_60_22;
    _zz_io_B_Valid_60_24 <= _zz_io_B_Valid_60_23;
    _zz_io_B_Valid_60_25 <= _zz_io_B_Valid_60_24;
    _zz_io_B_Valid_60_26 <= _zz_io_B_Valid_60_25;
    _zz_io_B_Valid_60_27 <= _zz_io_B_Valid_60_26;
    _zz_io_B_Valid_60_28 <= _zz_io_B_Valid_60_27;
    _zz_io_B_Valid_60_29 <= _zz_io_B_Valid_60_28;
    _zz_io_B_Valid_60_30 <= _zz_io_B_Valid_60_29;
    _zz_io_B_Valid_60_31 <= _zz_io_B_Valid_60_30;
    _zz_io_B_Valid_60_32 <= _zz_io_B_Valid_60_31;
    _zz_io_B_Valid_60_33 <= _zz_io_B_Valid_60_32;
    _zz_io_B_Valid_60_34 <= _zz_io_B_Valid_60_33;
    _zz_io_B_Valid_60_35 <= _zz_io_B_Valid_60_34;
    _zz_io_B_Valid_60_36 <= _zz_io_B_Valid_60_35;
    _zz_io_B_Valid_60_37 <= _zz_io_B_Valid_60_36;
    _zz_io_B_Valid_60_38 <= _zz_io_B_Valid_60_37;
    _zz_io_B_Valid_60_39 <= _zz_io_B_Valid_60_38;
    _zz_io_B_Valid_60_40 <= _zz_io_B_Valid_60_39;
    _zz_io_B_Valid_60_41 <= _zz_io_B_Valid_60_40;
    _zz_io_B_Valid_60_42 <= _zz_io_B_Valid_60_41;
    _zz_io_B_Valid_60_43 <= _zz_io_B_Valid_60_42;
    _zz_io_B_Valid_60_44 <= _zz_io_B_Valid_60_43;
    _zz_io_B_Valid_60_45 <= _zz_io_B_Valid_60_44;
    _zz_io_B_Valid_60_46 <= _zz_io_B_Valid_60_45;
    _zz_io_B_Valid_60_47 <= _zz_io_B_Valid_60_46;
    _zz_io_B_Valid_60_48 <= _zz_io_B_Valid_60_47;
    _zz_io_B_Valid_60_49 <= _zz_io_B_Valid_60_48;
    _zz_io_B_Valid_60_50 <= _zz_io_B_Valid_60_49;
    _zz_io_B_Valid_60_51 <= _zz_io_B_Valid_60_50;
    _zz_io_B_Valid_60_52 <= _zz_io_B_Valid_60_51;
    _zz_io_B_Valid_60_53 <= _zz_io_B_Valid_60_52;
    _zz_io_B_Valid_60_54 <= _zz_io_B_Valid_60_53;
    _zz_io_B_Valid_60_55 <= _zz_io_B_Valid_60_54;
    _zz_io_B_Valid_60_56 <= _zz_io_B_Valid_60_55;
    _zz_io_B_Valid_60_57 <= _zz_io_B_Valid_60_56;
    _zz_io_B_Valid_60_58 <= _zz_io_B_Valid_60_57;
    _zz_io_B_Valid_60_59 <= _zz_io_B_Valid_60_58;
    _zz_io_MatrixB_61 <= SubModule_WeightCache_mData_61;
    _zz_io_MatrixB_61_1 <= _zz_io_MatrixB_61;
    _zz_io_MatrixB_61_2 <= _zz_io_MatrixB_61_1;
    _zz_io_MatrixB_61_3 <= _zz_io_MatrixB_61_2;
    _zz_io_MatrixB_61_4 <= _zz_io_MatrixB_61_3;
    _zz_io_MatrixB_61_5 <= _zz_io_MatrixB_61_4;
    _zz_io_MatrixB_61_6 <= _zz_io_MatrixB_61_5;
    _zz_io_MatrixB_61_7 <= _zz_io_MatrixB_61_6;
    _zz_io_MatrixB_61_8 <= _zz_io_MatrixB_61_7;
    _zz_io_MatrixB_61_9 <= _zz_io_MatrixB_61_8;
    _zz_io_MatrixB_61_10 <= _zz_io_MatrixB_61_9;
    _zz_io_MatrixB_61_11 <= _zz_io_MatrixB_61_10;
    _zz_io_MatrixB_61_12 <= _zz_io_MatrixB_61_11;
    _zz_io_MatrixB_61_13 <= _zz_io_MatrixB_61_12;
    _zz_io_MatrixB_61_14 <= _zz_io_MatrixB_61_13;
    _zz_io_MatrixB_61_15 <= _zz_io_MatrixB_61_14;
    _zz_io_MatrixB_61_16 <= _zz_io_MatrixB_61_15;
    _zz_io_MatrixB_61_17 <= _zz_io_MatrixB_61_16;
    _zz_io_MatrixB_61_18 <= _zz_io_MatrixB_61_17;
    _zz_io_MatrixB_61_19 <= _zz_io_MatrixB_61_18;
    _zz_io_MatrixB_61_20 <= _zz_io_MatrixB_61_19;
    _zz_io_MatrixB_61_21 <= _zz_io_MatrixB_61_20;
    _zz_io_MatrixB_61_22 <= _zz_io_MatrixB_61_21;
    _zz_io_MatrixB_61_23 <= _zz_io_MatrixB_61_22;
    _zz_io_MatrixB_61_24 <= _zz_io_MatrixB_61_23;
    _zz_io_MatrixB_61_25 <= _zz_io_MatrixB_61_24;
    _zz_io_MatrixB_61_26 <= _zz_io_MatrixB_61_25;
    _zz_io_MatrixB_61_27 <= _zz_io_MatrixB_61_26;
    _zz_io_MatrixB_61_28 <= _zz_io_MatrixB_61_27;
    _zz_io_MatrixB_61_29 <= _zz_io_MatrixB_61_28;
    _zz_io_MatrixB_61_30 <= _zz_io_MatrixB_61_29;
    _zz_io_MatrixB_61_31 <= _zz_io_MatrixB_61_30;
    _zz_io_MatrixB_61_32 <= _zz_io_MatrixB_61_31;
    _zz_io_MatrixB_61_33 <= _zz_io_MatrixB_61_32;
    _zz_io_MatrixB_61_34 <= _zz_io_MatrixB_61_33;
    _zz_io_MatrixB_61_35 <= _zz_io_MatrixB_61_34;
    _zz_io_MatrixB_61_36 <= _zz_io_MatrixB_61_35;
    _zz_io_MatrixB_61_37 <= _zz_io_MatrixB_61_36;
    _zz_io_MatrixB_61_38 <= _zz_io_MatrixB_61_37;
    _zz_io_MatrixB_61_39 <= _zz_io_MatrixB_61_38;
    _zz_io_MatrixB_61_40 <= _zz_io_MatrixB_61_39;
    _zz_io_MatrixB_61_41 <= _zz_io_MatrixB_61_40;
    _zz_io_MatrixB_61_42 <= _zz_io_MatrixB_61_41;
    _zz_io_MatrixB_61_43 <= _zz_io_MatrixB_61_42;
    _zz_io_MatrixB_61_44 <= _zz_io_MatrixB_61_43;
    _zz_io_MatrixB_61_45 <= _zz_io_MatrixB_61_44;
    _zz_io_MatrixB_61_46 <= _zz_io_MatrixB_61_45;
    _zz_io_MatrixB_61_47 <= _zz_io_MatrixB_61_46;
    _zz_io_MatrixB_61_48 <= _zz_io_MatrixB_61_47;
    _zz_io_MatrixB_61_49 <= _zz_io_MatrixB_61_48;
    _zz_io_MatrixB_61_50 <= _zz_io_MatrixB_61_49;
    _zz_io_MatrixB_61_51 <= _zz_io_MatrixB_61_50;
    _zz_io_MatrixB_61_52 <= _zz_io_MatrixB_61_51;
    _zz_io_MatrixB_61_53 <= _zz_io_MatrixB_61_52;
    _zz_io_MatrixB_61_54 <= _zz_io_MatrixB_61_53;
    _zz_io_MatrixB_61_55 <= _zz_io_MatrixB_61_54;
    _zz_io_MatrixB_61_56 <= _zz_io_MatrixB_61_55;
    _zz_io_MatrixB_61_57 <= _zz_io_MatrixB_61_56;
    _zz_io_MatrixB_61_58 <= _zz_io_MatrixB_61_57;
    _zz_io_MatrixB_61_59 <= _zz_io_MatrixB_61_58;
    _zz_io_MatrixB_61_60 <= _zz_io_MatrixB_61_59;
    _zz_io_B_Valid_61 <= SubModule_WeightCache_MatrixCol_Switch[61];
    _zz_io_B_Valid_61_1 <= _zz_io_B_Valid_61;
    _zz_io_B_Valid_61_2 <= _zz_io_B_Valid_61_1;
    _zz_io_B_Valid_61_3 <= _zz_io_B_Valid_61_2;
    _zz_io_B_Valid_61_4 <= _zz_io_B_Valid_61_3;
    _zz_io_B_Valid_61_5 <= _zz_io_B_Valid_61_4;
    _zz_io_B_Valid_61_6 <= _zz_io_B_Valid_61_5;
    _zz_io_B_Valid_61_7 <= _zz_io_B_Valid_61_6;
    _zz_io_B_Valid_61_8 <= _zz_io_B_Valid_61_7;
    _zz_io_B_Valid_61_9 <= _zz_io_B_Valid_61_8;
    _zz_io_B_Valid_61_10 <= _zz_io_B_Valid_61_9;
    _zz_io_B_Valid_61_11 <= _zz_io_B_Valid_61_10;
    _zz_io_B_Valid_61_12 <= _zz_io_B_Valid_61_11;
    _zz_io_B_Valid_61_13 <= _zz_io_B_Valid_61_12;
    _zz_io_B_Valid_61_14 <= _zz_io_B_Valid_61_13;
    _zz_io_B_Valid_61_15 <= _zz_io_B_Valid_61_14;
    _zz_io_B_Valid_61_16 <= _zz_io_B_Valid_61_15;
    _zz_io_B_Valid_61_17 <= _zz_io_B_Valid_61_16;
    _zz_io_B_Valid_61_18 <= _zz_io_B_Valid_61_17;
    _zz_io_B_Valid_61_19 <= _zz_io_B_Valid_61_18;
    _zz_io_B_Valid_61_20 <= _zz_io_B_Valid_61_19;
    _zz_io_B_Valid_61_21 <= _zz_io_B_Valid_61_20;
    _zz_io_B_Valid_61_22 <= _zz_io_B_Valid_61_21;
    _zz_io_B_Valid_61_23 <= _zz_io_B_Valid_61_22;
    _zz_io_B_Valid_61_24 <= _zz_io_B_Valid_61_23;
    _zz_io_B_Valid_61_25 <= _zz_io_B_Valid_61_24;
    _zz_io_B_Valid_61_26 <= _zz_io_B_Valid_61_25;
    _zz_io_B_Valid_61_27 <= _zz_io_B_Valid_61_26;
    _zz_io_B_Valid_61_28 <= _zz_io_B_Valid_61_27;
    _zz_io_B_Valid_61_29 <= _zz_io_B_Valid_61_28;
    _zz_io_B_Valid_61_30 <= _zz_io_B_Valid_61_29;
    _zz_io_B_Valid_61_31 <= _zz_io_B_Valid_61_30;
    _zz_io_B_Valid_61_32 <= _zz_io_B_Valid_61_31;
    _zz_io_B_Valid_61_33 <= _zz_io_B_Valid_61_32;
    _zz_io_B_Valid_61_34 <= _zz_io_B_Valid_61_33;
    _zz_io_B_Valid_61_35 <= _zz_io_B_Valid_61_34;
    _zz_io_B_Valid_61_36 <= _zz_io_B_Valid_61_35;
    _zz_io_B_Valid_61_37 <= _zz_io_B_Valid_61_36;
    _zz_io_B_Valid_61_38 <= _zz_io_B_Valid_61_37;
    _zz_io_B_Valid_61_39 <= _zz_io_B_Valid_61_38;
    _zz_io_B_Valid_61_40 <= _zz_io_B_Valid_61_39;
    _zz_io_B_Valid_61_41 <= _zz_io_B_Valid_61_40;
    _zz_io_B_Valid_61_42 <= _zz_io_B_Valid_61_41;
    _zz_io_B_Valid_61_43 <= _zz_io_B_Valid_61_42;
    _zz_io_B_Valid_61_44 <= _zz_io_B_Valid_61_43;
    _zz_io_B_Valid_61_45 <= _zz_io_B_Valid_61_44;
    _zz_io_B_Valid_61_46 <= _zz_io_B_Valid_61_45;
    _zz_io_B_Valid_61_47 <= _zz_io_B_Valid_61_46;
    _zz_io_B_Valid_61_48 <= _zz_io_B_Valid_61_47;
    _zz_io_B_Valid_61_49 <= _zz_io_B_Valid_61_48;
    _zz_io_B_Valid_61_50 <= _zz_io_B_Valid_61_49;
    _zz_io_B_Valid_61_51 <= _zz_io_B_Valid_61_50;
    _zz_io_B_Valid_61_52 <= _zz_io_B_Valid_61_51;
    _zz_io_B_Valid_61_53 <= _zz_io_B_Valid_61_52;
    _zz_io_B_Valid_61_54 <= _zz_io_B_Valid_61_53;
    _zz_io_B_Valid_61_55 <= _zz_io_B_Valid_61_54;
    _zz_io_B_Valid_61_56 <= _zz_io_B_Valid_61_55;
    _zz_io_B_Valid_61_57 <= _zz_io_B_Valid_61_56;
    _zz_io_B_Valid_61_58 <= _zz_io_B_Valid_61_57;
    _zz_io_B_Valid_61_59 <= _zz_io_B_Valid_61_58;
    _zz_io_B_Valid_61_60 <= _zz_io_B_Valid_61_59;
    _zz_io_MatrixB_62 <= SubModule_WeightCache_mData_62;
    _zz_io_MatrixB_62_1 <= _zz_io_MatrixB_62;
    _zz_io_MatrixB_62_2 <= _zz_io_MatrixB_62_1;
    _zz_io_MatrixB_62_3 <= _zz_io_MatrixB_62_2;
    _zz_io_MatrixB_62_4 <= _zz_io_MatrixB_62_3;
    _zz_io_MatrixB_62_5 <= _zz_io_MatrixB_62_4;
    _zz_io_MatrixB_62_6 <= _zz_io_MatrixB_62_5;
    _zz_io_MatrixB_62_7 <= _zz_io_MatrixB_62_6;
    _zz_io_MatrixB_62_8 <= _zz_io_MatrixB_62_7;
    _zz_io_MatrixB_62_9 <= _zz_io_MatrixB_62_8;
    _zz_io_MatrixB_62_10 <= _zz_io_MatrixB_62_9;
    _zz_io_MatrixB_62_11 <= _zz_io_MatrixB_62_10;
    _zz_io_MatrixB_62_12 <= _zz_io_MatrixB_62_11;
    _zz_io_MatrixB_62_13 <= _zz_io_MatrixB_62_12;
    _zz_io_MatrixB_62_14 <= _zz_io_MatrixB_62_13;
    _zz_io_MatrixB_62_15 <= _zz_io_MatrixB_62_14;
    _zz_io_MatrixB_62_16 <= _zz_io_MatrixB_62_15;
    _zz_io_MatrixB_62_17 <= _zz_io_MatrixB_62_16;
    _zz_io_MatrixB_62_18 <= _zz_io_MatrixB_62_17;
    _zz_io_MatrixB_62_19 <= _zz_io_MatrixB_62_18;
    _zz_io_MatrixB_62_20 <= _zz_io_MatrixB_62_19;
    _zz_io_MatrixB_62_21 <= _zz_io_MatrixB_62_20;
    _zz_io_MatrixB_62_22 <= _zz_io_MatrixB_62_21;
    _zz_io_MatrixB_62_23 <= _zz_io_MatrixB_62_22;
    _zz_io_MatrixB_62_24 <= _zz_io_MatrixB_62_23;
    _zz_io_MatrixB_62_25 <= _zz_io_MatrixB_62_24;
    _zz_io_MatrixB_62_26 <= _zz_io_MatrixB_62_25;
    _zz_io_MatrixB_62_27 <= _zz_io_MatrixB_62_26;
    _zz_io_MatrixB_62_28 <= _zz_io_MatrixB_62_27;
    _zz_io_MatrixB_62_29 <= _zz_io_MatrixB_62_28;
    _zz_io_MatrixB_62_30 <= _zz_io_MatrixB_62_29;
    _zz_io_MatrixB_62_31 <= _zz_io_MatrixB_62_30;
    _zz_io_MatrixB_62_32 <= _zz_io_MatrixB_62_31;
    _zz_io_MatrixB_62_33 <= _zz_io_MatrixB_62_32;
    _zz_io_MatrixB_62_34 <= _zz_io_MatrixB_62_33;
    _zz_io_MatrixB_62_35 <= _zz_io_MatrixB_62_34;
    _zz_io_MatrixB_62_36 <= _zz_io_MatrixB_62_35;
    _zz_io_MatrixB_62_37 <= _zz_io_MatrixB_62_36;
    _zz_io_MatrixB_62_38 <= _zz_io_MatrixB_62_37;
    _zz_io_MatrixB_62_39 <= _zz_io_MatrixB_62_38;
    _zz_io_MatrixB_62_40 <= _zz_io_MatrixB_62_39;
    _zz_io_MatrixB_62_41 <= _zz_io_MatrixB_62_40;
    _zz_io_MatrixB_62_42 <= _zz_io_MatrixB_62_41;
    _zz_io_MatrixB_62_43 <= _zz_io_MatrixB_62_42;
    _zz_io_MatrixB_62_44 <= _zz_io_MatrixB_62_43;
    _zz_io_MatrixB_62_45 <= _zz_io_MatrixB_62_44;
    _zz_io_MatrixB_62_46 <= _zz_io_MatrixB_62_45;
    _zz_io_MatrixB_62_47 <= _zz_io_MatrixB_62_46;
    _zz_io_MatrixB_62_48 <= _zz_io_MatrixB_62_47;
    _zz_io_MatrixB_62_49 <= _zz_io_MatrixB_62_48;
    _zz_io_MatrixB_62_50 <= _zz_io_MatrixB_62_49;
    _zz_io_MatrixB_62_51 <= _zz_io_MatrixB_62_50;
    _zz_io_MatrixB_62_52 <= _zz_io_MatrixB_62_51;
    _zz_io_MatrixB_62_53 <= _zz_io_MatrixB_62_52;
    _zz_io_MatrixB_62_54 <= _zz_io_MatrixB_62_53;
    _zz_io_MatrixB_62_55 <= _zz_io_MatrixB_62_54;
    _zz_io_MatrixB_62_56 <= _zz_io_MatrixB_62_55;
    _zz_io_MatrixB_62_57 <= _zz_io_MatrixB_62_56;
    _zz_io_MatrixB_62_58 <= _zz_io_MatrixB_62_57;
    _zz_io_MatrixB_62_59 <= _zz_io_MatrixB_62_58;
    _zz_io_MatrixB_62_60 <= _zz_io_MatrixB_62_59;
    _zz_io_MatrixB_62_61 <= _zz_io_MatrixB_62_60;
    _zz_io_B_Valid_62 <= SubModule_WeightCache_MatrixCol_Switch[62];
    _zz_io_B_Valid_62_1 <= _zz_io_B_Valid_62;
    _zz_io_B_Valid_62_2 <= _zz_io_B_Valid_62_1;
    _zz_io_B_Valid_62_3 <= _zz_io_B_Valid_62_2;
    _zz_io_B_Valid_62_4 <= _zz_io_B_Valid_62_3;
    _zz_io_B_Valid_62_5 <= _zz_io_B_Valid_62_4;
    _zz_io_B_Valid_62_6 <= _zz_io_B_Valid_62_5;
    _zz_io_B_Valid_62_7 <= _zz_io_B_Valid_62_6;
    _zz_io_B_Valid_62_8 <= _zz_io_B_Valid_62_7;
    _zz_io_B_Valid_62_9 <= _zz_io_B_Valid_62_8;
    _zz_io_B_Valid_62_10 <= _zz_io_B_Valid_62_9;
    _zz_io_B_Valid_62_11 <= _zz_io_B_Valid_62_10;
    _zz_io_B_Valid_62_12 <= _zz_io_B_Valid_62_11;
    _zz_io_B_Valid_62_13 <= _zz_io_B_Valid_62_12;
    _zz_io_B_Valid_62_14 <= _zz_io_B_Valid_62_13;
    _zz_io_B_Valid_62_15 <= _zz_io_B_Valid_62_14;
    _zz_io_B_Valid_62_16 <= _zz_io_B_Valid_62_15;
    _zz_io_B_Valid_62_17 <= _zz_io_B_Valid_62_16;
    _zz_io_B_Valid_62_18 <= _zz_io_B_Valid_62_17;
    _zz_io_B_Valid_62_19 <= _zz_io_B_Valid_62_18;
    _zz_io_B_Valid_62_20 <= _zz_io_B_Valid_62_19;
    _zz_io_B_Valid_62_21 <= _zz_io_B_Valid_62_20;
    _zz_io_B_Valid_62_22 <= _zz_io_B_Valid_62_21;
    _zz_io_B_Valid_62_23 <= _zz_io_B_Valid_62_22;
    _zz_io_B_Valid_62_24 <= _zz_io_B_Valid_62_23;
    _zz_io_B_Valid_62_25 <= _zz_io_B_Valid_62_24;
    _zz_io_B_Valid_62_26 <= _zz_io_B_Valid_62_25;
    _zz_io_B_Valid_62_27 <= _zz_io_B_Valid_62_26;
    _zz_io_B_Valid_62_28 <= _zz_io_B_Valid_62_27;
    _zz_io_B_Valid_62_29 <= _zz_io_B_Valid_62_28;
    _zz_io_B_Valid_62_30 <= _zz_io_B_Valid_62_29;
    _zz_io_B_Valid_62_31 <= _zz_io_B_Valid_62_30;
    _zz_io_B_Valid_62_32 <= _zz_io_B_Valid_62_31;
    _zz_io_B_Valid_62_33 <= _zz_io_B_Valid_62_32;
    _zz_io_B_Valid_62_34 <= _zz_io_B_Valid_62_33;
    _zz_io_B_Valid_62_35 <= _zz_io_B_Valid_62_34;
    _zz_io_B_Valid_62_36 <= _zz_io_B_Valid_62_35;
    _zz_io_B_Valid_62_37 <= _zz_io_B_Valid_62_36;
    _zz_io_B_Valid_62_38 <= _zz_io_B_Valid_62_37;
    _zz_io_B_Valid_62_39 <= _zz_io_B_Valid_62_38;
    _zz_io_B_Valid_62_40 <= _zz_io_B_Valid_62_39;
    _zz_io_B_Valid_62_41 <= _zz_io_B_Valid_62_40;
    _zz_io_B_Valid_62_42 <= _zz_io_B_Valid_62_41;
    _zz_io_B_Valid_62_43 <= _zz_io_B_Valid_62_42;
    _zz_io_B_Valid_62_44 <= _zz_io_B_Valid_62_43;
    _zz_io_B_Valid_62_45 <= _zz_io_B_Valid_62_44;
    _zz_io_B_Valid_62_46 <= _zz_io_B_Valid_62_45;
    _zz_io_B_Valid_62_47 <= _zz_io_B_Valid_62_46;
    _zz_io_B_Valid_62_48 <= _zz_io_B_Valid_62_47;
    _zz_io_B_Valid_62_49 <= _zz_io_B_Valid_62_48;
    _zz_io_B_Valid_62_50 <= _zz_io_B_Valid_62_49;
    _zz_io_B_Valid_62_51 <= _zz_io_B_Valid_62_50;
    _zz_io_B_Valid_62_52 <= _zz_io_B_Valid_62_51;
    _zz_io_B_Valid_62_53 <= _zz_io_B_Valid_62_52;
    _zz_io_B_Valid_62_54 <= _zz_io_B_Valid_62_53;
    _zz_io_B_Valid_62_55 <= _zz_io_B_Valid_62_54;
    _zz_io_B_Valid_62_56 <= _zz_io_B_Valid_62_55;
    _zz_io_B_Valid_62_57 <= _zz_io_B_Valid_62_56;
    _zz_io_B_Valid_62_58 <= _zz_io_B_Valid_62_57;
    _zz_io_B_Valid_62_59 <= _zz_io_B_Valid_62_58;
    _zz_io_B_Valid_62_60 <= _zz_io_B_Valid_62_59;
    _zz_io_B_Valid_62_61 <= _zz_io_B_Valid_62_60;
    _zz_io_MatrixB_63 <= SubModule_WeightCache_mData_63;
    _zz_io_MatrixB_63_1 <= _zz_io_MatrixB_63;
    _zz_io_MatrixB_63_2 <= _zz_io_MatrixB_63_1;
    _zz_io_MatrixB_63_3 <= _zz_io_MatrixB_63_2;
    _zz_io_MatrixB_63_4 <= _zz_io_MatrixB_63_3;
    _zz_io_MatrixB_63_5 <= _zz_io_MatrixB_63_4;
    _zz_io_MatrixB_63_6 <= _zz_io_MatrixB_63_5;
    _zz_io_MatrixB_63_7 <= _zz_io_MatrixB_63_6;
    _zz_io_MatrixB_63_8 <= _zz_io_MatrixB_63_7;
    _zz_io_MatrixB_63_9 <= _zz_io_MatrixB_63_8;
    _zz_io_MatrixB_63_10 <= _zz_io_MatrixB_63_9;
    _zz_io_MatrixB_63_11 <= _zz_io_MatrixB_63_10;
    _zz_io_MatrixB_63_12 <= _zz_io_MatrixB_63_11;
    _zz_io_MatrixB_63_13 <= _zz_io_MatrixB_63_12;
    _zz_io_MatrixB_63_14 <= _zz_io_MatrixB_63_13;
    _zz_io_MatrixB_63_15 <= _zz_io_MatrixB_63_14;
    _zz_io_MatrixB_63_16 <= _zz_io_MatrixB_63_15;
    _zz_io_MatrixB_63_17 <= _zz_io_MatrixB_63_16;
    _zz_io_MatrixB_63_18 <= _zz_io_MatrixB_63_17;
    _zz_io_MatrixB_63_19 <= _zz_io_MatrixB_63_18;
    _zz_io_MatrixB_63_20 <= _zz_io_MatrixB_63_19;
    _zz_io_MatrixB_63_21 <= _zz_io_MatrixB_63_20;
    _zz_io_MatrixB_63_22 <= _zz_io_MatrixB_63_21;
    _zz_io_MatrixB_63_23 <= _zz_io_MatrixB_63_22;
    _zz_io_MatrixB_63_24 <= _zz_io_MatrixB_63_23;
    _zz_io_MatrixB_63_25 <= _zz_io_MatrixB_63_24;
    _zz_io_MatrixB_63_26 <= _zz_io_MatrixB_63_25;
    _zz_io_MatrixB_63_27 <= _zz_io_MatrixB_63_26;
    _zz_io_MatrixB_63_28 <= _zz_io_MatrixB_63_27;
    _zz_io_MatrixB_63_29 <= _zz_io_MatrixB_63_28;
    _zz_io_MatrixB_63_30 <= _zz_io_MatrixB_63_29;
    _zz_io_MatrixB_63_31 <= _zz_io_MatrixB_63_30;
    _zz_io_MatrixB_63_32 <= _zz_io_MatrixB_63_31;
    _zz_io_MatrixB_63_33 <= _zz_io_MatrixB_63_32;
    _zz_io_MatrixB_63_34 <= _zz_io_MatrixB_63_33;
    _zz_io_MatrixB_63_35 <= _zz_io_MatrixB_63_34;
    _zz_io_MatrixB_63_36 <= _zz_io_MatrixB_63_35;
    _zz_io_MatrixB_63_37 <= _zz_io_MatrixB_63_36;
    _zz_io_MatrixB_63_38 <= _zz_io_MatrixB_63_37;
    _zz_io_MatrixB_63_39 <= _zz_io_MatrixB_63_38;
    _zz_io_MatrixB_63_40 <= _zz_io_MatrixB_63_39;
    _zz_io_MatrixB_63_41 <= _zz_io_MatrixB_63_40;
    _zz_io_MatrixB_63_42 <= _zz_io_MatrixB_63_41;
    _zz_io_MatrixB_63_43 <= _zz_io_MatrixB_63_42;
    _zz_io_MatrixB_63_44 <= _zz_io_MatrixB_63_43;
    _zz_io_MatrixB_63_45 <= _zz_io_MatrixB_63_44;
    _zz_io_MatrixB_63_46 <= _zz_io_MatrixB_63_45;
    _zz_io_MatrixB_63_47 <= _zz_io_MatrixB_63_46;
    _zz_io_MatrixB_63_48 <= _zz_io_MatrixB_63_47;
    _zz_io_MatrixB_63_49 <= _zz_io_MatrixB_63_48;
    _zz_io_MatrixB_63_50 <= _zz_io_MatrixB_63_49;
    _zz_io_MatrixB_63_51 <= _zz_io_MatrixB_63_50;
    _zz_io_MatrixB_63_52 <= _zz_io_MatrixB_63_51;
    _zz_io_MatrixB_63_53 <= _zz_io_MatrixB_63_52;
    _zz_io_MatrixB_63_54 <= _zz_io_MatrixB_63_53;
    _zz_io_MatrixB_63_55 <= _zz_io_MatrixB_63_54;
    _zz_io_MatrixB_63_56 <= _zz_io_MatrixB_63_55;
    _zz_io_MatrixB_63_57 <= _zz_io_MatrixB_63_56;
    _zz_io_MatrixB_63_58 <= _zz_io_MatrixB_63_57;
    _zz_io_MatrixB_63_59 <= _zz_io_MatrixB_63_58;
    _zz_io_MatrixB_63_60 <= _zz_io_MatrixB_63_59;
    _zz_io_MatrixB_63_61 <= _zz_io_MatrixB_63_60;
    _zz_io_MatrixB_63_62 <= _zz_io_MatrixB_63_61;
    _zz_io_B_Valid_63 <= SubModule_WeightCache_MatrixCol_Switch[63];
    _zz_io_B_Valid_63_1 <= _zz_io_B_Valid_63;
    _zz_io_B_Valid_63_2 <= _zz_io_B_Valid_63_1;
    _zz_io_B_Valid_63_3 <= _zz_io_B_Valid_63_2;
    _zz_io_B_Valid_63_4 <= _zz_io_B_Valid_63_3;
    _zz_io_B_Valid_63_5 <= _zz_io_B_Valid_63_4;
    _zz_io_B_Valid_63_6 <= _zz_io_B_Valid_63_5;
    _zz_io_B_Valid_63_7 <= _zz_io_B_Valid_63_6;
    _zz_io_B_Valid_63_8 <= _zz_io_B_Valid_63_7;
    _zz_io_B_Valid_63_9 <= _zz_io_B_Valid_63_8;
    _zz_io_B_Valid_63_10 <= _zz_io_B_Valid_63_9;
    _zz_io_B_Valid_63_11 <= _zz_io_B_Valid_63_10;
    _zz_io_B_Valid_63_12 <= _zz_io_B_Valid_63_11;
    _zz_io_B_Valid_63_13 <= _zz_io_B_Valid_63_12;
    _zz_io_B_Valid_63_14 <= _zz_io_B_Valid_63_13;
    _zz_io_B_Valid_63_15 <= _zz_io_B_Valid_63_14;
    _zz_io_B_Valid_63_16 <= _zz_io_B_Valid_63_15;
    _zz_io_B_Valid_63_17 <= _zz_io_B_Valid_63_16;
    _zz_io_B_Valid_63_18 <= _zz_io_B_Valid_63_17;
    _zz_io_B_Valid_63_19 <= _zz_io_B_Valid_63_18;
    _zz_io_B_Valid_63_20 <= _zz_io_B_Valid_63_19;
    _zz_io_B_Valid_63_21 <= _zz_io_B_Valid_63_20;
    _zz_io_B_Valid_63_22 <= _zz_io_B_Valid_63_21;
    _zz_io_B_Valid_63_23 <= _zz_io_B_Valid_63_22;
    _zz_io_B_Valid_63_24 <= _zz_io_B_Valid_63_23;
    _zz_io_B_Valid_63_25 <= _zz_io_B_Valid_63_24;
    _zz_io_B_Valid_63_26 <= _zz_io_B_Valid_63_25;
    _zz_io_B_Valid_63_27 <= _zz_io_B_Valid_63_26;
    _zz_io_B_Valid_63_28 <= _zz_io_B_Valid_63_27;
    _zz_io_B_Valid_63_29 <= _zz_io_B_Valid_63_28;
    _zz_io_B_Valid_63_30 <= _zz_io_B_Valid_63_29;
    _zz_io_B_Valid_63_31 <= _zz_io_B_Valid_63_30;
    _zz_io_B_Valid_63_32 <= _zz_io_B_Valid_63_31;
    _zz_io_B_Valid_63_33 <= _zz_io_B_Valid_63_32;
    _zz_io_B_Valid_63_34 <= _zz_io_B_Valid_63_33;
    _zz_io_B_Valid_63_35 <= _zz_io_B_Valid_63_34;
    _zz_io_B_Valid_63_36 <= _zz_io_B_Valid_63_35;
    _zz_io_B_Valid_63_37 <= _zz_io_B_Valid_63_36;
    _zz_io_B_Valid_63_38 <= _zz_io_B_Valid_63_37;
    _zz_io_B_Valid_63_39 <= _zz_io_B_Valid_63_38;
    _zz_io_B_Valid_63_40 <= _zz_io_B_Valid_63_39;
    _zz_io_B_Valid_63_41 <= _zz_io_B_Valid_63_40;
    _zz_io_B_Valid_63_42 <= _zz_io_B_Valid_63_41;
    _zz_io_B_Valid_63_43 <= _zz_io_B_Valid_63_42;
    _zz_io_B_Valid_63_44 <= _zz_io_B_Valid_63_43;
    _zz_io_B_Valid_63_45 <= _zz_io_B_Valid_63_44;
    _zz_io_B_Valid_63_46 <= _zz_io_B_Valid_63_45;
    _zz_io_B_Valid_63_47 <= _zz_io_B_Valid_63_46;
    _zz_io_B_Valid_63_48 <= _zz_io_B_Valid_63_47;
    _zz_io_B_Valid_63_49 <= _zz_io_B_Valid_63_48;
    _zz_io_B_Valid_63_50 <= _zz_io_B_Valid_63_49;
    _zz_io_B_Valid_63_51 <= _zz_io_B_Valid_63_50;
    _zz_io_B_Valid_63_52 <= _zz_io_B_Valid_63_51;
    _zz_io_B_Valid_63_53 <= _zz_io_B_Valid_63_52;
    _zz_io_B_Valid_63_54 <= _zz_io_B_Valid_63_53;
    _zz_io_B_Valid_63_55 <= _zz_io_B_Valid_63_54;
    _zz_io_B_Valid_63_56 <= _zz_io_B_Valid_63_55;
    _zz_io_B_Valid_63_57 <= _zz_io_B_Valid_63_56;
    _zz_io_B_Valid_63_58 <= _zz_io_B_Valid_63_57;
    _zz_io_B_Valid_63_59 <= _zz_io_B_Valid_63_58;
    _zz_io_B_Valid_63_60 <= _zz_io_B_Valid_63_59;
    _zz_io_B_Valid_63_61 <= _zz_io_B_Valid_63_60;
    _zz_io_B_Valid_63_62 <= _zz_io_B_Valid_63_61;
    toplevel_SubModule_WeightCache_Weight_Cached_delay_1 <= SubModule_WeightCache_Weight_Cached;
    toplevel_SubModule_WeightCache_Weight_Cached_delay_2 <= toplevel_SubModule_WeightCache_Weight_Cached_delay_1;
    toplevel_SubModule_WeightCache_Weight_Cached_delay_3 <= toplevel_SubModule_WeightCache_Weight_Cached_delay_2;
    _zz_start <= ((Fsm_nextState & TopCtrl_Enum_WEIGHT_CACHE) != 6'b000000);
    _zz_start_1 <= _zz_start;
    _zz_start_2 <= _zz_start_1;
  end


endmodule

module ConvArrangeV3 (
  input      [7:0]    sData_0,
  input      [7:0]    sData_1,
  input      [7:0]    sData_2,
  input      [7:0]    sData_3,
  input      [7:0]    sData_4,
  input      [7:0]    sData_5,
  input      [7:0]    sData_6,
  input      [7:0]    sData_7,
  output              sReady,
  input      [7:0]    sValid,
  input      [11:0]   MatrixCol,
  input      [19:0]   MatrixRow,
  input      [9:0]    OutChannel,
  input      [15:0]   OutFeatureSize,
  output reg          mData_valid,
  input               mData_ready,
  output reg [63:0]   mData_payload,
  output              mLast,
  output              LayerEnd,
  input               start,
  input               SwitchConv,
  input               clk,
  input               reset
);
  localparam CONVOUTPUT_ENUM_IDLE = 4'd1;
  localparam CONVOUTPUT_ENUM_INIT = 4'd2;
  localparam CONVOUTPUT_ENUM_DATA_ARRANGEMENT = 4'd4;
  localparam CONVOUTPUT_ENUM_WAIT_END = 4'd8;

  wire                ConvCtrl_ResetCnt;
  wire                ConvCtrl_InData_Cnt_En;
  wire                ConvCtrl_OutData_Cnt_En;
  wire                GemmCtrl_ResetCnt;
  wire                GemmCtrl_InData_Cnt_En;
  wire                GemmCtrl_OutData_Cnt_En;
  reg                 streamFifo_io_pop_ready;
  wire                axisDataConverter_8_inStream_valid;
  reg                 streamFifo_1_io_pop_ready;
  wire                axisDataConverter_9_inStream_valid;
  reg                 streamFifo_2_io_pop_ready;
  wire                axisDataConverter_10_inStream_valid;
  reg                 streamFifo_3_io_pop_ready;
  wire                axisDataConverter_11_inStream_valid;
  reg                 streamFifo_4_io_pop_ready;
  wire                axisDataConverter_12_inStream_valid;
  reg                 streamFifo_5_io_pop_ready;
  wire                axisDataConverter_13_inStream_valid;
  reg                 streamFifo_6_io_pop_ready;
  wire                axisDataConverter_14_inStream_valid;
  reg                 streamFifo_7_io_pop_ready;
  wire                axisDataConverter_15_inStream_valid;
  wire                ConvCtrl_Fsm_LayerEnd;
  wire                ConvCtrl_Fsm_Data_AllOut;
  wire                ConvCtrl_OutSwitch_Rotate;
  wire                ConvCtrl_OutSwitch_Reset;
  wire                GemmCtrl_Fsm_LayerEnd;
  wire                GemmCtrl_Fsm_Data_AllOut;
  wire                GemmCtrl_OutSwitch_Rotate;
  wire                streamFifo_io_push_ready;
  wire                streamFifo_io_pop_valid;
  wire       [63:0]   streamFifo_io_pop_payload;
  wire       [9:0]    streamFifo_io_occupancy;
  wire       [9:0]    streamFifo_io_availability;
  wire                axisDataConverter_8_inStream_ready;
  wire                axisDataConverter_8_outStream_valid;
  wire       [63:0]   axisDataConverter_8_outStream_payload;
  wire                streamFifo_1_io_push_ready;
  wire                streamFifo_1_io_pop_valid;
  wire       [63:0]   streamFifo_1_io_pop_payload;
  wire       [9:0]    streamFifo_1_io_occupancy;
  wire       [9:0]    streamFifo_1_io_availability;
  wire                axisDataConverter_9_inStream_ready;
  wire                axisDataConverter_9_outStream_valid;
  wire       [63:0]   axisDataConverter_9_outStream_payload;
  wire                streamFifo_2_io_push_ready;
  wire                streamFifo_2_io_pop_valid;
  wire       [63:0]   streamFifo_2_io_pop_payload;
  wire       [9:0]    streamFifo_2_io_occupancy;
  wire       [9:0]    streamFifo_2_io_availability;
  wire                axisDataConverter_10_inStream_ready;
  wire                axisDataConverter_10_outStream_valid;
  wire       [63:0]   axisDataConverter_10_outStream_payload;
  wire                streamFifo_3_io_push_ready;
  wire                streamFifo_3_io_pop_valid;
  wire       [63:0]   streamFifo_3_io_pop_payload;
  wire       [9:0]    streamFifo_3_io_occupancy;
  wire       [9:0]    streamFifo_3_io_availability;
  wire                axisDataConverter_11_inStream_ready;
  wire                axisDataConverter_11_outStream_valid;
  wire       [63:0]   axisDataConverter_11_outStream_payload;
  wire                streamFifo_4_io_push_ready;
  wire                streamFifo_4_io_pop_valid;
  wire       [63:0]   streamFifo_4_io_pop_payload;
  wire       [9:0]    streamFifo_4_io_occupancy;
  wire       [9:0]    streamFifo_4_io_availability;
  wire                axisDataConverter_12_inStream_ready;
  wire                axisDataConverter_12_outStream_valid;
  wire       [63:0]   axisDataConverter_12_outStream_payload;
  wire                streamFifo_5_io_push_ready;
  wire                streamFifo_5_io_pop_valid;
  wire       [63:0]   streamFifo_5_io_pop_payload;
  wire       [9:0]    streamFifo_5_io_occupancy;
  wire       [9:0]    streamFifo_5_io_availability;
  wire                axisDataConverter_13_inStream_ready;
  wire                axisDataConverter_13_outStream_valid;
  wire       [63:0]   axisDataConverter_13_outStream_payload;
  wire                streamFifo_6_io_push_ready;
  wire                streamFifo_6_io_pop_valid;
  wire       [63:0]   streamFifo_6_io_pop_payload;
  wire       [9:0]    streamFifo_6_io_occupancy;
  wire       [9:0]    streamFifo_6_io_availability;
  wire                axisDataConverter_14_inStream_ready;
  wire                axisDataConverter_14_outStream_valid;
  wire       [63:0]   axisDataConverter_14_outStream_payload;
  wire                streamFifo_7_io_push_ready;
  wire                streamFifo_7_io_pop_valid;
  wire       [63:0]   streamFifo_7_io_pop_payload;
  wire       [9:0]    streamFifo_7_io_occupancy;
  wire       [9:0]    streamFifo_7_io_availability;
  wire                axisDataConverter_15_inStream_ready;
  wire                axisDataConverter_15_outStream_valid;
  wire       [63:0]   axisDataConverter_15_outStream_payload;
  wire       [0:0]    _zz_when_SA3D_DataArrange_l131;
  wire       [0:0]    _zz_when_SA3D_DataArrange_l131_1;
  wire       [0:0]    _zz_when_SA3D_DataArrange_l131_2;
  wire       [0:0]    _zz_when_SA3D_DataArrange_l131_3;
  wire       [0:0]    _zz_when_SA3D_DataArrange_l131_4;
  wire       [0:0]    _zz_when_SA3D_DataArrange_l131_5;
  wire       [0:0]    _zz_when_SA3D_DataArrange_l131_6;
  wire       [0:0]    _zz_when_SA3D_DataArrange_l131_7;
  reg        [3:0]    Fsm_currentState;
  reg        [3:0]    Fsm_nextState;
  wire                Fsm_Inited;
  wire                Fsm_LayerEnd;
  wire                Fsm_Data_AllOut;
  wire                mData_fire;
  wire                mData_fire_1;
  wire                when_WaCounter_l40;
  reg        [2:0]    Init_Cnt_count;
  wire                Init_Cnt_valid;
  reg        [7:0]    OutSwitch;
  wire                when_SA3D_DataArrange_l108;
  wire                when_SA3D_DataArrange_l112;
  wire                when_SA3D_DataArrange_l131;
  wire                when_SA3D_DataArrange_l131_1;
  wire                when_SA3D_DataArrange_l131_2;
  wire                when_SA3D_DataArrange_l131_3;
  wire                when_SA3D_DataArrange_l131_4;
  wire                when_SA3D_DataArrange_l131_5;
  wire                when_SA3D_DataArrange_l131_6;
  wire                when_SA3D_DataArrange_l131_7;
  `ifndef SYNTHESIS
  reg [127:0] Fsm_currentState_string;
  reg [127:0] Fsm_nextState_string;
  `endif


  assign _zz_when_SA3D_DataArrange_l131 = OutSwitch[0 : 0];
  assign _zz_when_SA3D_DataArrange_l131_1 = OutSwitch[1 : 1];
  assign _zz_when_SA3D_DataArrange_l131_2 = OutSwitch[2 : 2];
  assign _zz_when_SA3D_DataArrange_l131_3 = OutSwitch[3 : 3];
  assign _zz_when_SA3D_DataArrange_l131_4 = OutSwitch[4 : 4];
  assign _zz_when_SA3D_DataArrange_l131_5 = OutSwitch[5 : 5];
  assign _zz_when_SA3D_DataArrange_l131_6 = OutSwitch[6 : 6];
  assign _zz_when_SA3D_DataArrange_l131_7 = OutSwitch[7 : 7];
  ConvOutput_Ctrl ConvCtrl (
    .ResetCnt         (ConvCtrl_ResetCnt        ), //i
    .InData_Cnt_En    (ConvCtrl_InData_Cnt_En   ), //i
    .OutData_Cnt_En   (ConvCtrl_OutData_Cnt_En  ), //i
    .OutChannel       (OutChannel[9:0]          ), //i
    .OutFeatureSize   (OutFeatureSize[15:0]     ), //i
    .Fsm_LayerEnd     (ConvCtrl_Fsm_LayerEnd    ), //o
    .Fsm_Data_AllOut  (ConvCtrl_Fsm_Data_AllOut ), //o
    .OutSwitch_Rotate (ConvCtrl_OutSwitch_Rotate), //o
    .OutSwitch_Reset  (ConvCtrl_OutSwitch_Reset ), //o
    .clk              (clk                      ), //i
    .reset            (reset                    )  //i
  );
  GemmOutput_Ctrl GemmCtrl (
    .ResetCnt         (GemmCtrl_ResetCnt        ), //i
    .InData_Cnt_En    (GemmCtrl_InData_Cnt_En   ), //i
    .OutData_Cnt_En   (GemmCtrl_OutData_Cnt_En  ), //i
    .MatrixCol        (MatrixCol[11:0]          ), //i
    .MatrixRow        (MatrixRow[19:0]          ), //i
    .Fsm_LayerEnd     (GemmCtrl_Fsm_LayerEnd    ), //o
    .Fsm_Data_AllOut  (GemmCtrl_Fsm_Data_AllOut ), //o
    .OutSwitch_Rotate (GemmCtrl_OutSwitch_Rotate), //o
    .clk              (clk                      ), //i
    .reset            (reset                    )  //i
  );
  ConvOutput_Fifo streamFifo (
    .io_push_valid   (axisDataConverter_8_outStream_valid        ), //i
    .io_push_ready   (streamFifo_io_push_ready                   ), //o
    .io_push_payload (axisDataConverter_8_outStream_payload[63:0]), //i
    .io_pop_valid    (streamFifo_io_pop_valid                    ), //o
    .io_pop_ready    (streamFifo_io_pop_ready                    ), //i
    .io_pop_payload  (streamFifo_io_pop_payload[63:0]            ), //o
    .io_flush        (1'b0                                       ), //i
    .io_occupancy    (streamFifo_io_occupancy[9:0]               ), //o
    .io_availability (streamFifo_io_availability[9:0]            ), //o
    .clk             (clk                                        ), //i
    .reset           (reset                                      )  //i
  );
  ConvOutput_Converter axisDataConverter_8 (
    .inStream_valid    (axisDataConverter_8_inStream_valid         ), //i
    .inStream_ready    (axisDataConverter_8_inStream_ready         ), //o
    .inStream_payload  (sData_0[7:0]                               ), //i
    .outStream_valid   (axisDataConverter_8_outStream_valid        ), //o
    .outStream_ready   (streamFifo_io_push_ready                   ), //i
    .outStream_payload (axisDataConverter_8_outStream_payload[63:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  ConvOutput_Fifo streamFifo_1 (
    .io_push_valid   (axisDataConverter_9_outStream_valid        ), //i
    .io_push_ready   (streamFifo_1_io_push_ready                 ), //o
    .io_push_payload (axisDataConverter_9_outStream_payload[63:0]), //i
    .io_pop_valid    (streamFifo_1_io_pop_valid                  ), //o
    .io_pop_ready    (streamFifo_1_io_pop_ready                  ), //i
    .io_pop_payload  (streamFifo_1_io_pop_payload[63:0]          ), //o
    .io_flush        (1'b0                                       ), //i
    .io_occupancy    (streamFifo_1_io_occupancy[9:0]             ), //o
    .io_availability (streamFifo_1_io_availability[9:0]          ), //o
    .clk             (clk                                        ), //i
    .reset           (reset                                      )  //i
  );
  ConvOutput_Converter axisDataConverter_9 (
    .inStream_valid    (axisDataConverter_9_inStream_valid         ), //i
    .inStream_ready    (axisDataConverter_9_inStream_ready         ), //o
    .inStream_payload  (sData_1[7:0]                               ), //i
    .outStream_valid   (axisDataConverter_9_outStream_valid        ), //o
    .outStream_ready   (streamFifo_1_io_push_ready                 ), //i
    .outStream_payload (axisDataConverter_9_outStream_payload[63:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  ConvOutput_Fifo streamFifo_2 (
    .io_push_valid   (axisDataConverter_10_outStream_valid        ), //i
    .io_push_ready   (streamFifo_2_io_push_ready                  ), //o
    .io_push_payload (axisDataConverter_10_outStream_payload[63:0]), //i
    .io_pop_valid    (streamFifo_2_io_pop_valid                   ), //o
    .io_pop_ready    (streamFifo_2_io_pop_ready                   ), //i
    .io_pop_payload  (streamFifo_2_io_pop_payload[63:0]           ), //o
    .io_flush        (1'b0                                        ), //i
    .io_occupancy    (streamFifo_2_io_occupancy[9:0]              ), //o
    .io_availability (streamFifo_2_io_availability[9:0]           ), //o
    .clk             (clk                                         ), //i
    .reset           (reset                                       )  //i
  );
  ConvOutput_Converter axisDataConverter_10 (
    .inStream_valid    (axisDataConverter_10_inStream_valid         ), //i
    .inStream_ready    (axisDataConverter_10_inStream_ready         ), //o
    .inStream_payload  (sData_2[7:0]                                ), //i
    .outStream_valid   (axisDataConverter_10_outStream_valid        ), //o
    .outStream_ready   (streamFifo_2_io_push_ready                  ), //i
    .outStream_payload (axisDataConverter_10_outStream_payload[63:0]), //o
    .clk               (clk                                         ), //i
    .reset             (reset                                       )  //i
  );
  ConvOutput_Fifo streamFifo_3 (
    .io_push_valid   (axisDataConverter_11_outStream_valid        ), //i
    .io_push_ready   (streamFifo_3_io_push_ready                  ), //o
    .io_push_payload (axisDataConverter_11_outStream_payload[63:0]), //i
    .io_pop_valid    (streamFifo_3_io_pop_valid                   ), //o
    .io_pop_ready    (streamFifo_3_io_pop_ready                   ), //i
    .io_pop_payload  (streamFifo_3_io_pop_payload[63:0]           ), //o
    .io_flush        (1'b0                                        ), //i
    .io_occupancy    (streamFifo_3_io_occupancy[9:0]              ), //o
    .io_availability (streamFifo_3_io_availability[9:0]           ), //o
    .clk             (clk                                         ), //i
    .reset           (reset                                       )  //i
  );
  ConvOutput_Converter axisDataConverter_11 (
    .inStream_valid    (axisDataConverter_11_inStream_valid         ), //i
    .inStream_ready    (axisDataConverter_11_inStream_ready         ), //o
    .inStream_payload  (sData_3[7:0]                                ), //i
    .outStream_valid   (axisDataConverter_11_outStream_valid        ), //o
    .outStream_ready   (streamFifo_3_io_push_ready                  ), //i
    .outStream_payload (axisDataConverter_11_outStream_payload[63:0]), //o
    .clk               (clk                                         ), //i
    .reset             (reset                                       )  //i
  );
  ConvOutput_Fifo streamFifo_4 (
    .io_push_valid   (axisDataConverter_12_outStream_valid        ), //i
    .io_push_ready   (streamFifo_4_io_push_ready                  ), //o
    .io_push_payload (axisDataConverter_12_outStream_payload[63:0]), //i
    .io_pop_valid    (streamFifo_4_io_pop_valid                   ), //o
    .io_pop_ready    (streamFifo_4_io_pop_ready                   ), //i
    .io_pop_payload  (streamFifo_4_io_pop_payload[63:0]           ), //o
    .io_flush        (1'b0                                        ), //i
    .io_occupancy    (streamFifo_4_io_occupancy[9:0]              ), //o
    .io_availability (streamFifo_4_io_availability[9:0]           ), //o
    .clk             (clk                                         ), //i
    .reset           (reset                                       )  //i
  );
  ConvOutput_Converter axisDataConverter_12 (
    .inStream_valid    (axisDataConverter_12_inStream_valid         ), //i
    .inStream_ready    (axisDataConverter_12_inStream_ready         ), //o
    .inStream_payload  (sData_4[7:0]                                ), //i
    .outStream_valid   (axisDataConverter_12_outStream_valid        ), //o
    .outStream_ready   (streamFifo_4_io_push_ready                  ), //i
    .outStream_payload (axisDataConverter_12_outStream_payload[63:0]), //o
    .clk               (clk                                         ), //i
    .reset             (reset                                       )  //i
  );
  ConvOutput_Fifo streamFifo_5 (
    .io_push_valid   (axisDataConverter_13_outStream_valid        ), //i
    .io_push_ready   (streamFifo_5_io_push_ready                  ), //o
    .io_push_payload (axisDataConverter_13_outStream_payload[63:0]), //i
    .io_pop_valid    (streamFifo_5_io_pop_valid                   ), //o
    .io_pop_ready    (streamFifo_5_io_pop_ready                   ), //i
    .io_pop_payload  (streamFifo_5_io_pop_payload[63:0]           ), //o
    .io_flush        (1'b0                                        ), //i
    .io_occupancy    (streamFifo_5_io_occupancy[9:0]              ), //o
    .io_availability (streamFifo_5_io_availability[9:0]           ), //o
    .clk             (clk                                         ), //i
    .reset           (reset                                       )  //i
  );
  ConvOutput_Converter axisDataConverter_13 (
    .inStream_valid    (axisDataConverter_13_inStream_valid         ), //i
    .inStream_ready    (axisDataConverter_13_inStream_ready         ), //o
    .inStream_payload  (sData_5[7:0]                                ), //i
    .outStream_valid   (axisDataConverter_13_outStream_valid        ), //o
    .outStream_ready   (streamFifo_5_io_push_ready                  ), //i
    .outStream_payload (axisDataConverter_13_outStream_payload[63:0]), //o
    .clk               (clk                                         ), //i
    .reset             (reset                                       )  //i
  );
  ConvOutput_Fifo streamFifo_6 (
    .io_push_valid   (axisDataConverter_14_outStream_valid        ), //i
    .io_push_ready   (streamFifo_6_io_push_ready                  ), //o
    .io_push_payload (axisDataConverter_14_outStream_payload[63:0]), //i
    .io_pop_valid    (streamFifo_6_io_pop_valid                   ), //o
    .io_pop_ready    (streamFifo_6_io_pop_ready                   ), //i
    .io_pop_payload  (streamFifo_6_io_pop_payload[63:0]           ), //o
    .io_flush        (1'b0                                        ), //i
    .io_occupancy    (streamFifo_6_io_occupancy[9:0]              ), //o
    .io_availability (streamFifo_6_io_availability[9:0]           ), //o
    .clk             (clk                                         ), //i
    .reset           (reset                                       )  //i
  );
  ConvOutput_Converter axisDataConverter_14 (
    .inStream_valid    (axisDataConverter_14_inStream_valid         ), //i
    .inStream_ready    (axisDataConverter_14_inStream_ready         ), //o
    .inStream_payload  (sData_6[7:0]                                ), //i
    .outStream_valid   (axisDataConverter_14_outStream_valid        ), //o
    .outStream_ready   (streamFifo_6_io_push_ready                  ), //i
    .outStream_payload (axisDataConverter_14_outStream_payload[63:0]), //o
    .clk               (clk                                         ), //i
    .reset             (reset                                       )  //i
  );
  ConvOutput_Fifo streamFifo_7 (
    .io_push_valid   (axisDataConverter_15_outStream_valid        ), //i
    .io_push_ready   (streamFifo_7_io_push_ready                  ), //o
    .io_push_payload (axisDataConverter_15_outStream_payload[63:0]), //i
    .io_pop_valid    (streamFifo_7_io_pop_valid                   ), //o
    .io_pop_ready    (streamFifo_7_io_pop_ready                   ), //i
    .io_pop_payload  (streamFifo_7_io_pop_payload[63:0]           ), //o
    .io_flush        (1'b0                                        ), //i
    .io_occupancy    (streamFifo_7_io_occupancy[9:0]              ), //o
    .io_availability (streamFifo_7_io_availability[9:0]           ), //o
    .clk             (clk                                         ), //i
    .reset           (reset                                       )  //i
  );
  ConvOutput_Converter axisDataConverter_15 (
    .inStream_valid    (axisDataConverter_15_inStream_valid         ), //i
    .inStream_ready    (axisDataConverter_15_inStream_ready         ), //o
    .inStream_payload  (sData_7[7:0]                                ), //i
    .outStream_valid   (axisDataConverter_15_outStream_valid        ), //o
    .outStream_ready   (streamFifo_7_io_push_ready                  ), //i
    .outStream_payload (axisDataConverter_15_outStream_payload[63:0]), //o
    .clk               (clk                                         ), //i
    .reset             (reset                                       )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      CONVOUTPUT_ENUM_IDLE : Fsm_currentState_string = "IDLE            ";
      CONVOUTPUT_ENUM_INIT : Fsm_currentState_string = "INIT            ";
      CONVOUTPUT_ENUM_DATA_ARRANGEMENT : Fsm_currentState_string = "DATA_ARRANGEMENT";
      CONVOUTPUT_ENUM_WAIT_END : Fsm_currentState_string = "WAIT_END        ";
      default : Fsm_currentState_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      CONVOUTPUT_ENUM_IDLE : Fsm_nextState_string = "IDLE            ";
      CONVOUTPUT_ENUM_INIT : Fsm_nextState_string = "INIT            ";
      CONVOUTPUT_ENUM_DATA_ARRANGEMENT : Fsm_nextState_string = "DATA_ARRANGEMENT";
      CONVOUTPUT_ENUM_WAIT_END : Fsm_nextState_string = "WAIT_END        ";
      default : Fsm_nextState_string = "????????????????";
    endcase
  end
  `endif

  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & CONVOUTPUT_ENUM_IDLE) == CONVOUTPUT_ENUM_IDLE) : begin
        if(start) begin
          Fsm_nextState = CONVOUTPUT_ENUM_INIT;
        end else begin
          Fsm_nextState = CONVOUTPUT_ENUM_IDLE;
        end
      end
      (((Fsm_currentState) & CONVOUTPUT_ENUM_INIT) == CONVOUTPUT_ENUM_INIT) : begin
        if(Fsm_Inited) begin
          Fsm_nextState = CONVOUTPUT_ENUM_DATA_ARRANGEMENT;
        end else begin
          Fsm_nextState = CONVOUTPUT_ENUM_INIT;
        end
      end
      (((Fsm_currentState) & CONVOUTPUT_ENUM_DATA_ARRANGEMENT) == CONVOUTPUT_ENUM_DATA_ARRANGEMENT) : begin
        if(Fsm_LayerEnd) begin
          Fsm_nextState = CONVOUTPUT_ENUM_WAIT_END;
        end else begin
          Fsm_nextState = CONVOUTPUT_ENUM_DATA_ARRANGEMENT;
        end
      end
      default : begin
        if(Fsm_Data_AllOut) begin
          Fsm_nextState = CONVOUTPUT_ENUM_IDLE;
        end else begin
          Fsm_nextState = CONVOUTPUT_ENUM_WAIT_END;
        end
      end
    endcase
  end

  assign ConvCtrl_ResetCnt = ((Fsm_currentState & CONVOUTPUT_ENUM_INIT) != 4'b0000);
  assign ConvCtrl_InData_Cnt_En = ((sReady && sValid[0]) && SwitchConv);
  assign mData_fire = (mData_valid && mData_ready);
  assign ConvCtrl_OutData_Cnt_En = (mData_fire && SwitchConv);
  assign GemmCtrl_ResetCnt = ((Fsm_currentState & CONVOUTPUT_ENUM_INIT) != 4'b0000);
  assign GemmCtrl_InData_Cnt_En = ((sReady && sValid[0]) && (! SwitchConv));
  assign mData_fire_1 = (mData_valid && mData_ready);
  assign GemmCtrl_OutData_Cnt_En = (mData_fire_1 && (! SwitchConv));
  assign when_WaCounter_l40 = ((Fsm_currentState & CONVOUTPUT_ENUM_INIT) != 4'b0000);
  assign Init_Cnt_valid = ((Init_Cnt_count == 3'b101) && when_WaCounter_l40);
  assign Fsm_Inited = Init_Cnt_valid;
  assign Fsm_LayerEnd = ((ConvCtrl_Fsm_LayerEnd && SwitchConv) || (GemmCtrl_Fsm_LayerEnd && (! SwitchConv)));
  assign Fsm_Data_AllOut = ((ConvCtrl_Fsm_Data_AllOut && SwitchConv) || (GemmCtrl_Fsm_Data_AllOut && (! SwitchConv)));
  always @(*) begin
    mData_payload = 64'h0;
    if(when_SA3D_DataArrange_l131) begin
      mData_payload = streamFifo_io_pop_payload;
    end
    if(when_SA3D_DataArrange_l131_1) begin
      mData_payload = streamFifo_1_io_pop_payload;
    end
    if(when_SA3D_DataArrange_l131_2) begin
      mData_payload = streamFifo_2_io_pop_payload;
    end
    if(when_SA3D_DataArrange_l131_3) begin
      mData_payload = streamFifo_3_io_pop_payload;
    end
    if(when_SA3D_DataArrange_l131_4) begin
      mData_payload = streamFifo_4_io_pop_payload;
    end
    if(when_SA3D_DataArrange_l131_5) begin
      mData_payload = streamFifo_5_io_pop_payload;
    end
    if(when_SA3D_DataArrange_l131_6) begin
      mData_payload = streamFifo_6_io_pop_payload;
    end
    if(when_SA3D_DataArrange_l131_7) begin
      mData_payload = streamFifo_7_io_pop_payload;
    end
  end

  always @(*) begin
    mData_valid = 1'b0;
    if(when_SA3D_DataArrange_l131) begin
      mData_valid = streamFifo_io_pop_valid;
    end
    if(when_SA3D_DataArrange_l131_1) begin
      mData_valid = streamFifo_1_io_pop_valid;
    end
    if(when_SA3D_DataArrange_l131_2) begin
      mData_valid = streamFifo_2_io_pop_valid;
    end
    if(when_SA3D_DataArrange_l131_3) begin
      mData_valid = streamFifo_3_io_pop_valid;
    end
    if(when_SA3D_DataArrange_l131_4) begin
      mData_valid = streamFifo_4_io_pop_valid;
    end
    if(when_SA3D_DataArrange_l131_5) begin
      mData_valid = streamFifo_5_io_pop_valid;
    end
    if(when_SA3D_DataArrange_l131_6) begin
      mData_valid = streamFifo_6_io_pop_valid;
    end
    if(when_SA3D_DataArrange_l131_7) begin
      mData_valid = streamFifo_7_io_pop_valid;
    end
  end

  assign when_SA3D_DataArrange_l108 = ((Fsm_currentState & CONVOUTPUT_ENUM_INIT) != 4'b0000);
  assign when_SA3D_DataArrange_l112 = (ConvCtrl_OutSwitch_Rotate || GemmCtrl_OutSwitch_Rotate);
  assign sReady = (axisDataConverter_8_inStream_ready && ((Fsm_currentState & CONVOUTPUT_ENUM_DATA_ARRANGEMENT) != 4'b0000));
  assign axisDataConverter_8_inStream_valid = (sValid[0] && ((Fsm_currentState & CONVOUTPUT_ENUM_DATA_ARRANGEMENT) != 4'b0000));
  always @(*) begin
    streamFifo_io_pop_ready = 1'b0;
    if(when_SA3D_DataArrange_l131) begin
      streamFifo_io_pop_ready = mData_ready;
    end
  end

  assign when_SA3D_DataArrange_l131 = _zz_when_SA3D_DataArrange_l131[0];
  assign axisDataConverter_9_inStream_valid = (sValid[1] && ((Fsm_currentState & CONVOUTPUT_ENUM_DATA_ARRANGEMENT) != 4'b0000));
  always @(*) begin
    streamFifo_1_io_pop_ready = 1'b0;
    if(when_SA3D_DataArrange_l131_1) begin
      streamFifo_1_io_pop_ready = mData_ready;
    end
  end

  assign when_SA3D_DataArrange_l131_1 = _zz_when_SA3D_DataArrange_l131_1[0];
  assign axisDataConverter_10_inStream_valid = (sValid[2] && ((Fsm_currentState & CONVOUTPUT_ENUM_DATA_ARRANGEMENT) != 4'b0000));
  always @(*) begin
    streamFifo_2_io_pop_ready = 1'b0;
    if(when_SA3D_DataArrange_l131_2) begin
      streamFifo_2_io_pop_ready = mData_ready;
    end
  end

  assign when_SA3D_DataArrange_l131_2 = _zz_when_SA3D_DataArrange_l131_2[0];
  assign axisDataConverter_11_inStream_valid = (sValid[3] && ((Fsm_currentState & CONVOUTPUT_ENUM_DATA_ARRANGEMENT) != 4'b0000));
  always @(*) begin
    streamFifo_3_io_pop_ready = 1'b0;
    if(when_SA3D_DataArrange_l131_3) begin
      streamFifo_3_io_pop_ready = mData_ready;
    end
  end

  assign when_SA3D_DataArrange_l131_3 = _zz_when_SA3D_DataArrange_l131_3[0];
  assign axisDataConverter_12_inStream_valid = (sValid[4] && ((Fsm_currentState & CONVOUTPUT_ENUM_DATA_ARRANGEMENT) != 4'b0000));
  always @(*) begin
    streamFifo_4_io_pop_ready = 1'b0;
    if(when_SA3D_DataArrange_l131_4) begin
      streamFifo_4_io_pop_ready = mData_ready;
    end
  end

  assign when_SA3D_DataArrange_l131_4 = _zz_when_SA3D_DataArrange_l131_4[0];
  assign axisDataConverter_13_inStream_valid = (sValid[5] && ((Fsm_currentState & CONVOUTPUT_ENUM_DATA_ARRANGEMENT) != 4'b0000));
  always @(*) begin
    streamFifo_5_io_pop_ready = 1'b0;
    if(when_SA3D_DataArrange_l131_5) begin
      streamFifo_5_io_pop_ready = mData_ready;
    end
  end

  assign when_SA3D_DataArrange_l131_5 = _zz_when_SA3D_DataArrange_l131_5[0];
  assign axisDataConverter_14_inStream_valid = (sValid[6] && ((Fsm_currentState & CONVOUTPUT_ENUM_DATA_ARRANGEMENT) != 4'b0000));
  always @(*) begin
    streamFifo_6_io_pop_ready = 1'b0;
    if(when_SA3D_DataArrange_l131_6) begin
      streamFifo_6_io_pop_ready = mData_ready;
    end
  end

  assign when_SA3D_DataArrange_l131_6 = _zz_when_SA3D_DataArrange_l131_6[0];
  assign axisDataConverter_15_inStream_valid = (sValid[7] && ((Fsm_currentState & CONVOUTPUT_ENUM_DATA_ARRANGEMENT) != 4'b0000));
  always @(*) begin
    streamFifo_7_io_pop_ready = 1'b0;
    if(when_SA3D_DataArrange_l131_7) begin
      streamFifo_7_io_pop_ready = mData_ready;
    end
  end

  assign when_SA3D_DataArrange_l131_7 = _zz_when_SA3D_DataArrange_l131_7[0];
  assign mLast = Fsm_Data_AllOut;
  assign LayerEnd = Fsm_Data_AllOut;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= CONVOUTPUT_ENUM_IDLE;
      Init_Cnt_count <= 3'b000;
      OutSwitch <= 8'h01;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l40) begin
        if(Init_Cnt_valid) begin
          Init_Cnt_count <= 3'b000;
        end else begin
          Init_Cnt_count <= (Init_Cnt_count + 3'b001);
        end
      end
      if(when_SA3D_DataArrange_l108) begin
        OutSwitch <= 8'h01;
      end else begin
        if(ConvCtrl_OutSwitch_Reset) begin
          OutSwitch <= 8'h01;
        end else begin
          if(when_SA3D_DataArrange_l112) begin
            OutSwitch <= {OutSwitch[6 : 0],OutSwitch[7 : 7]};
          end
        end
      end
    end
  end


endmodule

module WeightCache_Stream (
  input      [63:0]   s_axis_s2mm_tdata,
  input      [7:0]    s_axis_s2mm_tkeep,
  input               s_axis_s2mm_tlast,
  output              s_axis_s2mm_tready,
  input               s_axis_s2mm_tvalid,
  input               start,
  input      [15:0]   Matrix_Row,
  input      [15:0]   Matrix_Col,
  output     [7:0]    mData_0,
  output     [7:0]    mData_1,
  output     [7:0]    mData_2,
  output     [7:0]    mData_3,
  output     [7:0]    mData_4,
  output     [7:0]    mData_5,
  output     [7:0]    mData_6,
  output     [7:0]    mData_7,
  output     [7:0]    mData_8,
  output     [7:0]    mData_9,
  output     [7:0]    mData_10,
  output     [7:0]    mData_11,
  output     [7:0]    mData_12,
  output     [7:0]    mData_13,
  output     [7:0]    mData_14,
  output     [7:0]    mData_15,
  output     [7:0]    mData_16,
  output     [7:0]    mData_17,
  output     [7:0]    mData_18,
  output     [7:0]    mData_19,
  output     [7:0]    mData_20,
  output     [7:0]    mData_21,
  output     [7:0]    mData_22,
  output     [7:0]    mData_23,
  output     [7:0]    mData_24,
  output     [7:0]    mData_25,
  output     [7:0]    mData_26,
  output     [7:0]    mData_27,
  output     [7:0]    mData_28,
  output     [7:0]    mData_29,
  output     [7:0]    mData_30,
  output     [7:0]    mData_31,
  output     [7:0]    mData_32,
  output     [7:0]    mData_33,
  output     [7:0]    mData_34,
  output     [7:0]    mData_35,
  output     [7:0]    mData_36,
  output     [7:0]    mData_37,
  output     [7:0]    mData_38,
  output     [7:0]    mData_39,
  output     [7:0]    mData_40,
  output     [7:0]    mData_41,
  output     [7:0]    mData_42,
  output     [7:0]    mData_43,
  output     [7:0]    mData_44,
  output     [7:0]    mData_45,
  output     [7:0]    mData_46,
  output     [7:0]    mData_47,
  output     [7:0]    mData_48,
  output     [7:0]    mData_49,
  output     [7:0]    mData_50,
  output     [7:0]    mData_51,
  output     [7:0]    mData_52,
  output     [7:0]    mData_53,
  output     [7:0]    mData_54,
  output     [7:0]    mData_55,
  output     [7:0]    mData_56,
  output     [7:0]    mData_57,
  output     [7:0]    mData_58,
  output     [7:0]    mData_59,
  output     [7:0]    mData_60,
  output     [7:0]    mData_61,
  output     [7:0]    mData_62,
  output     [7:0]    mData_63,
  input               Raddr_Valid,
  output              Weight_Cached,
  input               LayerEnd,
  output     [63:0]   MatrixCol_Switch,
  input               clk,
  input               reset
);

  wire                WeightCache_sData_ready;
  wire       [7:0]    WeightCache_mData_0;
  wire       [7:0]    WeightCache_mData_1;
  wire       [7:0]    WeightCache_mData_2;
  wire       [7:0]    WeightCache_mData_3;
  wire       [7:0]    WeightCache_mData_4;
  wire       [7:0]    WeightCache_mData_5;
  wire       [7:0]    WeightCache_mData_6;
  wire       [7:0]    WeightCache_mData_7;
  wire       [7:0]    WeightCache_mData_8;
  wire       [7:0]    WeightCache_mData_9;
  wire       [7:0]    WeightCache_mData_10;
  wire       [7:0]    WeightCache_mData_11;
  wire       [7:0]    WeightCache_mData_12;
  wire       [7:0]    WeightCache_mData_13;
  wire       [7:0]    WeightCache_mData_14;
  wire       [7:0]    WeightCache_mData_15;
  wire       [7:0]    WeightCache_mData_16;
  wire       [7:0]    WeightCache_mData_17;
  wire       [7:0]    WeightCache_mData_18;
  wire       [7:0]    WeightCache_mData_19;
  wire       [7:0]    WeightCache_mData_20;
  wire       [7:0]    WeightCache_mData_21;
  wire       [7:0]    WeightCache_mData_22;
  wire       [7:0]    WeightCache_mData_23;
  wire       [7:0]    WeightCache_mData_24;
  wire       [7:0]    WeightCache_mData_25;
  wire       [7:0]    WeightCache_mData_26;
  wire       [7:0]    WeightCache_mData_27;
  wire       [7:0]    WeightCache_mData_28;
  wire       [7:0]    WeightCache_mData_29;
  wire       [7:0]    WeightCache_mData_30;
  wire       [7:0]    WeightCache_mData_31;
  wire       [7:0]    WeightCache_mData_32;
  wire       [7:0]    WeightCache_mData_33;
  wire       [7:0]    WeightCache_mData_34;
  wire       [7:0]    WeightCache_mData_35;
  wire       [7:0]    WeightCache_mData_36;
  wire       [7:0]    WeightCache_mData_37;
  wire       [7:0]    WeightCache_mData_38;
  wire       [7:0]    WeightCache_mData_39;
  wire       [7:0]    WeightCache_mData_40;
  wire       [7:0]    WeightCache_mData_41;
  wire       [7:0]    WeightCache_mData_42;
  wire       [7:0]    WeightCache_mData_43;
  wire       [7:0]    WeightCache_mData_44;
  wire       [7:0]    WeightCache_mData_45;
  wire       [7:0]    WeightCache_mData_46;
  wire       [7:0]    WeightCache_mData_47;
  wire       [7:0]    WeightCache_mData_48;
  wire       [7:0]    WeightCache_mData_49;
  wire       [7:0]    WeightCache_mData_50;
  wire       [7:0]    WeightCache_mData_51;
  wire       [7:0]    WeightCache_mData_52;
  wire       [7:0]    WeightCache_mData_53;
  wire       [7:0]    WeightCache_mData_54;
  wire       [7:0]    WeightCache_mData_55;
  wire       [7:0]    WeightCache_mData_56;
  wire       [7:0]    WeightCache_mData_57;
  wire       [7:0]    WeightCache_mData_58;
  wire       [7:0]    WeightCache_mData_59;
  wire       [7:0]    WeightCache_mData_60;
  wire       [7:0]    WeightCache_mData_61;
  wire       [7:0]    WeightCache_mData_62;
  wire       [7:0]    WeightCache_mData_63;
  wire                WeightCache_Weight_Cached;
  wire       [63:0]   WeightCache_MatrixCol_Switch;

  Weight_Cache WeightCache (
    .start            (start                             ), //i
    .sData_valid      (s_axis_s2mm_tvalid                ), //i
    .sData_ready      (WeightCache_sData_ready           ), //o
    .sData_payload    (s_axis_s2mm_tdata[63:0]           ), //i
    .Matrix_Row       (Matrix_Row[15:0]                  ), //i
    .Matrix_Col       (Matrix_Col[15:0]                  ), //i
    .mData_0          (WeightCache_mData_0[7:0]          ), //o
    .mData_1          (WeightCache_mData_1[7:0]          ), //o
    .mData_2          (WeightCache_mData_2[7:0]          ), //o
    .mData_3          (WeightCache_mData_3[7:0]          ), //o
    .mData_4          (WeightCache_mData_4[7:0]          ), //o
    .mData_5          (WeightCache_mData_5[7:0]          ), //o
    .mData_6          (WeightCache_mData_6[7:0]          ), //o
    .mData_7          (WeightCache_mData_7[7:0]          ), //o
    .mData_8          (WeightCache_mData_8[7:0]          ), //o
    .mData_9          (WeightCache_mData_9[7:0]          ), //o
    .mData_10         (WeightCache_mData_10[7:0]         ), //o
    .mData_11         (WeightCache_mData_11[7:0]         ), //o
    .mData_12         (WeightCache_mData_12[7:0]         ), //o
    .mData_13         (WeightCache_mData_13[7:0]         ), //o
    .mData_14         (WeightCache_mData_14[7:0]         ), //o
    .mData_15         (WeightCache_mData_15[7:0]         ), //o
    .mData_16         (WeightCache_mData_16[7:0]         ), //o
    .mData_17         (WeightCache_mData_17[7:0]         ), //o
    .mData_18         (WeightCache_mData_18[7:0]         ), //o
    .mData_19         (WeightCache_mData_19[7:0]         ), //o
    .mData_20         (WeightCache_mData_20[7:0]         ), //o
    .mData_21         (WeightCache_mData_21[7:0]         ), //o
    .mData_22         (WeightCache_mData_22[7:0]         ), //o
    .mData_23         (WeightCache_mData_23[7:0]         ), //o
    .mData_24         (WeightCache_mData_24[7:0]         ), //o
    .mData_25         (WeightCache_mData_25[7:0]         ), //o
    .mData_26         (WeightCache_mData_26[7:0]         ), //o
    .mData_27         (WeightCache_mData_27[7:0]         ), //o
    .mData_28         (WeightCache_mData_28[7:0]         ), //o
    .mData_29         (WeightCache_mData_29[7:0]         ), //o
    .mData_30         (WeightCache_mData_30[7:0]         ), //o
    .mData_31         (WeightCache_mData_31[7:0]         ), //o
    .mData_32         (WeightCache_mData_32[7:0]         ), //o
    .mData_33         (WeightCache_mData_33[7:0]         ), //o
    .mData_34         (WeightCache_mData_34[7:0]         ), //o
    .mData_35         (WeightCache_mData_35[7:0]         ), //o
    .mData_36         (WeightCache_mData_36[7:0]         ), //o
    .mData_37         (WeightCache_mData_37[7:0]         ), //o
    .mData_38         (WeightCache_mData_38[7:0]         ), //o
    .mData_39         (WeightCache_mData_39[7:0]         ), //o
    .mData_40         (WeightCache_mData_40[7:0]         ), //o
    .mData_41         (WeightCache_mData_41[7:0]         ), //o
    .mData_42         (WeightCache_mData_42[7:0]         ), //o
    .mData_43         (WeightCache_mData_43[7:0]         ), //o
    .mData_44         (WeightCache_mData_44[7:0]         ), //o
    .mData_45         (WeightCache_mData_45[7:0]         ), //o
    .mData_46         (WeightCache_mData_46[7:0]         ), //o
    .mData_47         (WeightCache_mData_47[7:0]         ), //o
    .mData_48         (WeightCache_mData_48[7:0]         ), //o
    .mData_49         (WeightCache_mData_49[7:0]         ), //o
    .mData_50         (WeightCache_mData_50[7:0]         ), //o
    .mData_51         (WeightCache_mData_51[7:0]         ), //o
    .mData_52         (WeightCache_mData_52[7:0]         ), //o
    .mData_53         (WeightCache_mData_53[7:0]         ), //o
    .mData_54         (WeightCache_mData_54[7:0]         ), //o
    .mData_55         (WeightCache_mData_55[7:0]         ), //o
    .mData_56         (WeightCache_mData_56[7:0]         ), //o
    .mData_57         (WeightCache_mData_57[7:0]         ), //o
    .mData_58         (WeightCache_mData_58[7:0]         ), //o
    .mData_59         (WeightCache_mData_59[7:0]         ), //o
    .mData_60         (WeightCache_mData_60[7:0]         ), //o
    .mData_61         (WeightCache_mData_61[7:0]         ), //o
    .mData_62         (WeightCache_mData_62[7:0]         ), //o
    .mData_63         (WeightCache_mData_63[7:0]         ), //o
    .Raddr_Valid      (Raddr_Valid                       ), //i
    .Weight_Cached    (WeightCache_Weight_Cached         ), //o
    .LayerEnd         (LayerEnd                          ), //i
    .MatrixCol_Switch (WeightCache_MatrixCol_Switch[63:0]), //o
    .clk              (clk                               ), //i
    .reset            (reset                             )  //i
  );
  assign mData_0 = WeightCache_mData_0;
  assign mData_1 = WeightCache_mData_1;
  assign mData_2 = WeightCache_mData_2;
  assign mData_3 = WeightCache_mData_3;
  assign mData_4 = WeightCache_mData_4;
  assign mData_5 = WeightCache_mData_5;
  assign mData_6 = WeightCache_mData_6;
  assign mData_7 = WeightCache_mData_7;
  assign mData_8 = WeightCache_mData_8;
  assign mData_9 = WeightCache_mData_9;
  assign mData_10 = WeightCache_mData_10;
  assign mData_11 = WeightCache_mData_11;
  assign mData_12 = WeightCache_mData_12;
  assign mData_13 = WeightCache_mData_13;
  assign mData_14 = WeightCache_mData_14;
  assign mData_15 = WeightCache_mData_15;
  assign mData_16 = WeightCache_mData_16;
  assign mData_17 = WeightCache_mData_17;
  assign mData_18 = WeightCache_mData_18;
  assign mData_19 = WeightCache_mData_19;
  assign mData_20 = WeightCache_mData_20;
  assign mData_21 = WeightCache_mData_21;
  assign mData_22 = WeightCache_mData_22;
  assign mData_23 = WeightCache_mData_23;
  assign mData_24 = WeightCache_mData_24;
  assign mData_25 = WeightCache_mData_25;
  assign mData_26 = WeightCache_mData_26;
  assign mData_27 = WeightCache_mData_27;
  assign mData_28 = WeightCache_mData_28;
  assign mData_29 = WeightCache_mData_29;
  assign mData_30 = WeightCache_mData_30;
  assign mData_31 = WeightCache_mData_31;
  assign mData_32 = WeightCache_mData_32;
  assign mData_33 = WeightCache_mData_33;
  assign mData_34 = WeightCache_mData_34;
  assign mData_35 = WeightCache_mData_35;
  assign mData_36 = WeightCache_mData_36;
  assign mData_37 = WeightCache_mData_37;
  assign mData_38 = WeightCache_mData_38;
  assign mData_39 = WeightCache_mData_39;
  assign mData_40 = WeightCache_mData_40;
  assign mData_41 = WeightCache_mData_41;
  assign mData_42 = WeightCache_mData_42;
  assign mData_43 = WeightCache_mData_43;
  assign mData_44 = WeightCache_mData_44;
  assign mData_45 = WeightCache_mData_45;
  assign mData_46 = WeightCache_mData_46;
  assign mData_47 = WeightCache_mData_47;
  assign mData_48 = WeightCache_mData_48;
  assign mData_49 = WeightCache_mData_49;
  assign mData_50 = WeightCache_mData_50;
  assign mData_51 = WeightCache_mData_51;
  assign mData_52 = WeightCache_mData_52;
  assign mData_53 = WeightCache_mData_53;
  assign mData_54 = WeightCache_mData_54;
  assign mData_55 = WeightCache_mData_55;
  assign mData_56 = WeightCache_mData_56;
  assign mData_57 = WeightCache_mData_57;
  assign mData_58 = WeightCache_mData_58;
  assign mData_59 = WeightCache_mData_59;
  assign mData_60 = WeightCache_mData_60;
  assign mData_61 = WeightCache_mData_61;
  assign mData_62 = WeightCache_mData_62;
  assign mData_63 = WeightCache_mData_63;
  assign Weight_Cached = WeightCache_Weight_Cached;
  assign MatrixCol_Switch = WeightCache_MatrixCol_Switch;
  assign s_axis_s2mm_tready = WeightCache_sData_ready;

endmodule

module SA_3D (
  input               start,
  input      [7:0]    _zz_io_MatrixA_0,
  input      [7:0]    _zz_io_MatrixA_1,
  input      [7:0]    _zz_io_MatrixA_2,
  input      [7:0]    _zz_io_MatrixA_3,
  input      [7:0]    _zz_io_MatrixA_4,
  input      [7:0]    _zz_io_MatrixA_5,
  input      [7:0]    _zz_io_MatrixA_6,
  input      [7:0]    _zz_io_MatrixA_7,
  input      [7:0]    _zz_io_MatrixB_0,
  input      [7:0]    _zz_io_MatrixB_1,
  input      [7:0]    _zz_io_MatrixB_2,
  input      [7:0]    _zz_io_MatrixB_3,
  input      [7:0]    _zz_io_MatrixB_4,
  input      [7:0]    _zz_io_MatrixB_5,
  input      [7:0]    _zz_io_MatrixB_6,
  input      [7:0]    _zz_io_MatrixB_7,
  input      [7:0]    _zz_io_MatrixB_8,
  input      [7:0]    _zz_io_MatrixB_9,
  input      [7:0]    _zz_io_MatrixB_10,
  input      [7:0]    _zz_io_MatrixB_11,
  input      [7:0]    _zz_io_MatrixB_12,
  input      [7:0]    _zz_io_MatrixB_13,
  input      [7:0]    _zz_io_MatrixB_14,
  input      [7:0]    _zz_io_MatrixB_15,
  input      [7:0]    _zz_io_MatrixB_16,
  input      [7:0]    _zz_io_MatrixB_17,
  input      [7:0]    _zz_io_MatrixB_18,
  input      [7:0]    _zz_io_MatrixB_19,
  input      [7:0]    _zz_io_MatrixB_20,
  input      [7:0]    _zz_io_MatrixB_21,
  input      [7:0]    _zz_io_MatrixB_22,
  input      [7:0]    _zz_io_MatrixB_23,
  input      [7:0]    _zz_io_MatrixB_24,
  input      [7:0]    _zz_io_MatrixB_25,
  input      [7:0]    _zz_io_MatrixB_26,
  input      [7:0]    _zz_io_MatrixB_27,
  input      [7:0]    _zz_io_MatrixB_28,
  input      [7:0]    _zz_io_MatrixB_29,
  input      [7:0]    _zz_io_MatrixB_30,
  input      [7:0]    _zz_io_MatrixB_31,
  input      [7:0]    _zz_io_MatrixB_32,
  input      [7:0]    _zz_io_MatrixB_33,
  input      [7:0]    _zz_io_MatrixB_34,
  input      [7:0]    _zz_io_MatrixB_35,
  input      [7:0]    _zz_io_MatrixB_36,
  input      [7:0]    _zz_io_MatrixB_37,
  input      [7:0]    _zz_io_MatrixB_38,
  input      [7:0]    _zz_io_MatrixB_39,
  input      [7:0]    _zz_io_MatrixB_40,
  input      [7:0]    _zz_io_MatrixB_41,
  input      [7:0]    _zz_io_MatrixB_42,
  input      [7:0]    _zz_io_MatrixB_43,
  input      [7:0]    _zz_io_MatrixB_44,
  input      [7:0]    _zz_io_MatrixB_45,
  input      [7:0]    _zz_io_MatrixB_46,
  input      [7:0]    _zz_io_MatrixB_47,
  input      [7:0]    _zz_io_MatrixB_48,
  input      [7:0]    _zz_io_MatrixB_49,
  input      [7:0]    _zz_io_MatrixB_50,
  input      [7:0]    _zz_io_MatrixB_51,
  input      [7:0]    _zz_io_MatrixB_52,
  input      [7:0]    _zz_io_MatrixB_53,
  input      [7:0]    _zz_io_MatrixB_54,
  input      [7:0]    _zz_io_MatrixB_55,
  input      [7:0]    _zz_io_MatrixB_56,
  input      [7:0]    _zz_io_MatrixB_57,
  input      [7:0]    _zz_io_MatrixB_58,
  input      [7:0]    _zz_io_MatrixB_59,
  input      [7:0]    _zz_io_MatrixB_60,
  input      [7:0]    _zz_io_MatrixB_61,
  input      [7:0]    _zz_io_MatrixB_62,
  input      [7:0]    _zz_io_MatrixB_63,
  input               _zz_io_A_Valid_0,
  input               _zz_io_A_Valid_1,
  input               _zz_io_A_Valid_2,
  input               _zz_io_A_Valid_3,
  input               _zz_io_A_Valid_4,
  input               _zz_io_A_Valid_5,
  input               _zz_io_A_Valid_6,
  input               _zz_io_A_Valid_7,
  input               _zz_io_B_Valid_0,
  input               _zz_io_B_Valid_1,
  input               _zz_io_B_Valid_2,
  input               _zz_io_B_Valid_3,
  input               _zz_io_B_Valid_4,
  input               _zz_io_B_Valid_5,
  input               _zz_io_B_Valid_6,
  input               _zz_io_B_Valid_7,
  input               _zz_io_B_Valid_8,
  input               _zz_io_B_Valid_9,
  input               _zz_io_B_Valid_10,
  input               _zz_io_B_Valid_11,
  input               _zz_io_B_Valid_12,
  input               _zz_io_B_Valid_13,
  input               _zz_io_B_Valid_14,
  input               _zz_io_B_Valid_15,
  input               _zz_io_B_Valid_16,
  input               _zz_io_B_Valid_17,
  input               _zz_io_B_Valid_18,
  input               _zz_io_B_Valid_19,
  input               _zz_io_B_Valid_20,
  input               _zz_io_B_Valid_21,
  input               _zz_io_B_Valid_22,
  input               _zz_io_B_Valid_23,
  input               _zz_io_B_Valid_24,
  input               _zz_io_B_Valid_25,
  input               _zz_io_B_Valid_26,
  input               _zz_io_B_Valid_27,
  input               _zz_io_B_Valid_28,
  input               _zz_io_B_Valid_29,
  input               _zz_io_B_Valid_30,
  input               _zz_io_B_Valid_31,
  input               _zz_io_B_Valid_32,
  input               _zz_io_B_Valid_33,
  input               _zz_io_B_Valid_34,
  input               _zz_io_B_Valid_35,
  input               _zz_io_B_Valid_36,
  input               _zz_io_B_Valid_37,
  input               _zz_io_B_Valid_38,
  input               _zz_io_B_Valid_39,
  input               _zz_io_B_Valid_40,
  input               _zz_io_B_Valid_41,
  input               _zz_io_B_Valid_42,
  input               _zz_io_B_Valid_43,
  input               _zz_io_B_Valid_44,
  input               _zz_io_B_Valid_45,
  input               _zz_io_B_Valid_46,
  input               _zz_io_B_Valid_47,
  input               _zz_io_B_Valid_48,
  input               _zz_io_B_Valid_49,
  input               _zz_io_B_Valid_50,
  input               _zz_io_B_Valid_51,
  input               _zz_io_B_Valid_52,
  input               _zz_io_B_Valid_53,
  input               _zz_io_B_Valid_54,
  input               _zz_io_B_Valid_55,
  input               _zz_io_B_Valid_56,
  input               _zz_io_B_Valid_57,
  input               _zz_io_B_Valid_58,
  input               _zz_io_B_Valid_59,
  input               _zz_io_B_Valid_60,
  input               _zz_io_B_Valid_61,
  input               _zz_io_B_Valid_62,
  input               _zz_io_B_Valid_63,
  input      [15:0]   _zz_io_signCount,
  input               clk,
  output              Matrix_C_valid_0,
  output              Matrix_C_valid_1,
  output              Matrix_C_valid_2,
  output              Matrix_C_valid_3,
  output              Matrix_C_valid_4,
  output              Matrix_C_valid_5,
  output              Matrix_C_valid_6,
  output              Matrix_C_valid_7,
  output     [31:0]   Matrix_C_payload_0,
  output     [31:0]   Matrix_C_payload_1,
  output     [31:0]   Matrix_C_payload_2,
  output     [31:0]   Matrix_C_payload_3,
  output     [31:0]   Matrix_C_payload_4,
  output     [31:0]   Matrix_C_payload_5,
  output     [31:0]   Matrix_C_payload_6,
  output     [31:0]   Matrix_C_payload_7,
  input               reset
);

  wire       [31:0]   Slice0_MatrixC_0;
  wire       [31:0]   Slice0_MatrixC_1;
  wire       [31:0]   Slice0_MatrixC_2;
  wire       [31:0]   Slice0_MatrixC_3;
  wire       [31:0]   Slice0_MatrixC_4;
  wire       [31:0]   Slice0_MatrixC_5;
  wire       [31:0]   Slice0_MatrixC_6;
  wire       [31:0]   Slice0_MatrixC_7;
  wire                Slice0_C_Valid_0;
  wire                Slice0_C_Valid_1;
  wire                Slice0_C_Valid_2;
  wire                Slice0_C_Valid_3;
  wire                Slice0_C_Valid_4;
  wire                Slice0_C_Valid_5;
  wire                Slice0_C_Valid_6;
  wire                Slice0_C_Valid_7;
  reg                 SubModule_SA_3D_Slice0_C_Valid_0_delay_1;
  reg                 SubModule_SA_3D_Slice0_C_Valid_0_delay_2;
  reg                 SubModule_SA_3D_Slice0_C_Valid_0_delay_3;
  reg                 SubModule_SA_3D_Slice0_C_Valid_0_delay_4;
  reg                 SubModule_SA_3D_Slice0_C_Valid_0_delay_5;
  reg                 SubModule_SA_3D_Slice0_C_Valid_0_delay_6;
  reg                 SubModule_SA_3D_Slice0_C_Valid_0_delay_7;
  reg                 SubModule_SA_3D_Slice0_C_Valid_0_delay_8;
  reg                 SubModule_SA_3D_Slice0_C_Valid_0_delay_9;
  reg        [31:0]   _zz_Matrix_C_payload_0;
  reg        [31:0]   _zz_Matrix_C_payload_0_1;
  reg        [31:0]   _zz_Matrix_C_payload_0_2;
  reg        [31:0]   _zz_Matrix_C_payload_0_3;
  reg        [31:0]   _zz_Matrix_C_payload_0_4;
  reg        [31:0]   _zz_Matrix_C_payload_0_5;
  reg        [31:0]   _zz_Matrix_C_payload_0_6;
  reg        [31:0]   _zz_Matrix_C_payload_0_7;
  reg        [31:0]   _zz_Matrix_C_payload_0_8;
  reg                 SubModule_SA_3D_Slice0_C_Valid_1_delay_1;
  reg                 SubModule_SA_3D_Slice0_C_Valid_1_delay_2;
  reg                 SubModule_SA_3D_Slice0_C_Valid_1_delay_3;
  reg                 SubModule_SA_3D_Slice0_C_Valid_1_delay_4;
  reg                 SubModule_SA_3D_Slice0_C_Valid_1_delay_5;
  reg                 SubModule_SA_3D_Slice0_C_Valid_1_delay_6;
  reg                 SubModule_SA_3D_Slice0_C_Valid_1_delay_7;
  reg                 SubModule_SA_3D_Slice0_C_Valid_1_delay_8;
  reg        [31:0]   _zz_Matrix_C_payload_1;
  reg        [31:0]   _zz_Matrix_C_payload_1_1;
  reg        [31:0]   _zz_Matrix_C_payload_1_2;
  reg        [31:0]   _zz_Matrix_C_payload_1_3;
  reg        [31:0]   _zz_Matrix_C_payload_1_4;
  reg        [31:0]   _zz_Matrix_C_payload_1_5;
  reg        [31:0]   _zz_Matrix_C_payload_1_6;
  reg        [31:0]   _zz_Matrix_C_payload_1_7;
  reg                 SubModule_SA_3D_Slice0_C_Valid_2_delay_1;
  reg                 SubModule_SA_3D_Slice0_C_Valid_2_delay_2;
  reg                 SubModule_SA_3D_Slice0_C_Valid_2_delay_3;
  reg                 SubModule_SA_3D_Slice0_C_Valid_2_delay_4;
  reg                 SubModule_SA_3D_Slice0_C_Valid_2_delay_5;
  reg                 SubModule_SA_3D_Slice0_C_Valid_2_delay_6;
  reg                 SubModule_SA_3D_Slice0_C_Valid_2_delay_7;
  reg        [31:0]   _zz_Matrix_C_payload_2;
  reg        [31:0]   _zz_Matrix_C_payload_2_1;
  reg        [31:0]   _zz_Matrix_C_payload_2_2;
  reg        [31:0]   _zz_Matrix_C_payload_2_3;
  reg        [31:0]   _zz_Matrix_C_payload_2_4;
  reg        [31:0]   _zz_Matrix_C_payload_2_5;
  reg        [31:0]   _zz_Matrix_C_payload_2_6;
  reg                 SubModule_SA_3D_Slice0_C_Valid_3_delay_1;
  reg                 SubModule_SA_3D_Slice0_C_Valid_3_delay_2;
  reg                 SubModule_SA_3D_Slice0_C_Valid_3_delay_3;
  reg                 SubModule_SA_3D_Slice0_C_Valid_3_delay_4;
  reg                 SubModule_SA_3D_Slice0_C_Valid_3_delay_5;
  reg                 SubModule_SA_3D_Slice0_C_Valid_3_delay_6;
  reg        [31:0]   _zz_Matrix_C_payload_3;
  reg        [31:0]   _zz_Matrix_C_payload_3_1;
  reg        [31:0]   _zz_Matrix_C_payload_3_2;
  reg        [31:0]   _zz_Matrix_C_payload_3_3;
  reg        [31:0]   _zz_Matrix_C_payload_3_4;
  reg        [31:0]   _zz_Matrix_C_payload_3_5;
  reg                 SubModule_SA_3D_Slice0_C_Valid_4_delay_1;
  reg                 SubModule_SA_3D_Slice0_C_Valid_4_delay_2;
  reg                 SubModule_SA_3D_Slice0_C_Valid_4_delay_3;
  reg                 SubModule_SA_3D_Slice0_C_Valid_4_delay_4;
  reg                 SubModule_SA_3D_Slice0_C_Valid_4_delay_5;
  reg        [31:0]   _zz_Matrix_C_payload_4;
  reg        [31:0]   _zz_Matrix_C_payload_4_1;
  reg        [31:0]   _zz_Matrix_C_payload_4_2;
  reg        [31:0]   _zz_Matrix_C_payload_4_3;
  reg        [31:0]   _zz_Matrix_C_payload_4_4;
  reg                 SubModule_SA_3D_Slice0_C_Valid_5_delay_1;
  reg                 SubModule_SA_3D_Slice0_C_Valid_5_delay_2;
  reg                 SubModule_SA_3D_Slice0_C_Valid_5_delay_3;
  reg                 SubModule_SA_3D_Slice0_C_Valid_5_delay_4;
  reg        [31:0]   _zz_Matrix_C_payload_5;
  reg        [31:0]   _zz_Matrix_C_payload_5_1;
  reg        [31:0]   _zz_Matrix_C_payload_5_2;
  reg        [31:0]   _zz_Matrix_C_payload_5_3;
  reg                 SubModule_SA_3D_Slice0_C_Valid_6_delay_1;
  reg                 SubModule_SA_3D_Slice0_C_Valid_6_delay_2;
  reg                 SubModule_SA_3D_Slice0_C_Valid_6_delay_3;
  reg        [31:0]   _zz_Matrix_C_payload_6;
  reg        [31:0]   _zz_Matrix_C_payload_6_1;
  reg        [31:0]   _zz_Matrix_C_payload_6_2;
  reg                 SubModule_SA_3D_Slice0_C_Valid_7_delay_1;
  reg                 SubModule_SA_3D_Slice0_C_Valid_7_delay_2;
  reg        [31:0]   _zz_Matrix_C_payload_7;
  reg        [31:0]   _zz_Matrix_C_payload_7_1;

  SA_2D Slice0 (
    .io_MatrixA_0  (_zz_io_MatrixA_0[7:0] ), //i
    .io_MatrixA_1  (_zz_io_MatrixA_1[7:0] ), //i
    .io_MatrixA_2  (_zz_io_MatrixA_2[7:0] ), //i
    .io_MatrixA_3  (_zz_io_MatrixA_3[7:0] ), //i
    .io_MatrixA_4  (_zz_io_MatrixA_4[7:0] ), //i
    .io_MatrixA_5  (_zz_io_MatrixA_5[7:0] ), //i
    .io_MatrixA_6  (_zz_io_MatrixA_6[7:0] ), //i
    .io_MatrixA_7  (_zz_io_MatrixA_7[7:0] ), //i
    .io_MatrixB_0  (_zz_io_MatrixB_0[7:0] ), //i
    .io_MatrixB_1  (_zz_io_MatrixB_1[7:0] ), //i
    .io_MatrixB_2  (_zz_io_MatrixB_2[7:0] ), //i
    .io_MatrixB_3  (_zz_io_MatrixB_3[7:0] ), //i
    .io_MatrixB_4  (_zz_io_MatrixB_4[7:0] ), //i
    .io_MatrixB_5  (_zz_io_MatrixB_5[7:0] ), //i
    .io_MatrixB_6  (_zz_io_MatrixB_6[7:0] ), //i
    .io_MatrixB_7  (_zz_io_MatrixB_7[7:0] ), //i
    .io_MatrixB_8  (_zz_io_MatrixB_8[7:0] ), //i
    .io_MatrixB_9  (_zz_io_MatrixB_9[7:0] ), //i
    .io_MatrixB_10 (_zz_io_MatrixB_10[7:0]), //i
    .io_MatrixB_11 (_zz_io_MatrixB_11[7:0]), //i
    .io_MatrixB_12 (_zz_io_MatrixB_12[7:0]), //i
    .io_MatrixB_13 (_zz_io_MatrixB_13[7:0]), //i
    .io_MatrixB_14 (_zz_io_MatrixB_14[7:0]), //i
    .io_MatrixB_15 (_zz_io_MatrixB_15[7:0]), //i
    .io_MatrixB_16 (_zz_io_MatrixB_16[7:0]), //i
    .io_MatrixB_17 (_zz_io_MatrixB_17[7:0]), //i
    .io_MatrixB_18 (_zz_io_MatrixB_18[7:0]), //i
    .io_MatrixB_19 (_zz_io_MatrixB_19[7:0]), //i
    .io_MatrixB_20 (_zz_io_MatrixB_20[7:0]), //i
    .io_MatrixB_21 (_zz_io_MatrixB_21[7:0]), //i
    .io_MatrixB_22 (_zz_io_MatrixB_22[7:0]), //i
    .io_MatrixB_23 (_zz_io_MatrixB_23[7:0]), //i
    .io_MatrixB_24 (_zz_io_MatrixB_24[7:0]), //i
    .io_MatrixB_25 (_zz_io_MatrixB_25[7:0]), //i
    .io_MatrixB_26 (_zz_io_MatrixB_26[7:0]), //i
    .io_MatrixB_27 (_zz_io_MatrixB_27[7:0]), //i
    .io_MatrixB_28 (_zz_io_MatrixB_28[7:0]), //i
    .io_MatrixB_29 (_zz_io_MatrixB_29[7:0]), //i
    .io_MatrixB_30 (_zz_io_MatrixB_30[7:0]), //i
    .io_MatrixB_31 (_zz_io_MatrixB_31[7:0]), //i
    .io_MatrixB_32 (_zz_io_MatrixB_32[7:0]), //i
    .io_MatrixB_33 (_zz_io_MatrixB_33[7:0]), //i
    .io_MatrixB_34 (_zz_io_MatrixB_34[7:0]), //i
    .io_MatrixB_35 (_zz_io_MatrixB_35[7:0]), //i
    .io_MatrixB_36 (_zz_io_MatrixB_36[7:0]), //i
    .io_MatrixB_37 (_zz_io_MatrixB_37[7:0]), //i
    .io_MatrixB_38 (_zz_io_MatrixB_38[7:0]), //i
    .io_MatrixB_39 (_zz_io_MatrixB_39[7:0]), //i
    .io_MatrixB_40 (_zz_io_MatrixB_40[7:0]), //i
    .io_MatrixB_41 (_zz_io_MatrixB_41[7:0]), //i
    .io_MatrixB_42 (_zz_io_MatrixB_42[7:0]), //i
    .io_MatrixB_43 (_zz_io_MatrixB_43[7:0]), //i
    .io_MatrixB_44 (_zz_io_MatrixB_44[7:0]), //i
    .io_MatrixB_45 (_zz_io_MatrixB_45[7:0]), //i
    .io_MatrixB_46 (_zz_io_MatrixB_46[7:0]), //i
    .io_MatrixB_47 (_zz_io_MatrixB_47[7:0]), //i
    .io_MatrixB_48 (_zz_io_MatrixB_48[7:0]), //i
    .io_MatrixB_49 (_zz_io_MatrixB_49[7:0]), //i
    .io_MatrixB_50 (_zz_io_MatrixB_50[7:0]), //i
    .io_MatrixB_51 (_zz_io_MatrixB_51[7:0]), //i
    .io_MatrixB_52 (_zz_io_MatrixB_52[7:0]), //i
    .io_MatrixB_53 (_zz_io_MatrixB_53[7:0]), //i
    .io_MatrixB_54 (_zz_io_MatrixB_54[7:0]), //i
    .io_MatrixB_55 (_zz_io_MatrixB_55[7:0]), //i
    .io_MatrixB_56 (_zz_io_MatrixB_56[7:0]), //i
    .io_MatrixB_57 (_zz_io_MatrixB_57[7:0]), //i
    .io_MatrixB_58 (_zz_io_MatrixB_58[7:0]), //i
    .io_MatrixB_59 (_zz_io_MatrixB_59[7:0]), //i
    .io_MatrixB_60 (_zz_io_MatrixB_60[7:0]), //i
    .io_MatrixB_61 (_zz_io_MatrixB_61[7:0]), //i
    .io_MatrixB_62 (_zz_io_MatrixB_62[7:0]), //i
    .io_MatrixB_63 (_zz_io_MatrixB_63[7:0]), //i
    .io_A_Valid_0  (_zz_io_A_Valid_0      ), //i
    .io_A_Valid_1  (_zz_io_A_Valid_1      ), //i
    .io_A_Valid_2  (_zz_io_A_Valid_2      ), //i
    .io_A_Valid_3  (_zz_io_A_Valid_3      ), //i
    .io_A_Valid_4  (_zz_io_A_Valid_4      ), //i
    .io_A_Valid_5  (_zz_io_A_Valid_5      ), //i
    .io_A_Valid_6  (_zz_io_A_Valid_6      ), //i
    .io_A_Valid_7  (_zz_io_A_Valid_7      ), //i
    .io_B_Valid_0  (_zz_io_B_Valid_0      ), //i
    .io_B_Valid_1  (_zz_io_B_Valid_1      ), //i
    .io_B_Valid_2  (_zz_io_B_Valid_2      ), //i
    .io_B_Valid_3  (_zz_io_B_Valid_3      ), //i
    .io_B_Valid_4  (_zz_io_B_Valid_4      ), //i
    .io_B_Valid_5  (_zz_io_B_Valid_5      ), //i
    .io_B_Valid_6  (_zz_io_B_Valid_6      ), //i
    .io_B_Valid_7  (_zz_io_B_Valid_7      ), //i
    .io_B_Valid_8  (_zz_io_B_Valid_8      ), //i
    .io_B_Valid_9  (_zz_io_B_Valid_9      ), //i
    .io_B_Valid_10 (_zz_io_B_Valid_10     ), //i
    .io_B_Valid_11 (_zz_io_B_Valid_11     ), //i
    .io_B_Valid_12 (_zz_io_B_Valid_12     ), //i
    .io_B_Valid_13 (_zz_io_B_Valid_13     ), //i
    .io_B_Valid_14 (_zz_io_B_Valid_14     ), //i
    .io_B_Valid_15 (_zz_io_B_Valid_15     ), //i
    .io_B_Valid_16 (_zz_io_B_Valid_16     ), //i
    .io_B_Valid_17 (_zz_io_B_Valid_17     ), //i
    .io_B_Valid_18 (_zz_io_B_Valid_18     ), //i
    .io_B_Valid_19 (_zz_io_B_Valid_19     ), //i
    .io_B_Valid_20 (_zz_io_B_Valid_20     ), //i
    .io_B_Valid_21 (_zz_io_B_Valid_21     ), //i
    .io_B_Valid_22 (_zz_io_B_Valid_22     ), //i
    .io_B_Valid_23 (_zz_io_B_Valid_23     ), //i
    .io_B_Valid_24 (_zz_io_B_Valid_24     ), //i
    .io_B_Valid_25 (_zz_io_B_Valid_25     ), //i
    .io_B_Valid_26 (_zz_io_B_Valid_26     ), //i
    .io_B_Valid_27 (_zz_io_B_Valid_27     ), //i
    .io_B_Valid_28 (_zz_io_B_Valid_28     ), //i
    .io_B_Valid_29 (_zz_io_B_Valid_29     ), //i
    .io_B_Valid_30 (_zz_io_B_Valid_30     ), //i
    .io_B_Valid_31 (_zz_io_B_Valid_31     ), //i
    .io_B_Valid_32 (_zz_io_B_Valid_32     ), //i
    .io_B_Valid_33 (_zz_io_B_Valid_33     ), //i
    .io_B_Valid_34 (_zz_io_B_Valid_34     ), //i
    .io_B_Valid_35 (_zz_io_B_Valid_35     ), //i
    .io_B_Valid_36 (_zz_io_B_Valid_36     ), //i
    .io_B_Valid_37 (_zz_io_B_Valid_37     ), //i
    .io_B_Valid_38 (_zz_io_B_Valid_38     ), //i
    .io_B_Valid_39 (_zz_io_B_Valid_39     ), //i
    .io_B_Valid_40 (_zz_io_B_Valid_40     ), //i
    .io_B_Valid_41 (_zz_io_B_Valid_41     ), //i
    .io_B_Valid_42 (_zz_io_B_Valid_42     ), //i
    .io_B_Valid_43 (_zz_io_B_Valid_43     ), //i
    .io_B_Valid_44 (_zz_io_B_Valid_44     ), //i
    .io_B_Valid_45 (_zz_io_B_Valid_45     ), //i
    .io_B_Valid_46 (_zz_io_B_Valid_46     ), //i
    .io_B_Valid_47 (_zz_io_B_Valid_47     ), //i
    .io_B_Valid_48 (_zz_io_B_Valid_48     ), //i
    .io_B_Valid_49 (_zz_io_B_Valid_49     ), //i
    .io_B_Valid_50 (_zz_io_B_Valid_50     ), //i
    .io_B_Valid_51 (_zz_io_B_Valid_51     ), //i
    .io_B_Valid_52 (_zz_io_B_Valid_52     ), //i
    .io_B_Valid_53 (_zz_io_B_Valid_53     ), //i
    .io_B_Valid_54 (_zz_io_B_Valid_54     ), //i
    .io_B_Valid_55 (_zz_io_B_Valid_55     ), //i
    .io_B_Valid_56 (_zz_io_B_Valid_56     ), //i
    .io_B_Valid_57 (_zz_io_B_Valid_57     ), //i
    .io_B_Valid_58 (_zz_io_B_Valid_58     ), //i
    .io_B_Valid_59 (_zz_io_B_Valid_59     ), //i
    .io_B_Valid_60 (_zz_io_B_Valid_60     ), //i
    .io_B_Valid_61 (_zz_io_B_Valid_61     ), //i
    .io_B_Valid_62 (_zz_io_B_Valid_62     ), //i
    .io_B_Valid_63 (_zz_io_B_Valid_63     ), //i
    .io_signCount  (_zz_io_signCount[15:0]), //i
    .MatrixC_0     (Slice0_MatrixC_0[31:0]), //o
    .MatrixC_1     (Slice0_MatrixC_1[31:0]), //o
    .MatrixC_2     (Slice0_MatrixC_2[31:0]), //o
    .MatrixC_3     (Slice0_MatrixC_3[31:0]), //o
    .MatrixC_4     (Slice0_MatrixC_4[31:0]), //o
    .MatrixC_5     (Slice0_MatrixC_5[31:0]), //o
    .MatrixC_6     (Slice0_MatrixC_6[31:0]), //o
    .MatrixC_7     (Slice0_MatrixC_7[31:0]), //o
    .C_Valid_0     (Slice0_C_Valid_0      ), //o
    .C_Valid_1     (Slice0_C_Valid_1      ), //o
    .C_Valid_2     (Slice0_C_Valid_2      ), //o
    .C_Valid_3     (Slice0_C_Valid_3      ), //o
    .C_Valid_4     (Slice0_C_Valid_4      ), //o
    .C_Valid_5     (Slice0_C_Valid_5      ), //o
    .C_Valid_6     (Slice0_C_Valid_6      ), //o
    .C_Valid_7     (Slice0_C_Valid_7      ), //o
    .start         (start                 ), //i
    .clk           (clk                   ), //i
    .reset         (reset                 )  //i
  );
  assign Matrix_C_valid_0 = SubModule_SA_3D_Slice0_C_Valid_0_delay_9;
  assign Matrix_C_payload_0[31 : 0] = _zz_Matrix_C_payload_0_8;
  assign Matrix_C_valid_1 = SubModule_SA_3D_Slice0_C_Valid_1_delay_8;
  assign Matrix_C_payload_1[31 : 0] = _zz_Matrix_C_payload_1_7;
  assign Matrix_C_valid_2 = SubModule_SA_3D_Slice0_C_Valid_2_delay_7;
  assign Matrix_C_payload_2[31 : 0] = _zz_Matrix_C_payload_2_6;
  assign Matrix_C_valid_3 = SubModule_SA_3D_Slice0_C_Valid_3_delay_6;
  assign Matrix_C_payload_3[31 : 0] = _zz_Matrix_C_payload_3_5;
  assign Matrix_C_valid_4 = SubModule_SA_3D_Slice0_C_Valid_4_delay_5;
  assign Matrix_C_payload_4[31 : 0] = _zz_Matrix_C_payload_4_4;
  assign Matrix_C_valid_5 = SubModule_SA_3D_Slice0_C_Valid_5_delay_4;
  assign Matrix_C_payload_5[31 : 0] = _zz_Matrix_C_payload_5_3;
  assign Matrix_C_valid_6 = SubModule_SA_3D_Slice0_C_Valid_6_delay_3;
  assign Matrix_C_payload_6[31 : 0] = _zz_Matrix_C_payload_6_2;
  assign Matrix_C_valid_7 = SubModule_SA_3D_Slice0_C_Valid_7_delay_2;
  assign Matrix_C_payload_7[31 : 0] = _zz_Matrix_C_payload_7_1;
  always @(posedge clk) begin
    SubModule_SA_3D_Slice0_C_Valid_0_delay_1 <= Slice0_C_Valid_0;
    SubModule_SA_3D_Slice0_C_Valid_0_delay_2 <= SubModule_SA_3D_Slice0_C_Valid_0_delay_1;
    SubModule_SA_3D_Slice0_C_Valid_0_delay_3 <= SubModule_SA_3D_Slice0_C_Valid_0_delay_2;
    SubModule_SA_3D_Slice0_C_Valid_0_delay_4 <= SubModule_SA_3D_Slice0_C_Valid_0_delay_3;
    SubModule_SA_3D_Slice0_C_Valid_0_delay_5 <= SubModule_SA_3D_Slice0_C_Valid_0_delay_4;
    SubModule_SA_3D_Slice0_C_Valid_0_delay_6 <= SubModule_SA_3D_Slice0_C_Valid_0_delay_5;
    SubModule_SA_3D_Slice0_C_Valid_0_delay_7 <= SubModule_SA_3D_Slice0_C_Valid_0_delay_6;
    SubModule_SA_3D_Slice0_C_Valid_0_delay_8 <= SubModule_SA_3D_Slice0_C_Valid_0_delay_7;
    SubModule_SA_3D_Slice0_C_Valid_0_delay_9 <= SubModule_SA_3D_Slice0_C_Valid_0_delay_8;
    _zz_Matrix_C_payload_0 <= Slice0_MatrixC_0;
    _zz_Matrix_C_payload_0_1 <= _zz_Matrix_C_payload_0;
    _zz_Matrix_C_payload_0_2 <= _zz_Matrix_C_payload_0_1;
    _zz_Matrix_C_payload_0_3 <= _zz_Matrix_C_payload_0_2;
    _zz_Matrix_C_payload_0_4 <= _zz_Matrix_C_payload_0_3;
    _zz_Matrix_C_payload_0_5 <= _zz_Matrix_C_payload_0_4;
    _zz_Matrix_C_payload_0_6 <= _zz_Matrix_C_payload_0_5;
    _zz_Matrix_C_payload_0_7 <= _zz_Matrix_C_payload_0_6;
    _zz_Matrix_C_payload_0_8 <= _zz_Matrix_C_payload_0_7;
    SubModule_SA_3D_Slice0_C_Valid_1_delay_1 <= Slice0_C_Valid_1;
    SubModule_SA_3D_Slice0_C_Valid_1_delay_2 <= SubModule_SA_3D_Slice0_C_Valid_1_delay_1;
    SubModule_SA_3D_Slice0_C_Valid_1_delay_3 <= SubModule_SA_3D_Slice0_C_Valid_1_delay_2;
    SubModule_SA_3D_Slice0_C_Valid_1_delay_4 <= SubModule_SA_3D_Slice0_C_Valid_1_delay_3;
    SubModule_SA_3D_Slice0_C_Valid_1_delay_5 <= SubModule_SA_3D_Slice0_C_Valid_1_delay_4;
    SubModule_SA_3D_Slice0_C_Valid_1_delay_6 <= SubModule_SA_3D_Slice0_C_Valid_1_delay_5;
    SubModule_SA_3D_Slice0_C_Valid_1_delay_7 <= SubModule_SA_3D_Slice0_C_Valid_1_delay_6;
    SubModule_SA_3D_Slice0_C_Valid_1_delay_8 <= SubModule_SA_3D_Slice0_C_Valid_1_delay_7;
    _zz_Matrix_C_payload_1 <= Slice0_MatrixC_1;
    _zz_Matrix_C_payload_1_1 <= _zz_Matrix_C_payload_1;
    _zz_Matrix_C_payload_1_2 <= _zz_Matrix_C_payload_1_1;
    _zz_Matrix_C_payload_1_3 <= _zz_Matrix_C_payload_1_2;
    _zz_Matrix_C_payload_1_4 <= _zz_Matrix_C_payload_1_3;
    _zz_Matrix_C_payload_1_5 <= _zz_Matrix_C_payload_1_4;
    _zz_Matrix_C_payload_1_6 <= _zz_Matrix_C_payload_1_5;
    _zz_Matrix_C_payload_1_7 <= _zz_Matrix_C_payload_1_6;
    SubModule_SA_3D_Slice0_C_Valid_2_delay_1 <= Slice0_C_Valid_2;
    SubModule_SA_3D_Slice0_C_Valid_2_delay_2 <= SubModule_SA_3D_Slice0_C_Valid_2_delay_1;
    SubModule_SA_3D_Slice0_C_Valid_2_delay_3 <= SubModule_SA_3D_Slice0_C_Valid_2_delay_2;
    SubModule_SA_3D_Slice0_C_Valid_2_delay_4 <= SubModule_SA_3D_Slice0_C_Valid_2_delay_3;
    SubModule_SA_3D_Slice0_C_Valid_2_delay_5 <= SubModule_SA_3D_Slice0_C_Valid_2_delay_4;
    SubModule_SA_3D_Slice0_C_Valid_2_delay_6 <= SubModule_SA_3D_Slice0_C_Valid_2_delay_5;
    SubModule_SA_3D_Slice0_C_Valid_2_delay_7 <= SubModule_SA_3D_Slice0_C_Valid_2_delay_6;
    _zz_Matrix_C_payload_2 <= Slice0_MatrixC_2;
    _zz_Matrix_C_payload_2_1 <= _zz_Matrix_C_payload_2;
    _zz_Matrix_C_payload_2_2 <= _zz_Matrix_C_payload_2_1;
    _zz_Matrix_C_payload_2_3 <= _zz_Matrix_C_payload_2_2;
    _zz_Matrix_C_payload_2_4 <= _zz_Matrix_C_payload_2_3;
    _zz_Matrix_C_payload_2_5 <= _zz_Matrix_C_payload_2_4;
    _zz_Matrix_C_payload_2_6 <= _zz_Matrix_C_payload_2_5;
    SubModule_SA_3D_Slice0_C_Valid_3_delay_1 <= Slice0_C_Valid_3;
    SubModule_SA_3D_Slice0_C_Valid_3_delay_2 <= SubModule_SA_3D_Slice0_C_Valid_3_delay_1;
    SubModule_SA_3D_Slice0_C_Valid_3_delay_3 <= SubModule_SA_3D_Slice0_C_Valid_3_delay_2;
    SubModule_SA_3D_Slice0_C_Valid_3_delay_4 <= SubModule_SA_3D_Slice0_C_Valid_3_delay_3;
    SubModule_SA_3D_Slice0_C_Valid_3_delay_5 <= SubModule_SA_3D_Slice0_C_Valid_3_delay_4;
    SubModule_SA_3D_Slice0_C_Valid_3_delay_6 <= SubModule_SA_3D_Slice0_C_Valid_3_delay_5;
    _zz_Matrix_C_payload_3 <= Slice0_MatrixC_3;
    _zz_Matrix_C_payload_3_1 <= _zz_Matrix_C_payload_3;
    _zz_Matrix_C_payload_3_2 <= _zz_Matrix_C_payload_3_1;
    _zz_Matrix_C_payload_3_3 <= _zz_Matrix_C_payload_3_2;
    _zz_Matrix_C_payload_3_4 <= _zz_Matrix_C_payload_3_3;
    _zz_Matrix_C_payload_3_5 <= _zz_Matrix_C_payload_3_4;
    SubModule_SA_3D_Slice0_C_Valid_4_delay_1 <= Slice0_C_Valid_4;
    SubModule_SA_3D_Slice0_C_Valid_4_delay_2 <= SubModule_SA_3D_Slice0_C_Valid_4_delay_1;
    SubModule_SA_3D_Slice0_C_Valid_4_delay_3 <= SubModule_SA_3D_Slice0_C_Valid_4_delay_2;
    SubModule_SA_3D_Slice0_C_Valid_4_delay_4 <= SubModule_SA_3D_Slice0_C_Valid_4_delay_3;
    SubModule_SA_3D_Slice0_C_Valid_4_delay_5 <= SubModule_SA_3D_Slice0_C_Valid_4_delay_4;
    _zz_Matrix_C_payload_4 <= Slice0_MatrixC_4;
    _zz_Matrix_C_payload_4_1 <= _zz_Matrix_C_payload_4;
    _zz_Matrix_C_payload_4_2 <= _zz_Matrix_C_payload_4_1;
    _zz_Matrix_C_payload_4_3 <= _zz_Matrix_C_payload_4_2;
    _zz_Matrix_C_payload_4_4 <= _zz_Matrix_C_payload_4_3;
    SubModule_SA_3D_Slice0_C_Valid_5_delay_1 <= Slice0_C_Valid_5;
    SubModule_SA_3D_Slice0_C_Valid_5_delay_2 <= SubModule_SA_3D_Slice0_C_Valid_5_delay_1;
    SubModule_SA_3D_Slice0_C_Valid_5_delay_3 <= SubModule_SA_3D_Slice0_C_Valid_5_delay_2;
    SubModule_SA_3D_Slice0_C_Valid_5_delay_4 <= SubModule_SA_3D_Slice0_C_Valid_5_delay_3;
    _zz_Matrix_C_payload_5 <= Slice0_MatrixC_5;
    _zz_Matrix_C_payload_5_1 <= _zz_Matrix_C_payload_5;
    _zz_Matrix_C_payload_5_2 <= _zz_Matrix_C_payload_5_1;
    _zz_Matrix_C_payload_5_3 <= _zz_Matrix_C_payload_5_2;
    SubModule_SA_3D_Slice0_C_Valid_6_delay_1 <= Slice0_C_Valid_6;
    SubModule_SA_3D_Slice0_C_Valid_6_delay_2 <= SubModule_SA_3D_Slice0_C_Valid_6_delay_1;
    SubModule_SA_3D_Slice0_C_Valid_6_delay_3 <= SubModule_SA_3D_Slice0_C_Valid_6_delay_2;
    _zz_Matrix_C_payload_6 <= Slice0_MatrixC_6;
    _zz_Matrix_C_payload_6_1 <= _zz_Matrix_C_payload_6;
    _zz_Matrix_C_payload_6_2 <= _zz_Matrix_C_payload_6_1;
    SubModule_SA_3D_Slice0_C_Valid_7_delay_1 <= Slice0_C_Valid_7;
    SubModule_SA_3D_Slice0_C_Valid_7_delay_2 <= SubModule_SA_3D_Slice0_C_Valid_7_delay_1;
    _zz_Matrix_C_payload_7 <= Slice0_MatrixC_7;
    _zz_Matrix_C_payload_7_1 <= _zz_Matrix_C_payload_7;
  end


endmodule

module Img2ColStreamV2 (
  output reg [63:0]   mData,
  output reg [7:0]    mValid,
  input      [63:0]   s_axis_s2mm_tdata,
  input      [7:0]    s_axis_s2mm_tkeep,
  input               s_axis_s2mm_tlast,
  output              s_axis_s2mm_tready,
  input               s_axis_s2mm_tvalid,
  input               start,
  output              Raddr_Valid,
  output              LayerEnd,
  input      [4:0]    Stride,
  input      [4:0]    Kernel_Size,
  input      [15:0]   Window_Size,
  input      [15:0]   InFeature_Size,
  input      [15:0]   InFeature_Channel,
  input      [15:0]   OutFeature_Channel,
  input      [15:0]   OutFeature_Size,
  input      [15:0]   OutCol_Count_Times,
  input      [15:0]   InCol_Count_Times,
  input      [15:0]   OutRow_Count_Times,
  input      [15:0]   OutFeature_Channel_Count_Times,
  input      [12:0]   Sliding_Size,
  input               clk,
  input               reset
);

  wire                SubModule_Fifo_Clear;
  wire       [15:0]   SubModule_Test_Generate_Period;
  wire                streamFifo_io_push_valid;
  wire                streamFifo_1_io_push_valid;
  wire                streamFifo_2_io_push_valid;
  wire                streamFifo_3_io_push_valid;
  wire                streamFifo_4_io_push_valid;
  wire                streamFifo_5_io_push_valid;
  wire                streamFifo_6_io_push_valid;
  wire                streamFifo_7_io_push_valid;
  wire                SubModule_sData_ready;
  wire       [63:0]   SubModule_mData;
  wire                SubModule_mValid;
  wire                SubModule_mLast;
  wire                SubModule_Test_Signal;
  wire                SubModule_Test_End;
  wire                SubModule_Raddr_Valid;
  wire                SubModule_LayerEnd;
  wire                SubModule_SA_Row_Cnt_Valid;
  wire                streamFifo_io_push_ready;
  wire                streamFifo_io_pop_valid;
  wire       [63:0]   streamFifo_io_pop_payload;
  wire       [4:0]    streamFifo_io_occupancy;
  wire       [4:0]    streamFifo_io_availability;
  wire                axisDataConverter_8_inStream_ready;
  wire                axisDataConverter_8_outStream_valid;
  wire       [7:0]    axisDataConverter_8_outStream_payload;
  wire                streamFifo_1_io_push_ready;
  wire                streamFifo_1_io_pop_valid;
  wire       [63:0]   streamFifo_1_io_pop_payload;
  wire       [4:0]    streamFifo_1_io_occupancy;
  wire       [4:0]    streamFifo_1_io_availability;
  wire                axisDataConverter_9_inStream_ready;
  wire                axisDataConverter_9_outStream_valid;
  wire       [7:0]    axisDataConverter_9_outStream_payload;
  wire                streamFifo_2_io_push_ready;
  wire                streamFifo_2_io_pop_valid;
  wire       [63:0]   streamFifo_2_io_pop_payload;
  wire       [4:0]    streamFifo_2_io_occupancy;
  wire       [4:0]    streamFifo_2_io_availability;
  wire                axisDataConverter_10_inStream_ready;
  wire                axisDataConverter_10_outStream_valid;
  wire       [7:0]    axisDataConverter_10_outStream_payload;
  wire                streamFifo_3_io_push_ready;
  wire                streamFifo_3_io_pop_valid;
  wire       [63:0]   streamFifo_3_io_pop_payload;
  wire       [4:0]    streamFifo_3_io_occupancy;
  wire       [4:0]    streamFifo_3_io_availability;
  wire                axisDataConverter_11_inStream_ready;
  wire                axisDataConverter_11_outStream_valid;
  wire       [7:0]    axisDataConverter_11_outStream_payload;
  wire                streamFifo_4_io_push_ready;
  wire                streamFifo_4_io_pop_valid;
  wire       [63:0]   streamFifo_4_io_pop_payload;
  wire       [4:0]    streamFifo_4_io_occupancy;
  wire       [4:0]    streamFifo_4_io_availability;
  wire                axisDataConverter_12_inStream_ready;
  wire                axisDataConverter_12_outStream_valid;
  wire       [7:0]    axisDataConverter_12_outStream_payload;
  wire                streamFifo_5_io_push_ready;
  wire                streamFifo_5_io_pop_valid;
  wire       [63:0]   streamFifo_5_io_pop_payload;
  wire       [4:0]    streamFifo_5_io_occupancy;
  wire       [4:0]    streamFifo_5_io_availability;
  wire                axisDataConverter_13_inStream_ready;
  wire                axisDataConverter_13_outStream_valid;
  wire       [7:0]    axisDataConverter_13_outStream_payload;
  wire                streamFifo_6_io_push_ready;
  wire                streamFifo_6_io_pop_valid;
  wire       [63:0]   streamFifo_6_io_pop_payload;
  wire       [4:0]    streamFifo_6_io_occupancy;
  wire       [4:0]    streamFifo_6_io_availability;
  wire                axisDataConverter_14_inStream_ready;
  wire                axisDataConverter_14_outStream_valid;
  wire       [7:0]    axisDataConverter_14_outStream_payload;
  wire                streamFifo_7_io_push_ready;
  wire                streamFifo_7_io_pop_valid;
  wire       [63:0]   streamFifo_7_io_pop_payload;
  wire       [4:0]    streamFifo_7_io_occupancy;
  wire       [4:0]    streamFifo_7_io_availability;
  wire                axisDataConverter_15_inStream_ready;
  wire                axisDataConverter_15_outStream_valid;
  wire       [7:0]    axisDataConverter_15_outStream_payload;
  reg        [7:0]    OutData_Switch;
  reg                 Switch_Reset;
  wire                TestValid_Signal_0;
  wire                TestValid_Signal_1;
  wire                TestValid_Signal_2;
  wire                TestValid_Signal_3;
  wire                TestValid_Signal_4;
  wire                TestValid_Signal_5;
  wire                TestValid_Signal_6;
  wire                TestValid_Signal_7;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_8_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_8_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_9_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_9_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_10_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_10_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_11_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_11_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_12_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_12_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_13_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_13_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_14_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_14_outStream_valid_regNext;
  reg        [7:0]    SubModule_Img2Col_axisDataConverter_15_outStream_payload_regNext;
  reg                 SubModule_Img2Col_axisDataConverter_15_outStream_valid_regNext;
  reg                 SubModule_Img2Col_SubModule_LayerEnd_delay_1;
  reg                 SubModule_Img2Col_SubModule_LayerEnd_delay_2;
  reg                 SubModule_Img2Col_SubModule_LayerEnd_delay_3;

  Img2Col_Top SubModule (
    .start                          (start                               ), //i
    .sData_valid                    (s_axis_s2mm_tvalid                  ), //i
    .sData_ready                    (SubModule_sData_ready               ), //o
    .sData_payload                  (s_axis_s2mm_tdata[63:0]             ), //i
    .mData                          (SubModule_mData[63:0]               ), //o
    .mReady                         (streamFifo_io_push_ready            ), //i
    .mValid                         (SubModule_mValid                    ), //o
    .Fifo_Clear                     (SubModule_Fifo_Clear                ), //i
    .mLast                          (SubModule_mLast                     ), //o
    .Stride                         (Stride[4:0]                         ), //i
    .Kernel_Size                    (Kernel_Size[4:0]                    ), //i
    .Window_Size                    (Window_Size[15:0]                   ), //i
    .InFeature_Size                 (InFeature_Size[15:0]                ), //i
    .InFeature_Channel              (InFeature_Channel[15:0]             ), //i
    .OutFeature_Channel             (OutFeature_Channel[15:0]            ), //i
    .OutFeature_Size                (OutFeature_Size[15:0]               ), //i
    .OutCol_Count_Times             (OutCol_Count_Times[15:0]            ), //i
    .InCol_Count_Times              (InCol_Count_Times[15:0]             ), //i
    .OutRow_Count_Times             (OutRow_Count_Times[15:0]            ), //i
    .OutFeature_Channel_Count_Times (OutFeature_Channel_Count_Times[15:0]), //i
    .Sliding_Size                   (Sliding_Size[12:0]                  ), //i
    .Test_Signal                    (SubModule_Test_Signal               ), //o
    .Test_Generate_Period           (SubModule_Test_Generate_Period[15:0]), //i
    .Test_End                       (SubModule_Test_End                  ), //o
    .Raddr_Valid                    (SubModule_Raddr_Valid               ), //o
    .LayerEnd                       (SubModule_LayerEnd                  ), //o
    .SA_Row_Cnt_Valid               (SubModule_SA_Row_Cnt_Valid          ), //o
    .clk                            (clk                                 ), //i
    .reset                          (reset                               )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo (
    .io_push_valid   (streamFifo_io_push_valid          ), //i
    .io_push_ready   (streamFifo_io_push_ready          ), //o
    .io_push_payload (SubModule_mData[63:0]             ), //i
    .io_pop_valid    (streamFifo_io_pop_valid           ), //o
    .io_pop_ready    (axisDataConverter_8_inStream_ready), //i
    .io_pop_payload  (streamFifo_io_pop_payload[63:0]   ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (streamFifo_io_occupancy[4:0]      ), //o
    .io_availability (streamFifo_io_availability[4:0]   ), //o
    .clk             (clk                               ), //i
    .reset           (reset                             )  //i
  );
  AxisDataConverter axisDataConverter_8 (
    .inStream_valid    (streamFifo_io_pop_valid                   ), //i
    .inStream_ready    (axisDataConverter_8_inStream_ready        ), //o
    .inStream_payload  (streamFifo_io_pop_payload[63:0]           ), //i
    .outStream_valid   (axisDataConverter_8_outStream_valid       ), //o
    .outStream_ready   (1'b1                                      ), //i
    .outStream_payload (axisDataConverter_8_outStream_payload[7:0]), //o
    .clk               (clk                                       ), //i
    .reset             (reset                                     )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_1 (
    .io_push_valid   (streamFifo_1_io_push_valid        ), //i
    .io_push_ready   (streamFifo_1_io_push_ready        ), //o
    .io_push_payload (SubModule_mData[63:0]             ), //i
    .io_pop_valid    (streamFifo_1_io_pop_valid         ), //o
    .io_pop_ready    (axisDataConverter_9_inStream_ready), //i
    .io_pop_payload  (streamFifo_1_io_pop_payload[63:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (streamFifo_1_io_occupancy[4:0]    ), //o
    .io_availability (streamFifo_1_io_availability[4:0] ), //o
    .clk             (clk                               ), //i
    .reset           (reset                             )  //i
  );
  AxisDataConverter axisDataConverter_9 (
    .inStream_valid    (streamFifo_1_io_pop_valid                 ), //i
    .inStream_ready    (axisDataConverter_9_inStream_ready        ), //o
    .inStream_payload  (streamFifo_1_io_pop_payload[63:0]         ), //i
    .outStream_valid   (axisDataConverter_9_outStream_valid       ), //o
    .outStream_ready   (1'b1                                      ), //i
    .outStream_payload (axisDataConverter_9_outStream_payload[7:0]), //o
    .clk               (clk                                       ), //i
    .reset             (reset                                     )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_2 (
    .io_push_valid   (streamFifo_2_io_push_valid         ), //i
    .io_push_ready   (streamFifo_2_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_2_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_10_inStream_ready), //i
    .io_pop_payload  (streamFifo_2_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_2_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_2_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_10 (
    .inStream_valid    (streamFifo_2_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_10_inStream_ready        ), //o
    .inStream_payload  (streamFifo_2_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_10_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_10_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_3 (
    .io_push_valid   (streamFifo_3_io_push_valid         ), //i
    .io_push_ready   (streamFifo_3_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_3_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_11_inStream_ready), //i
    .io_pop_payload  (streamFifo_3_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_3_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_3_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_11 (
    .inStream_valid    (streamFifo_3_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_11_inStream_ready        ), //o
    .inStream_payload  (streamFifo_3_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_11_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_11_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_4 (
    .io_push_valid   (streamFifo_4_io_push_valid         ), //i
    .io_push_ready   (streamFifo_4_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_4_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_12_inStream_ready), //i
    .io_pop_payload  (streamFifo_4_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_4_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_4_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_12 (
    .inStream_valid    (streamFifo_4_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_12_inStream_ready        ), //o
    .inStream_payload  (streamFifo_4_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_12_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_12_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_5 (
    .io_push_valid   (streamFifo_5_io_push_valid         ), //i
    .io_push_ready   (streamFifo_5_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_5_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_13_inStream_ready), //i
    .io_pop_payload  (streamFifo_5_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_5_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_5_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_13 (
    .inStream_valid    (streamFifo_5_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_13_inStream_ready        ), //o
    .inStream_payload  (streamFifo_5_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_13_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_13_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_6 (
    .io_push_valid   (streamFifo_6_io_push_valid         ), //i
    .io_push_ready   (streamFifo_6_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_6_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_14_inStream_ready), //i
    .io_pop_payload  (streamFifo_6_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_6_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_6_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_14 (
    .inStream_valid    (streamFifo_6_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_14_inStream_ready        ), //o
    .inStream_payload  (streamFifo_6_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_14_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_14_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  Img2Col_WidthConverter_Fifo streamFifo_7 (
    .io_push_valid   (streamFifo_7_io_push_valid         ), //i
    .io_push_ready   (streamFifo_7_io_push_ready         ), //o
    .io_push_payload (SubModule_mData[63:0]              ), //i
    .io_pop_valid    (streamFifo_7_io_pop_valid          ), //o
    .io_pop_ready    (axisDataConverter_15_inStream_ready), //i
    .io_pop_payload  (streamFifo_7_io_pop_payload[63:0]  ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (streamFifo_7_io_occupancy[4:0]     ), //o
    .io_availability (streamFifo_7_io_availability[4:0]  ), //o
    .clk             (clk                                ), //i
    .reset           (reset                              )  //i
  );
  AxisDataConverter axisDataConverter_15 (
    .inStream_valid    (streamFifo_7_io_pop_valid                  ), //i
    .inStream_ready    (axisDataConverter_15_inStream_ready        ), //o
    .inStream_payload  (streamFifo_7_io_pop_payload[63:0]          ), //i
    .outStream_valid   (axisDataConverter_15_outStream_valid       ), //o
    .outStream_ready   (1'b1                                       ), //i
    .outStream_payload (axisDataConverter_15_outStream_payload[7:0]), //o
    .clk               (clk                                        ), //i
    .reset             (reset                                      )  //i
  );
  assign streamFifo_io_push_valid = (OutData_Switch[0] && SubModule_mValid);
  always @(*) begin
    mData[7 : 0] = SubModule_Img2Col_axisDataConverter_8_outStream_payload_regNext;
    mData[15 : 8] = SubModule_Img2Col_axisDataConverter_9_outStream_payload_regNext;
    mData[23 : 16] = SubModule_Img2Col_axisDataConverter_10_outStream_payload_regNext;
    mData[31 : 24] = SubModule_Img2Col_axisDataConverter_11_outStream_payload_regNext;
    mData[39 : 32] = SubModule_Img2Col_axisDataConverter_12_outStream_payload_regNext;
    mData[47 : 40] = SubModule_Img2Col_axisDataConverter_13_outStream_payload_regNext;
    mData[55 : 48] = SubModule_Img2Col_axisDataConverter_14_outStream_payload_regNext;
    mData[63 : 56] = SubModule_Img2Col_axisDataConverter_15_outStream_payload_regNext;
  end

  always @(*) begin
    mValid[0] = SubModule_Img2Col_axisDataConverter_8_outStream_valid_regNext;
    mValid[1] = SubModule_Img2Col_axisDataConverter_9_outStream_valid_regNext;
    mValid[2] = SubModule_Img2Col_axisDataConverter_10_outStream_valid_regNext;
    mValid[3] = SubModule_Img2Col_axisDataConverter_11_outStream_valid_regNext;
    mValid[4] = SubModule_Img2Col_axisDataConverter_12_outStream_valid_regNext;
    mValid[5] = SubModule_Img2Col_axisDataConverter_13_outStream_valid_regNext;
    mValid[6] = SubModule_Img2Col_axisDataConverter_14_outStream_valid_regNext;
    mValid[7] = SubModule_Img2Col_axisDataConverter_15_outStream_valid_regNext;
  end

  assign streamFifo_1_io_push_valid = (OutData_Switch[1] && SubModule_mValid);
  assign streamFifo_2_io_push_valid = (OutData_Switch[2] && SubModule_mValid);
  assign streamFifo_3_io_push_valid = (OutData_Switch[3] && SubModule_mValid);
  assign streamFifo_4_io_push_valid = (OutData_Switch[4] && SubModule_mValid);
  assign streamFifo_5_io_push_valid = (OutData_Switch[5] && SubModule_mValid);
  assign streamFifo_6_io_push_valid = (OutData_Switch[6] && SubModule_mValid);
  assign streamFifo_7_io_push_valid = (OutData_Switch[7] && SubModule_mValid);
  assign Raddr_Valid = axisDataConverter_8_outStream_valid;
  assign s_axis_s2mm_tready = SubModule_sData_ready;
  assign SubModule_Fifo_Clear = (! streamFifo_io_pop_valid);
  assign LayerEnd = SubModule_Img2Col_SubModule_LayerEnd_delay_3;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      OutData_Switch <= 8'h01;
    end else begin
      if(Switch_Reset) begin
        OutData_Switch <= 8'h01;
      end else begin
        if(SubModule_mValid) begin
          OutData_Switch <= {OutData_Switch[6 : 0],OutData_Switch[7 : 7]};
        end
      end
    end
  end

  always @(posedge clk) begin
    Switch_Reset <= SubModule_SA_Row_Cnt_Valid;
    SubModule_Img2Col_axisDataConverter_8_outStream_payload_regNext <= axisDataConverter_8_outStream_payload;
    SubModule_Img2Col_axisDataConverter_8_outStream_valid_regNext <= axisDataConverter_8_outStream_valid;
    SubModule_Img2Col_axisDataConverter_9_outStream_payload_regNext <= axisDataConverter_9_outStream_payload;
    SubModule_Img2Col_axisDataConverter_9_outStream_valid_regNext <= axisDataConverter_9_outStream_valid;
    SubModule_Img2Col_axisDataConverter_10_outStream_payload_regNext <= axisDataConverter_10_outStream_payload;
    SubModule_Img2Col_axisDataConverter_10_outStream_valid_regNext <= axisDataConverter_10_outStream_valid;
    SubModule_Img2Col_axisDataConverter_11_outStream_payload_regNext <= axisDataConverter_11_outStream_payload;
    SubModule_Img2Col_axisDataConverter_11_outStream_valid_regNext <= axisDataConverter_11_outStream_valid;
    SubModule_Img2Col_axisDataConverter_12_outStream_payload_regNext <= axisDataConverter_12_outStream_payload;
    SubModule_Img2Col_axisDataConverter_12_outStream_valid_regNext <= axisDataConverter_12_outStream_valid;
    SubModule_Img2Col_axisDataConverter_13_outStream_payload_regNext <= axisDataConverter_13_outStream_payload;
    SubModule_Img2Col_axisDataConverter_13_outStream_valid_regNext <= axisDataConverter_13_outStream_valid;
    SubModule_Img2Col_axisDataConverter_14_outStream_payload_regNext <= axisDataConverter_14_outStream_payload;
    SubModule_Img2Col_axisDataConverter_14_outStream_valid_regNext <= axisDataConverter_14_outStream_valid;
    SubModule_Img2Col_axisDataConverter_15_outStream_payload_regNext <= axisDataConverter_15_outStream_payload;
    SubModule_Img2Col_axisDataConverter_15_outStream_valid_regNext <= axisDataConverter_15_outStream_valid;
    SubModule_Img2Col_SubModule_LayerEnd_delay_1 <= SubModule_LayerEnd;
    SubModule_Img2Col_SubModule_LayerEnd_delay_2 <= SubModule_Img2Col_SubModule_LayerEnd_delay_1;
    SubModule_Img2Col_SubModule_LayerEnd_delay_3 <= SubModule_Img2Col_SubModule_LayerEnd_delay_2;
  end


endmodule

module Compute_DataIn_Switch (
  input      [1:0]    Switch,
  input      [63:0]   s0_axis_s2mm_tdata,
  input      [7:0]    s0_axis_s2mm_tkeep,
  input               s0_axis_s2mm_tlast,
  output reg          s0_axis_s2mm_tready,
  input               s0_axis_s2mm_tvalid,
  output reg [63:0]   m_0_axis_mm2s_tdata,
  output     [7:0]    m_0_axis_mm2s_tkeep,
  output reg          m_0_axis_mm2s_tlast,
  input               m_0_axis_mm2s_tready,
  output reg          m_0_axis_mm2s_tvalid,
  output reg [63:0]   m_1_axis_mm2s_tdata,
  output     [7:0]    m_1_axis_mm2s_tkeep,
  output reg          m_1_axis_mm2s_tlast,
  input               m_1_axis_mm2s_tready,
  output reg          m_1_axis_mm2s_tvalid
);

  wire                when_Axis_Switch_l103;
  wire                when_Axis_Switch_l103_1;

  assign m_0_axis_mm2s_tkeep = s0_axis_s2mm_tkeep;
  assign m_1_axis_mm2s_tkeep = s0_axis_s2mm_tkeep;
  always @(*) begin
    s0_axis_s2mm_tready = 1'b0;
    if(when_Axis_Switch_l103) begin
      s0_axis_s2mm_tready = m_0_axis_mm2s_tready;
    end
    if(when_Axis_Switch_l103_1) begin
      s0_axis_s2mm_tready = m_1_axis_mm2s_tready;
    end
  end

  assign when_Axis_Switch_l103 = (Switch == 2'b00);
  always @(*) begin
    if(when_Axis_Switch_l103) begin
      m_0_axis_mm2s_tdata = s0_axis_s2mm_tdata;
    end else begin
      m_0_axis_mm2s_tdata = 64'h0;
    end
  end

  always @(*) begin
    if(when_Axis_Switch_l103) begin
      m_0_axis_mm2s_tlast = s0_axis_s2mm_tlast;
    end else begin
      m_0_axis_mm2s_tlast = 1'b0;
    end
  end

  always @(*) begin
    if(when_Axis_Switch_l103) begin
      m_0_axis_mm2s_tvalid = s0_axis_s2mm_tvalid;
    end else begin
      m_0_axis_mm2s_tvalid = 1'b0;
    end
  end

  assign when_Axis_Switch_l103_1 = (Switch == 2'b01);
  always @(*) begin
    if(when_Axis_Switch_l103_1) begin
      m_1_axis_mm2s_tdata = s0_axis_s2mm_tdata;
    end else begin
      m_1_axis_mm2s_tdata = 64'h0;
    end
  end

  always @(*) begin
    if(when_Axis_Switch_l103_1) begin
      m_1_axis_mm2s_tlast = s0_axis_s2mm_tlast;
    end else begin
      m_1_axis_mm2s_tlast = 1'b0;
    end
  end

  always @(*) begin
    if(when_Axis_Switch_l103_1) begin
      m_1_axis_mm2s_tvalid = s0_axis_s2mm_tvalid;
    end else begin
      m_1_axis_mm2s_tvalid = 1'b0;
    end
  end


endmodule

//ConvOutput_Converter replaced by ConvOutput_Converter

//ConvOutput_Fifo replaced by ConvOutput_Fifo

//ConvOutput_Converter replaced by ConvOutput_Converter

//ConvOutput_Fifo replaced by ConvOutput_Fifo

//ConvOutput_Converter replaced by ConvOutput_Converter

//ConvOutput_Fifo replaced by ConvOutput_Fifo

//ConvOutput_Converter replaced by ConvOutput_Converter

//ConvOutput_Fifo replaced by ConvOutput_Fifo

//ConvOutput_Converter replaced by ConvOutput_Converter

//ConvOutput_Fifo replaced by ConvOutput_Fifo

//ConvOutput_Converter replaced by ConvOutput_Converter

//ConvOutput_Fifo replaced by ConvOutput_Fifo

//ConvOutput_Converter replaced by ConvOutput_Converter

//ConvOutput_Fifo replaced by ConvOutput_Fifo

module ConvOutput_Converter (
  input               inStream_valid,
  output              inStream_ready,
  input      [7:0]    inStream_payload,
  output              outStream_valid,
  input               outStream_ready,
  output     [63:0]   outStream_payload,
  input               clk,
  input               reset
);

  wire       [2:0]    _zz__zz_inStream_ready_1;
  wire       [0:0]    _zz__zz_inStream_ready_1_1;
  wire       [47:0]   _zz__zz_outStream_payload;
  wire       [63:0]   _zz_outStream_payload_1;
  wire       [63:0]   _zz_outStream_payload_2;
  wire                inStream_fire;
  reg                 _zz_inStream_ready;
  reg        [2:0]    _zz_inStream_ready_1;
  reg        [2:0]    _zz_inStream_ready_2;
  wire                _zz_inStream_ready_3;
  reg        [55:0]   _zz_outStream_payload;
  wire                inStream_fire_1;

  assign _zz__zz_inStream_ready_1_1 = _zz_inStream_ready;
  assign _zz__zz_inStream_ready_1 = {2'd0, _zz__zz_inStream_ready_1_1};
  assign _zz__zz_outStream_payload = (_zz_outStream_payload >>> 8);
  assign _zz_outStream_payload_2 = {inStream_payload,_zz_outStream_payload};
  assign _zz_outStream_payload_1 = _zz_outStream_payload_2;
  assign inStream_fire = (inStream_valid && inStream_ready);
  always @(*) begin
    _zz_inStream_ready = 1'b0;
    if(inStream_fire) begin
      _zz_inStream_ready = 1'b1;
    end
  end

  assign _zz_inStream_ready_3 = (_zz_inStream_ready_2 == 3'b111);
  always @(*) begin
    _zz_inStream_ready_1 = (_zz_inStream_ready_2 + _zz__zz_inStream_ready_1);
    if(1'b0) begin
      _zz_inStream_ready_1 = 3'b000;
    end
  end

  assign inStream_fire_1 = (inStream_valid && inStream_ready);
  assign outStream_valid = (inStream_valid && _zz_inStream_ready_3);
  assign outStream_payload = _zz_outStream_payload_1;
  assign inStream_ready = (! ((! outStream_ready) && _zz_inStream_ready_3));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _zz_inStream_ready_2 <= 3'b000;
    end else begin
      _zz_inStream_ready_2 <= _zz_inStream_ready_1;
    end
  end

  always @(posedge clk) begin
    if(inStream_fire_1) begin
      _zz_outStream_payload <= {inStream_payload,_zz__zz_outStream_payload};
    end
  end


endmodule

module ConvOutput_Fifo (
  input               io_push_valid,
  output              io_push_ready,
  input      [63:0]   io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [63:0]   io_pop_payload,
  input               io_flush,
  output     [9:0]    io_occupancy,
  output     [9:0]    io_availability,
  input               clk,
  input               reset
);

  reg        [63:0]   _zz_logic_ram_port0;
  wire       [8:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [8:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [63:0]   _zz_logic_ram_port_1;
  wire       [8:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [8:0]    logic_pushPtr_valueNext;
  reg        [8:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [8:0]    logic_popPtr_valueNext;
  reg        [8:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1122;
  wire       [8:0]    logic_ptrDif;
  reg [63:0] logic_ram [0:511];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {8'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {8'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  assign _zz_logic_ram_port_1 = io_push_payload;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 9'h1ff);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 9'h0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 9'h1ff);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 9'h0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1122 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_pushPtr_value <= 9'h0;
      logic_popPtr_value <= 9'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1122) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module GemmOutput_Ctrl (
  input               ResetCnt,
  input               InData_Cnt_En,
  input               OutData_Cnt_En,
  input      [11:0]   MatrixCol,
  input      [19:0]   MatrixRow,
  output              Fsm_LayerEnd,
  output              Fsm_Data_AllOut,
  output              OutSwitch_Rotate,
  input               clk,
  input               reset
);

  wire       [11:0]   _zz_In_Col_Cnt_valid;
  wire       [19:0]   _zz_In_Row_Cnt_valid;
  wire       [19:0]   _zz_In_Row_Cnt_count_1;
  wire       [8:0]    _zz_Out_Col_Cnt_valid;
  wire       [8:0]    _zz_Out_Col_Cnt_valid_1;
  wire       [19:0]   _zz_Out_Row_Cnt_valid;
  reg        [11:0]   In_Col_Cnt_count;
  wire                In_Col_Cnt_valid;
  wire       [3:0]    _zz_In_Row_Cnt_count;
  reg        [19:0]   In_Row_Cnt_count;
  reg                 In_Row_Cnt_valid;
  reg        [8:0]    Out_Col_Cnt_count;
  wire                Out_Col_Cnt_valid;
  reg        [19:0]   Out_Row_Cnt_count;
  wire                Out_Row_Cnt_valid;

  assign _zz_In_Col_Cnt_valid = (MatrixCol - 12'h001);
  assign _zz_In_Row_Cnt_valid = {16'd0, _zz_In_Row_Cnt_count};
  assign _zz_In_Row_Cnt_count_1 = {16'd0, _zz_In_Row_Cnt_count};
  assign _zz_Out_Col_Cnt_valid = (_zz_Out_Col_Cnt_valid_1 - 9'h001);
  assign _zz_Out_Col_Cnt_valid_1 = (MatrixCol >>> 3);
  assign _zz_Out_Row_Cnt_valid = (MatrixRow - 20'h00001);
  assign In_Col_Cnt_valid = ((In_Col_Cnt_count == _zz_In_Col_Cnt_valid) && InData_Cnt_En);
  assign _zz_In_Row_Cnt_count = 4'b1000;
  always @(*) begin
    In_Row_Cnt_valid = ((In_Row_Cnt_count <= _zz_In_Row_Cnt_valid) && In_Col_Cnt_valid);
    if(ResetCnt) begin
      In_Row_Cnt_valid = 1'b0;
    end
  end

  assign Out_Col_Cnt_valid = ((Out_Col_Cnt_count == _zz_Out_Col_Cnt_valid) && OutData_Cnt_En);
  assign Out_Row_Cnt_valid = ((Out_Row_Cnt_count == _zz_Out_Row_Cnt_valid) && Out_Col_Cnt_valid);
  assign Fsm_Data_AllOut = Out_Row_Cnt_valid;
  assign OutSwitch_Rotate = Out_Col_Cnt_valid;
  assign Fsm_LayerEnd = In_Row_Cnt_valid;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      In_Col_Cnt_count <= 12'h0;
      Out_Col_Cnt_count <= 9'h0;
      Out_Row_Cnt_count <= 20'h0;
    end else begin
      if(InData_Cnt_En) begin
        if(In_Col_Cnt_valid) begin
          In_Col_Cnt_count <= 12'h0;
        end else begin
          In_Col_Cnt_count <= (In_Col_Cnt_count + 12'h001);
        end
      end
      if(OutData_Cnt_En) begin
        if(Out_Col_Cnt_valid) begin
          Out_Col_Cnt_count <= 9'h0;
        end else begin
          Out_Col_Cnt_count <= (Out_Col_Cnt_count + 9'h001);
        end
      end
      if(Out_Col_Cnt_valid) begin
        if(Out_Row_Cnt_valid) begin
          Out_Row_Cnt_count <= 20'h0;
        end else begin
          Out_Row_Cnt_count <= (Out_Row_Cnt_count + 20'h00001);
        end
      end
    end
  end

  always @(posedge clk) begin
    if(In_Col_Cnt_valid) begin
      if(In_Row_Cnt_valid) begin
        In_Row_Cnt_count <= MatrixRow;
      end else begin
        In_Row_Cnt_count <= (In_Row_Cnt_count - _zz_In_Row_Cnt_count_1);
      end
    end
    if(ResetCnt) begin
      In_Row_Cnt_count <= MatrixRow;
    end
  end


endmodule

module ConvOutput_Ctrl (
  input               ResetCnt,
  input               InData_Cnt_En,
  input               OutData_Cnt_En,
  input      [9:0]    OutChannel,
  input      [15:0]   OutFeatureSize,
  output              Fsm_LayerEnd,
  output              Fsm_Data_AllOut,
  output              OutSwitch_Rotate,
  output              OutSwitch_Reset,
  input               clk,
  input               reset
);

  wire       [9:0]    _zz_InChannel_Cnt_valid;
  wire       [9:0]    _zz_InChannel_Cnt_valid_1;
  wire       [15:0]   _zz_In_Col_Cnt_valid;
  wire       [15:0]   _zz_In_Col_Cnt_count_1;
  wire       [19:0]   _zz_In_Row_Cnt_valid;
  wire       [15:0]   _zz_In_Row_Cnt_valid_1;
  wire       [8:0]    _zz_OutChannel_Cnt_valid;
  wire       [6:0]    _zz_OutChannel_Cnt_valid_1;
  wire       [6:0]    _zz_OutChannel_Cnt_valid_2;
  wire       [19:0]   _zz_Out_Col_Cnt_valid;
  wire       [15:0]   _zz_Out_Col_Cnt_valid_1;
  wire       [19:0]   _zz_Out_Row_Cnt_valid;
  wire       [15:0]   _zz_Out_Row_Cnt_valid_1;
  reg        [9:0]    InChannel_Cnt_count;
  wire                InChannel_Cnt_valid;
  wire       [3:0]    _zz_In_Col_Cnt_count;
  reg        [15:0]   In_Col_Cnt_count;
  reg                 In_Col_Cnt_valid;
  reg        [19:0]   In_Row_Cnt_count;
  wire                In_Row_Cnt_valid;
  reg        [8:0]    OutChannel_Cnt_count;
  wire                OutChannel_Cnt_valid;
  reg        [19:0]   Out_Col_Cnt_count;
  wire                Out_Col_Cnt_valid;
  reg        [19:0]   Out_Row_Cnt_count;
  wire                Out_Row_Cnt_valid;

  assign _zz_InChannel_Cnt_valid = (_zz_InChannel_Cnt_valid_1 >>> 0);
  assign _zz_InChannel_Cnt_valid_1 = (OutChannel - 10'h001);
  assign _zz_In_Col_Cnt_valid = {12'd0, _zz_In_Col_Cnt_count};
  assign _zz_In_Col_Cnt_count_1 = {12'd0, _zz_In_Col_Cnt_count};
  assign _zz_In_Row_Cnt_valid_1 = (OutFeatureSize - 16'h0001);
  assign _zz_In_Row_Cnt_valid = {4'd0, _zz_In_Row_Cnt_valid_1};
  assign _zz_OutChannel_Cnt_valid_1 = (_zz_OutChannel_Cnt_valid_2 - 7'h01);
  assign _zz_OutChannel_Cnt_valid = {2'd0, _zz_OutChannel_Cnt_valid_1};
  assign _zz_OutChannel_Cnt_valid_2 = (OutChannel >>> 3);
  assign _zz_Out_Col_Cnt_valid_1 = (OutFeatureSize - 16'h0001);
  assign _zz_Out_Col_Cnt_valid = {4'd0, _zz_Out_Col_Cnt_valid_1};
  assign _zz_Out_Row_Cnt_valid_1 = (OutFeatureSize - 16'h0001);
  assign _zz_Out_Row_Cnt_valid = {4'd0, _zz_Out_Row_Cnt_valid_1};
  assign InChannel_Cnt_valid = ((InChannel_Cnt_count == _zz_InChannel_Cnt_valid) && InData_Cnt_En);
  assign _zz_In_Col_Cnt_count = 4'b1000;
  always @(*) begin
    In_Col_Cnt_valid = ((In_Col_Cnt_count <= _zz_In_Col_Cnt_valid) && InChannel_Cnt_valid);
    if(ResetCnt) begin
      In_Col_Cnt_valid = 1'b0;
    end
  end

  assign In_Row_Cnt_valid = ((In_Row_Cnt_count == _zz_In_Row_Cnt_valid) && In_Col_Cnt_valid);
  assign Fsm_LayerEnd = In_Row_Cnt_valid;
  assign OutChannel_Cnt_valid = ((OutChannel_Cnt_count == _zz_OutChannel_Cnt_valid) && OutData_Cnt_En);
  assign Out_Col_Cnt_valid = ((Out_Col_Cnt_count == _zz_Out_Col_Cnt_valid) && OutChannel_Cnt_valid);
  assign Out_Row_Cnt_valid = ((Out_Row_Cnt_count == _zz_Out_Row_Cnt_valid) && Out_Col_Cnt_valid);
  assign Fsm_Data_AllOut = Out_Row_Cnt_valid;
  assign OutSwitch_Reset = Out_Col_Cnt_valid;
  assign OutSwitch_Rotate = OutChannel_Cnt_valid;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      InChannel_Cnt_count <= 10'h0;
      In_Row_Cnt_count <= 20'h0;
      OutChannel_Cnt_count <= 9'h0;
      Out_Col_Cnt_count <= 20'h0;
      Out_Row_Cnt_count <= 20'h0;
    end else begin
      if(InData_Cnt_En) begin
        if(InChannel_Cnt_valid) begin
          InChannel_Cnt_count <= 10'h0;
        end else begin
          InChannel_Cnt_count <= (InChannel_Cnt_count + 10'h001);
        end
      end
      if(In_Col_Cnt_valid) begin
        if(In_Row_Cnt_valid) begin
          In_Row_Cnt_count <= 20'h0;
        end else begin
          In_Row_Cnt_count <= (In_Row_Cnt_count + 20'h00001);
        end
      end
      if(OutData_Cnt_En) begin
        if(OutChannel_Cnt_valid) begin
          OutChannel_Cnt_count <= 9'h0;
        end else begin
          OutChannel_Cnt_count <= (OutChannel_Cnt_count + 9'h001);
        end
      end
      if(OutChannel_Cnt_valid) begin
        if(Out_Col_Cnt_valid) begin
          Out_Col_Cnt_count <= 20'h0;
        end else begin
          Out_Col_Cnt_count <= (Out_Col_Cnt_count + 20'h00001);
        end
      end
      if(Out_Col_Cnt_valid) begin
        if(Out_Row_Cnt_valid) begin
          Out_Row_Cnt_count <= 20'h0;
        end else begin
          Out_Row_Cnt_count <= (Out_Row_Cnt_count + 20'h00001);
        end
      end
    end
  end

  always @(posedge clk) begin
    if(InChannel_Cnt_valid) begin
      if(In_Col_Cnt_valid) begin
        In_Col_Cnt_count <= OutFeatureSize;
      end else begin
        In_Col_Cnt_count <= (In_Col_Cnt_count - _zz_In_Col_Cnt_count_1);
      end
    end
    if(ResetCnt) begin
      In_Col_Cnt_count <= OutFeatureSize;
    end
  end


endmodule

module Weight_Cache (
  input               start,
  input               sData_valid,
  output              sData_ready,
  input      [63:0]   sData_payload,
  input      [15:0]   Matrix_Row,
  input      [15:0]   Matrix_Col,
  output     [7:0]    mData_0,
  output     [7:0]    mData_1,
  output     [7:0]    mData_2,
  output     [7:0]    mData_3,
  output     [7:0]    mData_4,
  output     [7:0]    mData_5,
  output     [7:0]    mData_6,
  output     [7:0]    mData_7,
  output     [7:0]    mData_8,
  output     [7:0]    mData_9,
  output     [7:0]    mData_10,
  output     [7:0]    mData_11,
  output     [7:0]    mData_12,
  output     [7:0]    mData_13,
  output     [7:0]    mData_14,
  output     [7:0]    mData_15,
  output     [7:0]    mData_16,
  output     [7:0]    mData_17,
  output     [7:0]    mData_18,
  output     [7:0]    mData_19,
  output     [7:0]    mData_20,
  output     [7:0]    mData_21,
  output     [7:0]    mData_22,
  output     [7:0]    mData_23,
  output     [7:0]    mData_24,
  output     [7:0]    mData_25,
  output     [7:0]    mData_26,
  output     [7:0]    mData_27,
  output     [7:0]    mData_28,
  output     [7:0]    mData_29,
  output     [7:0]    mData_30,
  output     [7:0]    mData_31,
  output     [7:0]    mData_32,
  output     [7:0]    mData_33,
  output     [7:0]    mData_34,
  output     [7:0]    mData_35,
  output     [7:0]    mData_36,
  output     [7:0]    mData_37,
  output     [7:0]    mData_38,
  output     [7:0]    mData_39,
  output     [7:0]    mData_40,
  output     [7:0]    mData_41,
  output     [7:0]    mData_42,
  output     [7:0]    mData_43,
  output     [7:0]    mData_44,
  output     [7:0]    mData_45,
  output     [7:0]    mData_46,
  output     [7:0]    mData_47,
  output     [7:0]    mData_48,
  output     [7:0]    mData_49,
  output     [7:0]    mData_50,
  output     [7:0]    mData_51,
  output     [7:0]    mData_52,
  output     [7:0]    mData_53,
  output     [7:0]    mData_54,
  output     [7:0]    mData_55,
  output     [7:0]    mData_56,
  output     [7:0]    mData_57,
  output     [7:0]    mData_58,
  output     [7:0]    mData_59,
  output     [7:0]    mData_60,
  output     [7:0]    mData_61,
  output     [7:0]    mData_62,
  output     [7:0]    mData_63,
  input               Raddr_Valid,
  output              Weight_Cached,
  input               LayerEnd,
  output     [63:0]   MatrixCol_Switch,
  input               clk,
  input               reset
);
  localparam WEIGHT_CACHE_STATUS_IDLE = 4'd1;
  localparam WEIGHT_CACHE_STATUS_INIT = 4'd2;
  localparam WEIGHT_CACHE_STATUS_CACHE_WEIGHT = 4'd4;
  localparam WEIGHT_CACHE_STATUS_SA_COMPUTE = 4'd8;

  wire       [10:0]   xil_SimpleDualBram_addra;
  wire                xil_SimpleDualBram_ena;
  wire       [13:0]   xil_SimpleDualBram_addrb;
  wire       [10:0]   xil_SimpleDualBram_1_addra;
  wire                xil_SimpleDualBram_1_ena;
  wire       [13:0]   xil_SimpleDualBram_1_addrb;
  wire       [10:0]   xil_SimpleDualBram_2_addra;
  wire                xil_SimpleDualBram_2_ena;
  wire       [13:0]   xil_SimpleDualBram_2_addrb;
  wire       [10:0]   xil_SimpleDualBram_3_addra;
  wire                xil_SimpleDualBram_3_ena;
  wire       [13:0]   xil_SimpleDualBram_3_addrb;
  wire       [10:0]   xil_SimpleDualBram_4_addra;
  wire                xil_SimpleDualBram_4_ena;
  wire       [13:0]   xil_SimpleDualBram_4_addrb;
  wire       [10:0]   xil_SimpleDualBram_5_addra;
  wire                xil_SimpleDualBram_5_ena;
  wire       [13:0]   xil_SimpleDualBram_5_addrb;
  wire       [10:0]   xil_SimpleDualBram_6_addra;
  wire                xil_SimpleDualBram_6_ena;
  wire       [13:0]   xil_SimpleDualBram_6_addrb;
  wire       [10:0]   xil_SimpleDualBram_7_addra;
  wire                xil_SimpleDualBram_7_ena;
  wire       [13:0]   xil_SimpleDualBram_7_addrb;
  wire       [10:0]   xil_SimpleDualBram_8_addra;
  wire                xil_SimpleDualBram_8_ena;
  wire       [13:0]   xil_SimpleDualBram_8_addrb;
  wire       [10:0]   xil_SimpleDualBram_9_addra;
  wire                xil_SimpleDualBram_9_ena;
  wire       [13:0]   xil_SimpleDualBram_9_addrb;
  wire       [10:0]   xil_SimpleDualBram_10_addra;
  wire                xil_SimpleDualBram_10_ena;
  wire       [13:0]   xil_SimpleDualBram_10_addrb;
  wire       [10:0]   xil_SimpleDualBram_11_addra;
  wire                xil_SimpleDualBram_11_ena;
  wire       [13:0]   xil_SimpleDualBram_11_addrb;
  wire       [10:0]   xil_SimpleDualBram_12_addra;
  wire                xil_SimpleDualBram_12_ena;
  wire       [13:0]   xil_SimpleDualBram_12_addrb;
  wire       [10:0]   xil_SimpleDualBram_13_addra;
  wire                xil_SimpleDualBram_13_ena;
  wire       [13:0]   xil_SimpleDualBram_13_addrb;
  wire       [10:0]   xil_SimpleDualBram_14_addra;
  wire                xil_SimpleDualBram_14_ena;
  wire       [13:0]   xil_SimpleDualBram_14_addrb;
  wire       [10:0]   xil_SimpleDualBram_15_addra;
  wire                xil_SimpleDualBram_15_ena;
  wire       [13:0]   xil_SimpleDualBram_15_addrb;
  wire       [10:0]   xil_SimpleDualBram_16_addra;
  wire                xil_SimpleDualBram_16_ena;
  wire       [13:0]   xil_SimpleDualBram_16_addrb;
  wire       [10:0]   xil_SimpleDualBram_17_addra;
  wire                xil_SimpleDualBram_17_ena;
  wire       [13:0]   xil_SimpleDualBram_17_addrb;
  wire       [10:0]   xil_SimpleDualBram_18_addra;
  wire                xil_SimpleDualBram_18_ena;
  wire       [13:0]   xil_SimpleDualBram_18_addrb;
  wire       [10:0]   xil_SimpleDualBram_19_addra;
  wire                xil_SimpleDualBram_19_ena;
  wire       [13:0]   xil_SimpleDualBram_19_addrb;
  wire       [10:0]   xil_SimpleDualBram_20_addra;
  wire                xil_SimpleDualBram_20_ena;
  wire       [13:0]   xil_SimpleDualBram_20_addrb;
  wire       [10:0]   xil_SimpleDualBram_21_addra;
  wire                xil_SimpleDualBram_21_ena;
  wire       [13:0]   xil_SimpleDualBram_21_addrb;
  wire       [10:0]   xil_SimpleDualBram_22_addra;
  wire                xil_SimpleDualBram_22_ena;
  wire       [13:0]   xil_SimpleDualBram_22_addrb;
  wire       [10:0]   xil_SimpleDualBram_23_addra;
  wire                xil_SimpleDualBram_23_ena;
  wire       [13:0]   xil_SimpleDualBram_23_addrb;
  wire       [10:0]   xil_SimpleDualBram_24_addra;
  wire                xil_SimpleDualBram_24_ena;
  wire       [13:0]   xil_SimpleDualBram_24_addrb;
  wire       [10:0]   xil_SimpleDualBram_25_addra;
  wire                xil_SimpleDualBram_25_ena;
  wire       [13:0]   xil_SimpleDualBram_25_addrb;
  wire       [10:0]   xil_SimpleDualBram_26_addra;
  wire                xil_SimpleDualBram_26_ena;
  wire       [13:0]   xil_SimpleDualBram_26_addrb;
  wire       [10:0]   xil_SimpleDualBram_27_addra;
  wire                xil_SimpleDualBram_27_ena;
  wire       [13:0]   xil_SimpleDualBram_27_addrb;
  wire       [10:0]   xil_SimpleDualBram_28_addra;
  wire                xil_SimpleDualBram_28_ena;
  wire       [13:0]   xil_SimpleDualBram_28_addrb;
  wire       [10:0]   xil_SimpleDualBram_29_addra;
  wire                xil_SimpleDualBram_29_ena;
  wire       [13:0]   xil_SimpleDualBram_29_addrb;
  wire       [10:0]   xil_SimpleDualBram_30_addra;
  wire                xil_SimpleDualBram_30_ena;
  wire       [13:0]   xil_SimpleDualBram_30_addrb;
  wire       [10:0]   xil_SimpleDualBram_31_addra;
  wire                xil_SimpleDualBram_31_ena;
  wire       [13:0]   xil_SimpleDualBram_31_addrb;
  wire       [10:0]   xil_SimpleDualBram_32_addra;
  wire                xil_SimpleDualBram_32_ena;
  wire       [13:0]   xil_SimpleDualBram_32_addrb;
  wire       [10:0]   xil_SimpleDualBram_33_addra;
  wire                xil_SimpleDualBram_33_ena;
  wire       [13:0]   xil_SimpleDualBram_33_addrb;
  wire       [10:0]   xil_SimpleDualBram_34_addra;
  wire                xil_SimpleDualBram_34_ena;
  wire       [13:0]   xil_SimpleDualBram_34_addrb;
  wire       [10:0]   xil_SimpleDualBram_35_addra;
  wire                xil_SimpleDualBram_35_ena;
  wire       [13:0]   xil_SimpleDualBram_35_addrb;
  wire       [10:0]   xil_SimpleDualBram_36_addra;
  wire                xil_SimpleDualBram_36_ena;
  wire       [13:0]   xil_SimpleDualBram_36_addrb;
  wire       [10:0]   xil_SimpleDualBram_37_addra;
  wire                xil_SimpleDualBram_37_ena;
  wire       [13:0]   xil_SimpleDualBram_37_addrb;
  wire       [10:0]   xil_SimpleDualBram_38_addra;
  wire                xil_SimpleDualBram_38_ena;
  wire       [13:0]   xil_SimpleDualBram_38_addrb;
  wire       [10:0]   xil_SimpleDualBram_39_addra;
  wire                xil_SimpleDualBram_39_ena;
  wire       [13:0]   xil_SimpleDualBram_39_addrb;
  wire       [10:0]   xil_SimpleDualBram_40_addra;
  wire                xil_SimpleDualBram_40_ena;
  wire       [13:0]   xil_SimpleDualBram_40_addrb;
  wire       [10:0]   xil_SimpleDualBram_41_addra;
  wire                xil_SimpleDualBram_41_ena;
  wire       [13:0]   xil_SimpleDualBram_41_addrb;
  wire       [10:0]   xil_SimpleDualBram_42_addra;
  wire                xil_SimpleDualBram_42_ena;
  wire       [13:0]   xil_SimpleDualBram_42_addrb;
  wire       [10:0]   xil_SimpleDualBram_43_addra;
  wire                xil_SimpleDualBram_43_ena;
  wire       [13:0]   xil_SimpleDualBram_43_addrb;
  wire       [10:0]   xil_SimpleDualBram_44_addra;
  wire                xil_SimpleDualBram_44_ena;
  wire       [13:0]   xil_SimpleDualBram_44_addrb;
  wire       [10:0]   xil_SimpleDualBram_45_addra;
  wire                xil_SimpleDualBram_45_ena;
  wire       [13:0]   xil_SimpleDualBram_45_addrb;
  wire       [10:0]   xil_SimpleDualBram_46_addra;
  wire                xil_SimpleDualBram_46_ena;
  wire       [13:0]   xil_SimpleDualBram_46_addrb;
  wire       [10:0]   xil_SimpleDualBram_47_addra;
  wire                xil_SimpleDualBram_47_ena;
  wire       [13:0]   xil_SimpleDualBram_47_addrb;
  wire       [10:0]   xil_SimpleDualBram_48_addra;
  wire                xil_SimpleDualBram_48_ena;
  wire       [13:0]   xil_SimpleDualBram_48_addrb;
  wire       [10:0]   xil_SimpleDualBram_49_addra;
  wire                xil_SimpleDualBram_49_ena;
  wire       [13:0]   xil_SimpleDualBram_49_addrb;
  wire       [10:0]   xil_SimpleDualBram_50_addra;
  wire                xil_SimpleDualBram_50_ena;
  wire       [13:0]   xil_SimpleDualBram_50_addrb;
  wire       [10:0]   xil_SimpleDualBram_51_addra;
  wire                xil_SimpleDualBram_51_ena;
  wire       [13:0]   xil_SimpleDualBram_51_addrb;
  wire       [10:0]   xil_SimpleDualBram_52_addra;
  wire                xil_SimpleDualBram_52_ena;
  wire       [13:0]   xil_SimpleDualBram_52_addrb;
  wire       [10:0]   xil_SimpleDualBram_53_addra;
  wire                xil_SimpleDualBram_53_ena;
  wire       [13:0]   xil_SimpleDualBram_53_addrb;
  wire       [10:0]   xil_SimpleDualBram_54_addra;
  wire                xil_SimpleDualBram_54_ena;
  wire       [13:0]   xil_SimpleDualBram_54_addrb;
  wire       [10:0]   xil_SimpleDualBram_55_addra;
  wire                xil_SimpleDualBram_55_ena;
  wire       [13:0]   xil_SimpleDualBram_55_addrb;
  wire       [10:0]   xil_SimpleDualBram_56_addra;
  wire                xil_SimpleDualBram_56_ena;
  wire       [13:0]   xil_SimpleDualBram_56_addrb;
  wire       [10:0]   xil_SimpleDualBram_57_addra;
  wire                xil_SimpleDualBram_57_ena;
  wire       [13:0]   xil_SimpleDualBram_57_addrb;
  wire       [10:0]   xil_SimpleDualBram_58_addra;
  wire                xil_SimpleDualBram_58_ena;
  wire       [13:0]   xil_SimpleDualBram_58_addrb;
  wire       [10:0]   xil_SimpleDualBram_59_addra;
  wire                xil_SimpleDualBram_59_ena;
  wire       [13:0]   xil_SimpleDualBram_59_addrb;
  wire       [10:0]   xil_SimpleDualBram_60_addra;
  wire                xil_SimpleDualBram_60_ena;
  wire       [13:0]   xil_SimpleDualBram_60_addrb;
  wire       [10:0]   xil_SimpleDualBram_61_addra;
  wire                xil_SimpleDualBram_61_ena;
  wire       [13:0]   xil_SimpleDualBram_61_addrb;
  wire       [10:0]   xil_SimpleDualBram_62_addra;
  wire                xil_SimpleDualBram_62_ena;
  wire       [13:0]   xil_SimpleDualBram_62_addrb;
  wire       [10:0]   xil_SimpleDualBram_63_addra;
  wire                xil_SimpleDualBram_63_ena;
  wire       [13:0]   xil_SimpleDualBram_63_addrb;
  wire       [7:0]    xil_SimpleDualBram_doutb;
  wire       [7:0]    xil_SimpleDualBram_1_doutb;
  wire       [7:0]    xil_SimpleDualBram_2_doutb;
  wire       [7:0]    xil_SimpleDualBram_3_doutb;
  wire       [7:0]    xil_SimpleDualBram_4_doutb;
  wire       [7:0]    xil_SimpleDualBram_5_doutb;
  wire       [7:0]    xil_SimpleDualBram_6_doutb;
  wire       [7:0]    xil_SimpleDualBram_7_doutb;
  wire       [7:0]    xil_SimpleDualBram_8_doutb;
  wire       [7:0]    xil_SimpleDualBram_9_doutb;
  wire       [7:0]    xil_SimpleDualBram_10_doutb;
  wire       [7:0]    xil_SimpleDualBram_11_doutb;
  wire       [7:0]    xil_SimpleDualBram_12_doutb;
  wire       [7:0]    xil_SimpleDualBram_13_doutb;
  wire       [7:0]    xil_SimpleDualBram_14_doutb;
  wire       [7:0]    xil_SimpleDualBram_15_doutb;
  wire       [7:0]    xil_SimpleDualBram_16_doutb;
  wire       [7:0]    xil_SimpleDualBram_17_doutb;
  wire       [7:0]    xil_SimpleDualBram_18_doutb;
  wire       [7:0]    xil_SimpleDualBram_19_doutb;
  wire       [7:0]    xil_SimpleDualBram_20_doutb;
  wire       [7:0]    xil_SimpleDualBram_21_doutb;
  wire       [7:0]    xil_SimpleDualBram_22_doutb;
  wire       [7:0]    xil_SimpleDualBram_23_doutb;
  wire       [7:0]    xil_SimpleDualBram_24_doutb;
  wire       [7:0]    xil_SimpleDualBram_25_doutb;
  wire       [7:0]    xil_SimpleDualBram_26_doutb;
  wire       [7:0]    xil_SimpleDualBram_27_doutb;
  wire       [7:0]    xil_SimpleDualBram_28_doutb;
  wire       [7:0]    xil_SimpleDualBram_29_doutb;
  wire       [7:0]    xil_SimpleDualBram_30_doutb;
  wire       [7:0]    xil_SimpleDualBram_31_doutb;
  wire       [7:0]    xil_SimpleDualBram_32_doutb;
  wire       [7:0]    xil_SimpleDualBram_33_doutb;
  wire       [7:0]    xil_SimpleDualBram_34_doutb;
  wire       [7:0]    xil_SimpleDualBram_35_doutb;
  wire       [7:0]    xil_SimpleDualBram_36_doutb;
  wire       [7:0]    xil_SimpleDualBram_37_doutb;
  wire       [7:0]    xil_SimpleDualBram_38_doutb;
  wire       [7:0]    xil_SimpleDualBram_39_doutb;
  wire       [7:0]    xil_SimpleDualBram_40_doutb;
  wire       [7:0]    xil_SimpleDualBram_41_doutb;
  wire       [7:0]    xil_SimpleDualBram_42_doutb;
  wire       [7:0]    xil_SimpleDualBram_43_doutb;
  wire       [7:0]    xil_SimpleDualBram_44_doutb;
  wire       [7:0]    xil_SimpleDualBram_45_doutb;
  wire       [7:0]    xil_SimpleDualBram_46_doutb;
  wire       [7:0]    xil_SimpleDualBram_47_doutb;
  wire       [7:0]    xil_SimpleDualBram_48_doutb;
  wire       [7:0]    xil_SimpleDualBram_49_doutb;
  wire       [7:0]    xil_SimpleDualBram_50_doutb;
  wire       [7:0]    xil_SimpleDualBram_51_doutb;
  wire       [7:0]    xil_SimpleDualBram_52_doutb;
  wire       [7:0]    xil_SimpleDualBram_53_doutb;
  wire       [7:0]    xil_SimpleDualBram_54_doutb;
  wire       [7:0]    xil_SimpleDualBram_55_doutb;
  wire       [7:0]    xil_SimpleDualBram_56_doutb;
  wire       [7:0]    xil_SimpleDualBram_57_doutb;
  wire       [7:0]    xil_SimpleDualBram_58_doutb;
  wire       [7:0]    xil_SimpleDualBram_59_doutb;
  wire       [7:0]    xil_SimpleDualBram_60_doutb;
  wire       [7:0]    xil_SimpleDualBram_61_doutb;
  wire       [7:0]    xil_SimpleDualBram_62_doutb;
  wire       [7:0]    xil_SimpleDualBram_63_doutb;
  wire       [15:0]   _zz_In_Row_Cnt_valid;
  wire       [12:0]   _zz_In_Row_Cnt_valid_1;
  wire       [15:0]   _zz_In_Col_Cnt_valid;
  wire       [15:0]   _zz_OutRow_Cnt_valid;
  wire       [15:0]   _zz_OutCol_Cnt_valid;
  wire       [15:0]   _zz_OutCol_Cnt_count_1;
  wire       [15:0]   _zz_Write_Row_Base_Addr;
  wire       [15:0]   _zz_addra;
  wire       [15:0]   _zz_addrb;
  wire       [0:0]    _zz_ena;
  wire       [15:0]   _zz_addra_1;
  wire       [15:0]   _zz_addrb_1;
  wire       [0:0]    _zz_ena_1;
  wire       [15:0]   _zz_addra_2;
  wire       [15:0]   _zz_addrb_2;
  wire       [0:0]    _zz_ena_2;
  wire       [15:0]   _zz_addra_3;
  wire       [15:0]   _zz_addrb_3;
  wire       [0:0]    _zz_ena_3;
  wire       [15:0]   _zz_addra_4;
  wire       [15:0]   _zz_addrb_4;
  wire       [0:0]    _zz_ena_4;
  wire       [15:0]   _zz_addra_5;
  wire       [15:0]   _zz_addrb_5;
  wire       [0:0]    _zz_ena_5;
  wire       [15:0]   _zz_addra_6;
  wire       [15:0]   _zz_addrb_6;
  wire       [0:0]    _zz_ena_6;
  wire       [15:0]   _zz_addra_7;
  wire       [15:0]   _zz_addrb_7;
  wire       [0:0]    _zz_ena_7;
  wire       [15:0]   _zz_addra_8;
  wire       [15:0]   _zz_addrb_8;
  wire       [0:0]    _zz_ena_8;
  wire       [15:0]   _zz_addra_9;
  wire       [15:0]   _zz_addrb_9;
  wire       [0:0]    _zz_ena_9;
  wire       [15:0]   _zz_addra_10;
  wire       [15:0]   _zz_addrb_10;
  wire       [0:0]    _zz_ena_10;
  wire       [15:0]   _zz_addra_11;
  wire       [15:0]   _zz_addrb_11;
  wire       [0:0]    _zz_ena_11;
  wire       [15:0]   _zz_addra_12;
  wire       [15:0]   _zz_addrb_12;
  wire       [0:0]    _zz_ena_12;
  wire       [15:0]   _zz_addra_13;
  wire       [15:0]   _zz_addrb_13;
  wire       [0:0]    _zz_ena_13;
  wire       [15:0]   _zz_addra_14;
  wire       [15:0]   _zz_addrb_14;
  wire       [0:0]    _zz_ena_14;
  wire       [15:0]   _zz_addra_15;
  wire       [15:0]   _zz_addrb_15;
  wire       [0:0]    _zz_ena_15;
  wire       [15:0]   _zz_addra_16;
  wire       [15:0]   _zz_addrb_16;
  wire       [0:0]    _zz_ena_16;
  wire       [15:0]   _zz_addra_17;
  wire       [15:0]   _zz_addrb_17;
  wire       [0:0]    _zz_ena_17;
  wire       [15:0]   _zz_addra_18;
  wire       [15:0]   _zz_addrb_18;
  wire       [0:0]    _zz_ena_18;
  wire       [15:0]   _zz_addra_19;
  wire       [15:0]   _zz_addrb_19;
  wire       [0:0]    _zz_ena_19;
  wire       [15:0]   _zz_addra_20;
  wire       [15:0]   _zz_addrb_20;
  wire       [0:0]    _zz_ena_20;
  wire       [15:0]   _zz_addra_21;
  wire       [15:0]   _zz_addrb_21;
  wire       [0:0]    _zz_ena_21;
  wire       [15:0]   _zz_addra_22;
  wire       [15:0]   _zz_addrb_22;
  wire       [0:0]    _zz_ena_22;
  wire       [15:0]   _zz_addra_23;
  wire       [15:0]   _zz_addrb_23;
  wire       [0:0]    _zz_ena_23;
  wire       [15:0]   _zz_addra_24;
  wire       [15:0]   _zz_addrb_24;
  wire       [0:0]    _zz_ena_24;
  wire       [15:0]   _zz_addra_25;
  wire       [15:0]   _zz_addrb_25;
  wire       [0:0]    _zz_ena_25;
  wire       [15:0]   _zz_addra_26;
  wire       [15:0]   _zz_addrb_26;
  wire       [0:0]    _zz_ena_26;
  wire       [15:0]   _zz_addra_27;
  wire       [15:0]   _zz_addrb_27;
  wire       [0:0]    _zz_ena_27;
  wire       [15:0]   _zz_addra_28;
  wire       [15:0]   _zz_addrb_28;
  wire       [0:0]    _zz_ena_28;
  wire       [15:0]   _zz_addra_29;
  wire       [15:0]   _zz_addrb_29;
  wire       [0:0]    _zz_ena_29;
  wire       [15:0]   _zz_addra_30;
  wire       [15:0]   _zz_addrb_30;
  wire       [0:0]    _zz_ena_30;
  wire       [15:0]   _zz_addra_31;
  wire       [15:0]   _zz_addrb_31;
  wire       [0:0]    _zz_ena_31;
  wire       [15:0]   _zz_addra_32;
  wire       [15:0]   _zz_addrb_32;
  wire       [0:0]    _zz_ena_32;
  wire       [15:0]   _zz_addra_33;
  wire       [15:0]   _zz_addrb_33;
  wire       [0:0]    _zz_ena_33;
  wire       [15:0]   _zz_addra_34;
  wire       [15:0]   _zz_addrb_34;
  wire       [0:0]    _zz_ena_34;
  wire       [15:0]   _zz_addra_35;
  wire       [15:0]   _zz_addrb_35;
  wire       [0:0]    _zz_ena_35;
  wire       [15:0]   _zz_addra_36;
  wire       [15:0]   _zz_addrb_36;
  wire       [0:0]    _zz_ena_36;
  wire       [15:0]   _zz_addra_37;
  wire       [15:0]   _zz_addrb_37;
  wire       [0:0]    _zz_ena_37;
  wire       [15:0]   _zz_addra_38;
  wire       [15:0]   _zz_addrb_38;
  wire       [0:0]    _zz_ena_38;
  wire       [15:0]   _zz_addra_39;
  wire       [15:0]   _zz_addrb_39;
  wire       [0:0]    _zz_ena_39;
  wire       [15:0]   _zz_addra_40;
  wire       [15:0]   _zz_addrb_40;
  wire       [0:0]    _zz_ena_40;
  wire       [15:0]   _zz_addra_41;
  wire       [15:0]   _zz_addrb_41;
  wire       [0:0]    _zz_ena_41;
  wire       [15:0]   _zz_addra_42;
  wire       [15:0]   _zz_addrb_42;
  wire       [0:0]    _zz_ena_42;
  wire       [15:0]   _zz_addra_43;
  wire       [15:0]   _zz_addrb_43;
  wire       [0:0]    _zz_ena_43;
  wire       [15:0]   _zz_addra_44;
  wire       [15:0]   _zz_addrb_44;
  wire       [0:0]    _zz_ena_44;
  wire       [15:0]   _zz_addra_45;
  wire       [15:0]   _zz_addrb_45;
  wire       [0:0]    _zz_ena_45;
  wire       [15:0]   _zz_addra_46;
  wire       [15:0]   _zz_addrb_46;
  wire       [0:0]    _zz_ena_46;
  wire       [15:0]   _zz_addra_47;
  wire       [15:0]   _zz_addrb_47;
  wire       [0:0]    _zz_ena_47;
  wire       [15:0]   _zz_addra_48;
  wire       [15:0]   _zz_addrb_48;
  wire       [0:0]    _zz_ena_48;
  wire       [15:0]   _zz_addra_49;
  wire       [15:0]   _zz_addrb_49;
  wire       [0:0]    _zz_ena_49;
  wire       [15:0]   _zz_addra_50;
  wire       [15:0]   _zz_addrb_50;
  wire       [0:0]    _zz_ena_50;
  wire       [15:0]   _zz_addra_51;
  wire       [15:0]   _zz_addrb_51;
  wire       [0:0]    _zz_ena_51;
  wire       [15:0]   _zz_addra_52;
  wire       [15:0]   _zz_addrb_52;
  wire       [0:0]    _zz_ena_52;
  wire       [15:0]   _zz_addra_53;
  wire       [15:0]   _zz_addrb_53;
  wire       [0:0]    _zz_ena_53;
  wire       [15:0]   _zz_addra_54;
  wire       [15:0]   _zz_addrb_54;
  wire       [0:0]    _zz_ena_54;
  wire       [15:0]   _zz_addra_55;
  wire       [15:0]   _zz_addrb_55;
  wire       [0:0]    _zz_ena_55;
  wire       [15:0]   _zz_addra_56;
  wire       [15:0]   _zz_addrb_56;
  wire       [0:0]    _zz_ena_56;
  wire       [15:0]   _zz_addra_57;
  wire       [15:0]   _zz_addrb_57;
  wire       [0:0]    _zz_ena_57;
  wire       [15:0]   _zz_addra_58;
  wire       [15:0]   _zz_addrb_58;
  wire       [0:0]    _zz_ena_58;
  wire       [15:0]   _zz_addra_59;
  wire       [15:0]   _zz_addrb_59;
  wire       [0:0]    _zz_ena_59;
  wire       [15:0]   _zz_addra_60;
  wire       [15:0]   _zz_addrb_60;
  wire       [0:0]    _zz_ena_60;
  wire       [15:0]   _zz_addra_61;
  wire       [15:0]   _zz_addrb_61;
  wire       [0:0]    _zz_ena_61;
  wire       [15:0]   _zz_addra_62;
  wire       [15:0]   _zz_addrb_62;
  wire       [0:0]    _zz_ena_62;
  wire       [15:0]   _zz_addra_63;
  wire       [15:0]   _zz_addrb_63;
  wire       [0:0]    _zz_ena_63;
  reg                 start_regNext;
  wire                when_SA3D_WeightCache_l33;
  reg        [3:0]    Fsm_currentState;
  reg        [3:0]    Fsm_nextState;
  wire                Fsm_Init_End;
  wire                Fsm_Weight_All_Cached;
  wire                Fsm_SA_Computed;
  wire                when_WaCounter_l19;
  reg        [2:0]    Init_Count_count;
  reg                 Init_Count_valid;
  wire                when_WaCounter_l14;
  reg        [63:0]   InData_Switch;
  wire       [12:0]   Matrix_In_MaxCnt;
  wire                sData_fire;
  reg        [15:0]   In_Row_Cnt_count;
  wire                In_Row_Cnt_valid;
  reg        [15:0]   In_Col_Cnt_count;
  wire                In_Col_Cnt_valid;
  reg        [15:0]   Read_Row_Base_Addr;
  reg        [15:0]   Write_Row_Base_Addr;
  wire                when_WaCounter_l40;
  reg        [15:0]   OutRow_Cnt_count;
  wire                OutRow_Cnt_valid;
  wire       [6:0]    _zz_OutCol_Cnt_count;
  reg        [15:0]   OutCol_Cnt_count;
  reg                 OutCol_Cnt_valid;
  reg        [5:0]    Col_In_8_Cnt_count;
  reg                 Col_In_8_Cnt_valid;
  wire                when_SA3D_WeightCache_l131;
  wire                when_SA3D_WeightCache_l136;
  wire                sData_fire_1;
  wire                sData_fire_2;
  wire                sData_fire_3;
  wire                sData_fire_4;
  wire                sData_fire_5;
  wire                sData_fire_6;
  wire                sData_fire_7;
  wire                sData_fire_8;
  wire                sData_fire_9;
  wire                sData_fire_10;
  wire                sData_fire_11;
  wire                sData_fire_12;
  wire                sData_fire_13;
  wire                sData_fire_14;
  wire                sData_fire_15;
  wire                sData_fire_16;
  wire                sData_fire_17;
  wire                sData_fire_18;
  wire                sData_fire_19;
  wire                sData_fire_20;
  wire                sData_fire_21;
  wire                sData_fire_22;
  wire                sData_fire_23;
  wire                sData_fire_24;
  wire                sData_fire_25;
  wire                sData_fire_26;
  wire                sData_fire_27;
  wire                sData_fire_28;
  wire                sData_fire_29;
  wire                sData_fire_30;
  wire                sData_fire_31;
  wire                sData_fire_32;
  wire                sData_fire_33;
  wire                sData_fire_34;
  wire                sData_fire_35;
  wire                sData_fire_36;
  wire                sData_fire_37;
  wire                sData_fire_38;
  wire                sData_fire_39;
  wire                sData_fire_40;
  wire                sData_fire_41;
  wire                sData_fire_42;
  wire                sData_fire_43;
  wire                sData_fire_44;
  wire                sData_fire_45;
  wire                sData_fire_46;
  wire                sData_fire_47;
  wire                sData_fire_48;
  wire                sData_fire_49;
  wire                sData_fire_50;
  wire                sData_fire_51;
  wire                sData_fire_52;
  wire                sData_fire_53;
  wire                sData_fire_54;
  wire                sData_fire_55;
  wire                sData_fire_56;
  wire                sData_fire_57;
  wire                sData_fire_58;
  wire                sData_fire_59;
  wire                sData_fire_60;
  wire                sData_fire_61;
  wire                sData_fire_62;
  wire                sData_fire_63;
  wire                sData_fire_64;
  reg        [63:0]   MatrixCol_Switch_1;
  reg        [63:0]   MatrixCol_Switch_1_regNext;
  `ifndef SYNTHESIS
  reg [95:0] Fsm_currentState_string;
  reg [95:0] Fsm_nextState_string;
  `endif


  assign _zz_In_Row_Cnt_valid_1 = (Matrix_In_MaxCnt - 13'h0001);
  assign _zz_In_Row_Cnt_valid = {3'd0, _zz_In_Row_Cnt_valid_1};
  assign _zz_In_Col_Cnt_valid = (Matrix_Col - 16'h0001);
  assign _zz_OutRow_Cnt_valid = (Matrix_Row - 16'h0001);
  assign _zz_OutCol_Cnt_valid = {9'd0, _zz_OutCol_Cnt_count};
  assign _zz_OutCol_Cnt_count_1 = {9'd0, _zz_OutCol_Cnt_count};
  assign _zz_Write_Row_Base_Addr = {3'd0, Matrix_In_MaxCnt};
  assign _zz_addra = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena = InData_Switch[0 : 0];
  assign _zz_addra_1 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_1 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_1 = InData_Switch[1 : 1];
  assign _zz_addra_2 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_2 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_2 = InData_Switch[2 : 2];
  assign _zz_addra_3 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_3 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_3 = InData_Switch[3 : 3];
  assign _zz_addra_4 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_4 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_4 = InData_Switch[4 : 4];
  assign _zz_addra_5 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_5 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_5 = InData_Switch[5 : 5];
  assign _zz_addra_6 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_6 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_6 = InData_Switch[6 : 6];
  assign _zz_addra_7 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_7 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_7 = InData_Switch[7 : 7];
  assign _zz_addra_8 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_8 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_8 = InData_Switch[8 : 8];
  assign _zz_addra_9 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_9 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_9 = InData_Switch[9 : 9];
  assign _zz_addra_10 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_10 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_10 = InData_Switch[10 : 10];
  assign _zz_addra_11 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_11 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_11 = InData_Switch[11 : 11];
  assign _zz_addra_12 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_12 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_12 = InData_Switch[12 : 12];
  assign _zz_addra_13 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_13 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_13 = InData_Switch[13 : 13];
  assign _zz_addra_14 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_14 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_14 = InData_Switch[14 : 14];
  assign _zz_addra_15 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_15 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_15 = InData_Switch[15 : 15];
  assign _zz_addra_16 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_16 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_16 = InData_Switch[16 : 16];
  assign _zz_addra_17 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_17 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_17 = InData_Switch[17 : 17];
  assign _zz_addra_18 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_18 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_18 = InData_Switch[18 : 18];
  assign _zz_addra_19 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_19 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_19 = InData_Switch[19 : 19];
  assign _zz_addra_20 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_20 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_20 = InData_Switch[20 : 20];
  assign _zz_addra_21 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_21 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_21 = InData_Switch[21 : 21];
  assign _zz_addra_22 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_22 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_22 = InData_Switch[22 : 22];
  assign _zz_addra_23 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_23 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_23 = InData_Switch[23 : 23];
  assign _zz_addra_24 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_24 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_24 = InData_Switch[24 : 24];
  assign _zz_addra_25 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_25 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_25 = InData_Switch[25 : 25];
  assign _zz_addra_26 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_26 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_26 = InData_Switch[26 : 26];
  assign _zz_addra_27 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_27 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_27 = InData_Switch[27 : 27];
  assign _zz_addra_28 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_28 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_28 = InData_Switch[28 : 28];
  assign _zz_addra_29 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_29 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_29 = InData_Switch[29 : 29];
  assign _zz_addra_30 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_30 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_30 = InData_Switch[30 : 30];
  assign _zz_addra_31 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_31 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_31 = InData_Switch[31 : 31];
  assign _zz_addra_32 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_32 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_32 = InData_Switch[32 : 32];
  assign _zz_addra_33 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_33 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_33 = InData_Switch[33 : 33];
  assign _zz_addra_34 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_34 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_34 = InData_Switch[34 : 34];
  assign _zz_addra_35 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_35 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_35 = InData_Switch[35 : 35];
  assign _zz_addra_36 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_36 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_36 = InData_Switch[36 : 36];
  assign _zz_addra_37 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_37 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_37 = InData_Switch[37 : 37];
  assign _zz_addra_38 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_38 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_38 = InData_Switch[38 : 38];
  assign _zz_addra_39 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_39 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_39 = InData_Switch[39 : 39];
  assign _zz_addra_40 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_40 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_40 = InData_Switch[40 : 40];
  assign _zz_addra_41 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_41 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_41 = InData_Switch[41 : 41];
  assign _zz_addra_42 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_42 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_42 = InData_Switch[42 : 42];
  assign _zz_addra_43 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_43 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_43 = InData_Switch[43 : 43];
  assign _zz_addra_44 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_44 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_44 = InData_Switch[44 : 44];
  assign _zz_addra_45 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_45 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_45 = InData_Switch[45 : 45];
  assign _zz_addra_46 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_46 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_46 = InData_Switch[46 : 46];
  assign _zz_addra_47 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_47 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_47 = InData_Switch[47 : 47];
  assign _zz_addra_48 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_48 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_48 = InData_Switch[48 : 48];
  assign _zz_addra_49 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_49 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_49 = InData_Switch[49 : 49];
  assign _zz_addra_50 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_50 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_50 = InData_Switch[50 : 50];
  assign _zz_addra_51 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_51 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_51 = InData_Switch[51 : 51];
  assign _zz_addra_52 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_52 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_52 = InData_Switch[52 : 52];
  assign _zz_addra_53 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_53 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_53 = InData_Switch[53 : 53];
  assign _zz_addra_54 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_54 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_54 = InData_Switch[54 : 54];
  assign _zz_addra_55 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_55 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_55 = InData_Switch[55 : 55];
  assign _zz_addra_56 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_56 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_56 = InData_Switch[56 : 56];
  assign _zz_addra_57 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_57 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_57 = InData_Switch[57 : 57];
  assign _zz_addra_58 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_58 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_58 = InData_Switch[58 : 58];
  assign _zz_addra_59 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_59 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_59 = InData_Switch[59 : 59];
  assign _zz_addra_60 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_60 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_60 = InData_Switch[60 : 60];
  assign _zz_addra_61 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_61 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_61 = InData_Switch[61 : 61];
  assign _zz_addra_62 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_62 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_62 = InData_Switch[62 : 62];
  assign _zz_addra_63 = (In_Row_Cnt_count + Write_Row_Base_Addr);
  assign _zz_addrb_63 = (Read_Row_Base_Addr + OutRow_Cnt_count);
  assign _zz_ena_63 = InData_Switch[63 : 63];
  Weight_Bram xil_SimpleDualBram (
    .clka  (clk                           ), //i
    .addra (xil_SimpleDualBram_addra[10:0]), //i
    .dina  (sData_payload[63:0]           ), //i
    .ena   (xil_SimpleDualBram_ena        ), //i
    .wea   (1'b1                          ), //i
    .addrb (xil_SimpleDualBram_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_doutb[7:0] ), //o
    .clkb  (clk                           )  //i
  );
  Weight_Bram xil_SimpleDualBram_1 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_1_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_1_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_1_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_1_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_2 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_2_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_2_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_2_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_2_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_3 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_3_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_3_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_3_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_3_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_4 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_4_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_4_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_4_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_4_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_5 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_5_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_5_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_5_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_5_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_6 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_6_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_6_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_6_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_6_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_7 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_7_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_7_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_7_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_7_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_8 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_8_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_8_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_8_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_8_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_9 (
    .clka  (clk                             ), //i
    .addra (xil_SimpleDualBram_9_addra[10:0]), //i
    .dina  (sData_payload[63:0]             ), //i
    .ena   (xil_SimpleDualBram_9_ena        ), //i
    .wea   (1'b1                            ), //i
    .addrb (xil_SimpleDualBram_9_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_9_doutb[7:0] ), //o
    .clkb  (clk                             )  //i
  );
  Weight_Bram xil_SimpleDualBram_10 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_10_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_10_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_10_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_10_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_11 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_11_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_11_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_11_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_11_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_12 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_12_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_12_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_12_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_12_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_13 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_13_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_13_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_13_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_13_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_14 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_14_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_14_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_14_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_14_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_15 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_15_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_15_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_15_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_15_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_16 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_16_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_16_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_16_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_16_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_17 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_17_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_17_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_17_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_17_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_18 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_18_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_18_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_18_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_18_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_19 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_19_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_19_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_19_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_19_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_20 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_20_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_20_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_20_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_20_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_21 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_21_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_21_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_21_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_21_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_22 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_22_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_22_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_22_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_22_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_23 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_23_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_23_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_23_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_23_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_24 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_24_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_24_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_24_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_24_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_25 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_25_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_25_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_25_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_25_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_26 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_26_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_26_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_26_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_26_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_27 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_27_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_27_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_27_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_27_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_28 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_28_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_28_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_28_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_28_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_29 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_29_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_29_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_29_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_29_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_30 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_30_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_30_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_30_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_30_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_31 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_31_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_31_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_31_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_31_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_32 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_32_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_32_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_32_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_32_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_33 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_33_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_33_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_33_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_33_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_34 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_34_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_34_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_34_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_34_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_35 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_35_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_35_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_35_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_35_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_36 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_36_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_36_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_36_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_36_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_37 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_37_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_37_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_37_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_37_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_38 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_38_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_38_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_38_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_38_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_39 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_39_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_39_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_39_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_39_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_40 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_40_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_40_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_40_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_40_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_41 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_41_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_41_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_41_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_41_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_42 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_42_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_42_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_42_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_42_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_43 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_43_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_43_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_43_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_43_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_44 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_44_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_44_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_44_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_44_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_45 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_45_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_45_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_45_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_45_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_46 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_46_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_46_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_46_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_46_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_47 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_47_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_47_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_47_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_47_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_48 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_48_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_48_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_48_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_48_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_49 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_49_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_49_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_49_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_49_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_50 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_50_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_50_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_50_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_50_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_51 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_51_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_51_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_51_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_51_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_52 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_52_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_52_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_52_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_52_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_53 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_53_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_53_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_53_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_53_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_54 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_54_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_54_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_54_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_54_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_55 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_55_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_55_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_55_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_55_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_56 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_56_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_56_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_56_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_56_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_57 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_57_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_57_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_57_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_57_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_58 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_58_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_58_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_58_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_58_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_59 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_59_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_59_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_59_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_59_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_60 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_60_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_60_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_60_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_60_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_61 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_61_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_61_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_61_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_61_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_62 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_62_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_62_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_62_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_62_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  Weight_Bram xil_SimpleDualBram_63 (
    .clka  (clk                              ), //i
    .addra (xil_SimpleDualBram_63_addra[10:0]), //i
    .dina  (sData_payload[63:0]              ), //i
    .ena   (xil_SimpleDualBram_63_ena        ), //i
    .wea   (1'b1                             ), //i
    .addrb (xil_SimpleDualBram_63_addrb[13:0]), //i
    .doutb (xil_SimpleDualBram_63_doutb[7:0] ), //o
    .clkb  (clk                              )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      WEIGHT_CACHE_STATUS_IDLE : Fsm_currentState_string = "IDLE        ";
      WEIGHT_CACHE_STATUS_INIT : Fsm_currentState_string = "INIT        ";
      WEIGHT_CACHE_STATUS_CACHE_WEIGHT : Fsm_currentState_string = "CACHE_WEIGHT";
      WEIGHT_CACHE_STATUS_SA_COMPUTE : Fsm_currentState_string = "SA_COMPUTE  ";
      default : Fsm_currentState_string = "????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      WEIGHT_CACHE_STATUS_IDLE : Fsm_nextState_string = "IDLE        ";
      WEIGHT_CACHE_STATUS_INIT : Fsm_nextState_string = "INIT        ";
      WEIGHT_CACHE_STATUS_CACHE_WEIGHT : Fsm_nextState_string = "CACHE_WEIGHT";
      WEIGHT_CACHE_STATUS_SA_COMPUTE : Fsm_nextState_string = "SA_COMPUTE  ";
      default : Fsm_nextState_string = "????????????";
    endcase
  end
  `endif

  assign when_SA3D_WeightCache_l33 = (start && (! start_regNext));
  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & WEIGHT_CACHE_STATUS_IDLE) == WEIGHT_CACHE_STATUS_IDLE) : begin
        if(when_SA3D_WeightCache_l33) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_INIT;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_IDLE;
        end
      end
      (((Fsm_currentState) & WEIGHT_CACHE_STATUS_INIT) == WEIGHT_CACHE_STATUS_INIT) : begin
        if(Fsm_Init_End) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_CACHE_WEIGHT;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_INIT;
        end
      end
      (((Fsm_currentState) & WEIGHT_CACHE_STATUS_CACHE_WEIGHT) == WEIGHT_CACHE_STATUS_CACHE_WEIGHT) : begin
        if(Fsm_Weight_All_Cached) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_SA_COMPUTE;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_CACHE_WEIGHT;
        end
      end
      default : begin
        if(Fsm_SA_Computed) begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_IDLE;
        end else begin
          Fsm_nextState = WEIGHT_CACHE_STATUS_SA_COMPUTE;
        end
      end
    endcase
  end

  assign when_WaCounter_l19 = ((Fsm_currentState & WEIGHT_CACHE_STATUS_INIT) != 4'b0000);
  assign when_WaCounter_l14 = (Init_Count_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l14) begin
      Init_Count_valid = 1'b1;
    end else begin
      Init_Count_valid = 1'b0;
    end
  end

  assign Fsm_Init_End = Init_Count_valid;
  assign Matrix_In_MaxCnt = (Matrix_Row >>> 3);
  assign sData_fire = (sData_valid && sData_ready);
  assign In_Row_Cnt_valid = ((In_Row_Cnt_count == _zz_In_Row_Cnt_valid) && sData_fire);
  assign In_Col_Cnt_valid = ((In_Col_Cnt_count == _zz_In_Col_Cnt_valid) && In_Row_Cnt_valid);
  assign when_WaCounter_l40 = (Raddr_Valid && ((Fsm_currentState & WEIGHT_CACHE_STATUS_SA_COMPUTE) != 4'b0000));
  assign OutRow_Cnt_valid = ((OutRow_Cnt_count == _zz_OutRow_Cnt_valid) && when_WaCounter_l40);
  assign _zz_OutCol_Cnt_count = 7'h40;
  always @(*) begin
    OutCol_Cnt_valid = ((OutCol_Cnt_count <= _zz_OutCol_Cnt_valid) && OutRow_Cnt_valid);
    if(start) begin
      OutCol_Cnt_valid = 1'b0;
    end
  end

  always @(*) begin
    Col_In_8_Cnt_valid = ((Col_In_8_Cnt_count == 6'h3f) && In_Row_Cnt_valid);
    if(OutCol_Cnt_valid) begin
      Col_In_8_Cnt_valid = 1'b0;
    end
  end

  assign when_SA3D_WeightCache_l131 = ((Fsm_currentState & WEIGHT_CACHE_STATUS_INIT) != 4'b0000);
  assign when_SA3D_WeightCache_l136 = ((Fsm_currentState & WEIGHT_CACHE_STATUS_INIT) != 4'b0000);
  assign Fsm_Weight_All_Cached = In_Col_Cnt_valid;
  assign Weight_Cached = In_Col_Cnt_valid;
  assign xil_SimpleDualBram_addra = _zz_addra[10:0];
  assign xil_SimpleDualBram_addrb = _zz_addrb[13:0];
  assign sData_fire_1 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_ena = (_zz_ena[0] && sData_fire_1);
  assign mData_0 = xil_SimpleDualBram_doutb;
  assign xil_SimpleDualBram_1_addra = _zz_addra_1[10:0];
  assign xil_SimpleDualBram_1_addrb = _zz_addrb_1[13:0];
  assign sData_fire_2 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_1_ena = (_zz_ena_1[0] && sData_fire_2);
  assign mData_1 = xil_SimpleDualBram_1_doutb;
  assign xil_SimpleDualBram_2_addra = _zz_addra_2[10:0];
  assign xil_SimpleDualBram_2_addrb = _zz_addrb_2[13:0];
  assign sData_fire_3 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_2_ena = (_zz_ena_2[0] && sData_fire_3);
  assign mData_2 = xil_SimpleDualBram_2_doutb;
  assign xil_SimpleDualBram_3_addra = _zz_addra_3[10:0];
  assign xil_SimpleDualBram_3_addrb = _zz_addrb_3[13:0];
  assign sData_fire_4 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_3_ena = (_zz_ena_3[0] && sData_fire_4);
  assign mData_3 = xil_SimpleDualBram_3_doutb;
  assign xil_SimpleDualBram_4_addra = _zz_addra_4[10:0];
  assign xil_SimpleDualBram_4_addrb = _zz_addrb_4[13:0];
  assign sData_fire_5 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_4_ena = (_zz_ena_4[0] && sData_fire_5);
  assign mData_4 = xil_SimpleDualBram_4_doutb;
  assign xil_SimpleDualBram_5_addra = _zz_addra_5[10:0];
  assign xil_SimpleDualBram_5_addrb = _zz_addrb_5[13:0];
  assign sData_fire_6 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_5_ena = (_zz_ena_5[0] && sData_fire_6);
  assign mData_5 = xil_SimpleDualBram_5_doutb;
  assign xil_SimpleDualBram_6_addra = _zz_addra_6[10:0];
  assign xil_SimpleDualBram_6_addrb = _zz_addrb_6[13:0];
  assign sData_fire_7 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_6_ena = (_zz_ena_6[0] && sData_fire_7);
  assign mData_6 = xil_SimpleDualBram_6_doutb;
  assign xil_SimpleDualBram_7_addra = _zz_addra_7[10:0];
  assign xil_SimpleDualBram_7_addrb = _zz_addrb_7[13:0];
  assign sData_fire_8 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_7_ena = (_zz_ena_7[0] && sData_fire_8);
  assign mData_7 = xil_SimpleDualBram_7_doutb;
  assign xil_SimpleDualBram_8_addra = _zz_addra_8[10:0];
  assign xil_SimpleDualBram_8_addrb = _zz_addrb_8[13:0];
  assign sData_fire_9 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_8_ena = (_zz_ena_8[0] && sData_fire_9);
  assign mData_8 = xil_SimpleDualBram_8_doutb;
  assign xil_SimpleDualBram_9_addra = _zz_addra_9[10:0];
  assign xil_SimpleDualBram_9_addrb = _zz_addrb_9[13:0];
  assign sData_fire_10 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_9_ena = (_zz_ena_9[0] && sData_fire_10);
  assign mData_9 = xil_SimpleDualBram_9_doutb;
  assign xil_SimpleDualBram_10_addra = _zz_addra_10[10:0];
  assign xil_SimpleDualBram_10_addrb = _zz_addrb_10[13:0];
  assign sData_fire_11 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_10_ena = (_zz_ena_10[0] && sData_fire_11);
  assign mData_10 = xil_SimpleDualBram_10_doutb;
  assign xil_SimpleDualBram_11_addra = _zz_addra_11[10:0];
  assign xil_SimpleDualBram_11_addrb = _zz_addrb_11[13:0];
  assign sData_fire_12 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_11_ena = (_zz_ena_11[0] && sData_fire_12);
  assign mData_11 = xil_SimpleDualBram_11_doutb;
  assign xil_SimpleDualBram_12_addra = _zz_addra_12[10:0];
  assign xil_SimpleDualBram_12_addrb = _zz_addrb_12[13:0];
  assign sData_fire_13 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_12_ena = (_zz_ena_12[0] && sData_fire_13);
  assign mData_12 = xil_SimpleDualBram_12_doutb;
  assign xil_SimpleDualBram_13_addra = _zz_addra_13[10:0];
  assign xil_SimpleDualBram_13_addrb = _zz_addrb_13[13:0];
  assign sData_fire_14 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_13_ena = (_zz_ena_13[0] && sData_fire_14);
  assign mData_13 = xil_SimpleDualBram_13_doutb;
  assign xil_SimpleDualBram_14_addra = _zz_addra_14[10:0];
  assign xil_SimpleDualBram_14_addrb = _zz_addrb_14[13:0];
  assign sData_fire_15 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_14_ena = (_zz_ena_14[0] && sData_fire_15);
  assign mData_14 = xil_SimpleDualBram_14_doutb;
  assign xil_SimpleDualBram_15_addra = _zz_addra_15[10:0];
  assign xil_SimpleDualBram_15_addrb = _zz_addrb_15[13:0];
  assign sData_fire_16 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_15_ena = (_zz_ena_15[0] && sData_fire_16);
  assign mData_15 = xil_SimpleDualBram_15_doutb;
  assign xil_SimpleDualBram_16_addra = _zz_addra_16[10:0];
  assign xil_SimpleDualBram_16_addrb = _zz_addrb_16[13:0];
  assign sData_fire_17 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_16_ena = (_zz_ena_16[0] && sData_fire_17);
  assign mData_16 = xil_SimpleDualBram_16_doutb;
  assign xil_SimpleDualBram_17_addra = _zz_addra_17[10:0];
  assign xil_SimpleDualBram_17_addrb = _zz_addrb_17[13:0];
  assign sData_fire_18 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_17_ena = (_zz_ena_17[0] && sData_fire_18);
  assign mData_17 = xil_SimpleDualBram_17_doutb;
  assign xil_SimpleDualBram_18_addra = _zz_addra_18[10:0];
  assign xil_SimpleDualBram_18_addrb = _zz_addrb_18[13:0];
  assign sData_fire_19 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_18_ena = (_zz_ena_18[0] && sData_fire_19);
  assign mData_18 = xil_SimpleDualBram_18_doutb;
  assign xil_SimpleDualBram_19_addra = _zz_addra_19[10:0];
  assign xil_SimpleDualBram_19_addrb = _zz_addrb_19[13:0];
  assign sData_fire_20 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_19_ena = (_zz_ena_19[0] && sData_fire_20);
  assign mData_19 = xil_SimpleDualBram_19_doutb;
  assign xil_SimpleDualBram_20_addra = _zz_addra_20[10:0];
  assign xil_SimpleDualBram_20_addrb = _zz_addrb_20[13:0];
  assign sData_fire_21 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_20_ena = (_zz_ena_20[0] && sData_fire_21);
  assign mData_20 = xil_SimpleDualBram_20_doutb;
  assign xil_SimpleDualBram_21_addra = _zz_addra_21[10:0];
  assign xil_SimpleDualBram_21_addrb = _zz_addrb_21[13:0];
  assign sData_fire_22 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_21_ena = (_zz_ena_21[0] && sData_fire_22);
  assign mData_21 = xil_SimpleDualBram_21_doutb;
  assign xil_SimpleDualBram_22_addra = _zz_addra_22[10:0];
  assign xil_SimpleDualBram_22_addrb = _zz_addrb_22[13:0];
  assign sData_fire_23 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_22_ena = (_zz_ena_22[0] && sData_fire_23);
  assign mData_22 = xil_SimpleDualBram_22_doutb;
  assign xil_SimpleDualBram_23_addra = _zz_addra_23[10:0];
  assign xil_SimpleDualBram_23_addrb = _zz_addrb_23[13:0];
  assign sData_fire_24 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_23_ena = (_zz_ena_23[0] && sData_fire_24);
  assign mData_23 = xil_SimpleDualBram_23_doutb;
  assign xil_SimpleDualBram_24_addra = _zz_addra_24[10:0];
  assign xil_SimpleDualBram_24_addrb = _zz_addrb_24[13:0];
  assign sData_fire_25 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_24_ena = (_zz_ena_24[0] && sData_fire_25);
  assign mData_24 = xil_SimpleDualBram_24_doutb;
  assign xil_SimpleDualBram_25_addra = _zz_addra_25[10:0];
  assign xil_SimpleDualBram_25_addrb = _zz_addrb_25[13:0];
  assign sData_fire_26 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_25_ena = (_zz_ena_25[0] && sData_fire_26);
  assign mData_25 = xil_SimpleDualBram_25_doutb;
  assign xil_SimpleDualBram_26_addra = _zz_addra_26[10:0];
  assign xil_SimpleDualBram_26_addrb = _zz_addrb_26[13:0];
  assign sData_fire_27 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_26_ena = (_zz_ena_26[0] && sData_fire_27);
  assign mData_26 = xil_SimpleDualBram_26_doutb;
  assign xil_SimpleDualBram_27_addra = _zz_addra_27[10:0];
  assign xil_SimpleDualBram_27_addrb = _zz_addrb_27[13:0];
  assign sData_fire_28 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_27_ena = (_zz_ena_27[0] && sData_fire_28);
  assign mData_27 = xil_SimpleDualBram_27_doutb;
  assign xil_SimpleDualBram_28_addra = _zz_addra_28[10:0];
  assign xil_SimpleDualBram_28_addrb = _zz_addrb_28[13:0];
  assign sData_fire_29 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_28_ena = (_zz_ena_28[0] && sData_fire_29);
  assign mData_28 = xil_SimpleDualBram_28_doutb;
  assign xil_SimpleDualBram_29_addra = _zz_addra_29[10:0];
  assign xil_SimpleDualBram_29_addrb = _zz_addrb_29[13:0];
  assign sData_fire_30 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_29_ena = (_zz_ena_29[0] && sData_fire_30);
  assign mData_29 = xil_SimpleDualBram_29_doutb;
  assign xil_SimpleDualBram_30_addra = _zz_addra_30[10:0];
  assign xil_SimpleDualBram_30_addrb = _zz_addrb_30[13:0];
  assign sData_fire_31 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_30_ena = (_zz_ena_30[0] && sData_fire_31);
  assign mData_30 = xil_SimpleDualBram_30_doutb;
  assign xil_SimpleDualBram_31_addra = _zz_addra_31[10:0];
  assign xil_SimpleDualBram_31_addrb = _zz_addrb_31[13:0];
  assign sData_fire_32 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_31_ena = (_zz_ena_31[0] && sData_fire_32);
  assign mData_31 = xil_SimpleDualBram_31_doutb;
  assign xil_SimpleDualBram_32_addra = _zz_addra_32[10:0];
  assign xil_SimpleDualBram_32_addrb = _zz_addrb_32[13:0];
  assign sData_fire_33 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_32_ena = (_zz_ena_32[0] && sData_fire_33);
  assign mData_32 = xil_SimpleDualBram_32_doutb;
  assign xil_SimpleDualBram_33_addra = _zz_addra_33[10:0];
  assign xil_SimpleDualBram_33_addrb = _zz_addrb_33[13:0];
  assign sData_fire_34 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_33_ena = (_zz_ena_33[0] && sData_fire_34);
  assign mData_33 = xil_SimpleDualBram_33_doutb;
  assign xil_SimpleDualBram_34_addra = _zz_addra_34[10:0];
  assign xil_SimpleDualBram_34_addrb = _zz_addrb_34[13:0];
  assign sData_fire_35 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_34_ena = (_zz_ena_34[0] && sData_fire_35);
  assign mData_34 = xil_SimpleDualBram_34_doutb;
  assign xil_SimpleDualBram_35_addra = _zz_addra_35[10:0];
  assign xil_SimpleDualBram_35_addrb = _zz_addrb_35[13:0];
  assign sData_fire_36 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_35_ena = (_zz_ena_35[0] && sData_fire_36);
  assign mData_35 = xil_SimpleDualBram_35_doutb;
  assign xil_SimpleDualBram_36_addra = _zz_addra_36[10:0];
  assign xil_SimpleDualBram_36_addrb = _zz_addrb_36[13:0];
  assign sData_fire_37 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_36_ena = (_zz_ena_36[0] && sData_fire_37);
  assign mData_36 = xil_SimpleDualBram_36_doutb;
  assign xil_SimpleDualBram_37_addra = _zz_addra_37[10:0];
  assign xil_SimpleDualBram_37_addrb = _zz_addrb_37[13:0];
  assign sData_fire_38 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_37_ena = (_zz_ena_37[0] && sData_fire_38);
  assign mData_37 = xil_SimpleDualBram_37_doutb;
  assign xil_SimpleDualBram_38_addra = _zz_addra_38[10:0];
  assign xil_SimpleDualBram_38_addrb = _zz_addrb_38[13:0];
  assign sData_fire_39 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_38_ena = (_zz_ena_38[0] && sData_fire_39);
  assign mData_38 = xil_SimpleDualBram_38_doutb;
  assign xil_SimpleDualBram_39_addra = _zz_addra_39[10:0];
  assign xil_SimpleDualBram_39_addrb = _zz_addrb_39[13:0];
  assign sData_fire_40 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_39_ena = (_zz_ena_39[0] && sData_fire_40);
  assign mData_39 = xil_SimpleDualBram_39_doutb;
  assign xil_SimpleDualBram_40_addra = _zz_addra_40[10:0];
  assign xil_SimpleDualBram_40_addrb = _zz_addrb_40[13:0];
  assign sData_fire_41 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_40_ena = (_zz_ena_40[0] && sData_fire_41);
  assign mData_40 = xil_SimpleDualBram_40_doutb;
  assign xil_SimpleDualBram_41_addra = _zz_addra_41[10:0];
  assign xil_SimpleDualBram_41_addrb = _zz_addrb_41[13:0];
  assign sData_fire_42 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_41_ena = (_zz_ena_41[0] && sData_fire_42);
  assign mData_41 = xil_SimpleDualBram_41_doutb;
  assign xil_SimpleDualBram_42_addra = _zz_addra_42[10:0];
  assign xil_SimpleDualBram_42_addrb = _zz_addrb_42[13:0];
  assign sData_fire_43 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_42_ena = (_zz_ena_42[0] && sData_fire_43);
  assign mData_42 = xil_SimpleDualBram_42_doutb;
  assign xil_SimpleDualBram_43_addra = _zz_addra_43[10:0];
  assign xil_SimpleDualBram_43_addrb = _zz_addrb_43[13:0];
  assign sData_fire_44 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_43_ena = (_zz_ena_43[0] && sData_fire_44);
  assign mData_43 = xil_SimpleDualBram_43_doutb;
  assign xil_SimpleDualBram_44_addra = _zz_addra_44[10:0];
  assign xil_SimpleDualBram_44_addrb = _zz_addrb_44[13:0];
  assign sData_fire_45 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_44_ena = (_zz_ena_44[0] && sData_fire_45);
  assign mData_44 = xil_SimpleDualBram_44_doutb;
  assign xil_SimpleDualBram_45_addra = _zz_addra_45[10:0];
  assign xil_SimpleDualBram_45_addrb = _zz_addrb_45[13:0];
  assign sData_fire_46 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_45_ena = (_zz_ena_45[0] && sData_fire_46);
  assign mData_45 = xil_SimpleDualBram_45_doutb;
  assign xil_SimpleDualBram_46_addra = _zz_addra_46[10:0];
  assign xil_SimpleDualBram_46_addrb = _zz_addrb_46[13:0];
  assign sData_fire_47 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_46_ena = (_zz_ena_46[0] && sData_fire_47);
  assign mData_46 = xil_SimpleDualBram_46_doutb;
  assign xil_SimpleDualBram_47_addra = _zz_addra_47[10:0];
  assign xil_SimpleDualBram_47_addrb = _zz_addrb_47[13:0];
  assign sData_fire_48 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_47_ena = (_zz_ena_47[0] && sData_fire_48);
  assign mData_47 = xil_SimpleDualBram_47_doutb;
  assign xil_SimpleDualBram_48_addra = _zz_addra_48[10:0];
  assign xil_SimpleDualBram_48_addrb = _zz_addrb_48[13:0];
  assign sData_fire_49 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_48_ena = (_zz_ena_48[0] && sData_fire_49);
  assign mData_48 = xil_SimpleDualBram_48_doutb;
  assign xil_SimpleDualBram_49_addra = _zz_addra_49[10:0];
  assign xil_SimpleDualBram_49_addrb = _zz_addrb_49[13:0];
  assign sData_fire_50 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_49_ena = (_zz_ena_49[0] && sData_fire_50);
  assign mData_49 = xil_SimpleDualBram_49_doutb;
  assign xil_SimpleDualBram_50_addra = _zz_addra_50[10:0];
  assign xil_SimpleDualBram_50_addrb = _zz_addrb_50[13:0];
  assign sData_fire_51 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_50_ena = (_zz_ena_50[0] && sData_fire_51);
  assign mData_50 = xil_SimpleDualBram_50_doutb;
  assign xil_SimpleDualBram_51_addra = _zz_addra_51[10:0];
  assign xil_SimpleDualBram_51_addrb = _zz_addrb_51[13:0];
  assign sData_fire_52 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_51_ena = (_zz_ena_51[0] && sData_fire_52);
  assign mData_51 = xil_SimpleDualBram_51_doutb;
  assign xil_SimpleDualBram_52_addra = _zz_addra_52[10:0];
  assign xil_SimpleDualBram_52_addrb = _zz_addrb_52[13:0];
  assign sData_fire_53 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_52_ena = (_zz_ena_52[0] && sData_fire_53);
  assign mData_52 = xil_SimpleDualBram_52_doutb;
  assign xil_SimpleDualBram_53_addra = _zz_addra_53[10:0];
  assign xil_SimpleDualBram_53_addrb = _zz_addrb_53[13:0];
  assign sData_fire_54 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_53_ena = (_zz_ena_53[0] && sData_fire_54);
  assign mData_53 = xil_SimpleDualBram_53_doutb;
  assign xil_SimpleDualBram_54_addra = _zz_addra_54[10:0];
  assign xil_SimpleDualBram_54_addrb = _zz_addrb_54[13:0];
  assign sData_fire_55 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_54_ena = (_zz_ena_54[0] && sData_fire_55);
  assign mData_54 = xil_SimpleDualBram_54_doutb;
  assign xil_SimpleDualBram_55_addra = _zz_addra_55[10:0];
  assign xil_SimpleDualBram_55_addrb = _zz_addrb_55[13:0];
  assign sData_fire_56 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_55_ena = (_zz_ena_55[0] && sData_fire_56);
  assign mData_55 = xil_SimpleDualBram_55_doutb;
  assign xil_SimpleDualBram_56_addra = _zz_addra_56[10:0];
  assign xil_SimpleDualBram_56_addrb = _zz_addrb_56[13:0];
  assign sData_fire_57 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_56_ena = (_zz_ena_56[0] && sData_fire_57);
  assign mData_56 = xil_SimpleDualBram_56_doutb;
  assign xil_SimpleDualBram_57_addra = _zz_addra_57[10:0];
  assign xil_SimpleDualBram_57_addrb = _zz_addrb_57[13:0];
  assign sData_fire_58 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_57_ena = (_zz_ena_57[0] && sData_fire_58);
  assign mData_57 = xil_SimpleDualBram_57_doutb;
  assign xil_SimpleDualBram_58_addra = _zz_addra_58[10:0];
  assign xil_SimpleDualBram_58_addrb = _zz_addrb_58[13:0];
  assign sData_fire_59 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_58_ena = (_zz_ena_58[0] && sData_fire_59);
  assign mData_58 = xil_SimpleDualBram_58_doutb;
  assign xil_SimpleDualBram_59_addra = _zz_addra_59[10:0];
  assign xil_SimpleDualBram_59_addrb = _zz_addrb_59[13:0];
  assign sData_fire_60 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_59_ena = (_zz_ena_59[0] && sData_fire_60);
  assign mData_59 = xil_SimpleDualBram_59_doutb;
  assign xil_SimpleDualBram_60_addra = _zz_addra_60[10:0];
  assign xil_SimpleDualBram_60_addrb = _zz_addrb_60[13:0];
  assign sData_fire_61 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_60_ena = (_zz_ena_60[0] && sData_fire_61);
  assign mData_60 = xil_SimpleDualBram_60_doutb;
  assign xil_SimpleDualBram_61_addra = _zz_addra_61[10:0];
  assign xil_SimpleDualBram_61_addrb = _zz_addrb_61[13:0];
  assign sData_fire_62 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_61_ena = (_zz_ena_61[0] && sData_fire_62);
  assign mData_61 = xil_SimpleDualBram_61_doutb;
  assign xil_SimpleDualBram_62_addra = _zz_addra_62[10:0];
  assign xil_SimpleDualBram_62_addrb = _zz_addrb_62[13:0];
  assign sData_fire_63 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_62_ena = (_zz_ena_62[0] && sData_fire_63);
  assign mData_62 = xil_SimpleDualBram_62_doutb;
  assign xil_SimpleDualBram_63_addra = _zz_addra_63[10:0];
  assign xil_SimpleDualBram_63_addrb = _zz_addrb_63[13:0];
  assign sData_fire_64 = (sData_valid && sData_ready);
  assign xil_SimpleDualBram_63_ena = (_zz_ena_63[0] && sData_fire_64);
  assign mData_63 = xil_SimpleDualBram_63_doutb;
  assign sData_ready = ((Fsm_currentState & WEIGHT_CACHE_STATUS_CACHE_WEIGHT) != 4'b0000);
  assign Fsm_SA_Computed = LayerEnd;
  always @(*) begin
    case(OutCol_Cnt_count)
      16'h0001 : begin
        MatrixCol_Switch_1[0 : 0] = 1'b1;
        MatrixCol_Switch_1[63 : 1] = 63'h0;
      end
      16'h0002 : begin
        MatrixCol_Switch_1[1 : 0] = 2'b11;
        MatrixCol_Switch_1[63 : 2] = 62'h0;
      end
      16'h0003 : begin
        MatrixCol_Switch_1[2 : 0] = 3'b111;
        MatrixCol_Switch_1[63 : 3] = 61'h0;
      end
      16'h0004 : begin
        MatrixCol_Switch_1[3 : 0] = 4'b1111;
        MatrixCol_Switch_1[63 : 4] = 60'h0;
      end
      16'h0005 : begin
        MatrixCol_Switch_1[4 : 0] = 5'h1f;
        MatrixCol_Switch_1[63 : 5] = 59'h0;
      end
      16'h0006 : begin
        MatrixCol_Switch_1[5 : 0] = 6'h3f;
        MatrixCol_Switch_1[63 : 6] = 58'h0;
      end
      16'h0007 : begin
        MatrixCol_Switch_1[6 : 0] = 7'h7f;
        MatrixCol_Switch_1[63 : 7] = 57'h0;
      end
      16'h0008 : begin
        MatrixCol_Switch_1[7 : 0] = 8'hff;
        MatrixCol_Switch_1[63 : 8] = 56'h0;
      end
      16'h0009 : begin
        MatrixCol_Switch_1[8 : 0] = 9'h1ff;
        MatrixCol_Switch_1[63 : 9] = 55'h0;
      end
      16'h000a : begin
        MatrixCol_Switch_1[9 : 0] = 10'h3ff;
        MatrixCol_Switch_1[63 : 10] = 54'h0;
      end
      16'h000b : begin
        MatrixCol_Switch_1[10 : 0] = 11'h7ff;
        MatrixCol_Switch_1[63 : 11] = 53'h0;
      end
      16'h000c : begin
        MatrixCol_Switch_1[11 : 0] = 12'hfff;
        MatrixCol_Switch_1[63 : 12] = 52'h0;
      end
      16'h000d : begin
        MatrixCol_Switch_1[12 : 0] = 13'h1fff;
        MatrixCol_Switch_1[63 : 13] = 51'h0;
      end
      16'h000e : begin
        MatrixCol_Switch_1[13 : 0] = 14'h3fff;
        MatrixCol_Switch_1[63 : 14] = 50'h0;
      end
      16'h000f : begin
        MatrixCol_Switch_1[14 : 0] = 15'h7fff;
        MatrixCol_Switch_1[63 : 15] = 49'h0;
      end
      16'h0010 : begin
        MatrixCol_Switch_1[15 : 0] = 16'hffff;
        MatrixCol_Switch_1[63 : 16] = 48'h0;
      end
      16'h0011 : begin
        MatrixCol_Switch_1[16 : 0] = 17'h1ffff;
        MatrixCol_Switch_1[63 : 17] = 47'h0;
      end
      16'h0012 : begin
        MatrixCol_Switch_1[17 : 0] = 18'h3ffff;
        MatrixCol_Switch_1[63 : 18] = 46'h0;
      end
      16'h0013 : begin
        MatrixCol_Switch_1[18 : 0] = 19'h7ffff;
        MatrixCol_Switch_1[63 : 19] = 45'h0;
      end
      16'h0014 : begin
        MatrixCol_Switch_1[19 : 0] = 20'hfffff;
        MatrixCol_Switch_1[63 : 20] = 44'h0;
      end
      16'h0015 : begin
        MatrixCol_Switch_1[20 : 0] = 21'h1fffff;
        MatrixCol_Switch_1[63 : 21] = 43'h0;
      end
      16'h0016 : begin
        MatrixCol_Switch_1[21 : 0] = 22'h3fffff;
        MatrixCol_Switch_1[63 : 22] = 42'h0;
      end
      16'h0017 : begin
        MatrixCol_Switch_1[22 : 0] = 23'h7fffff;
        MatrixCol_Switch_1[63 : 23] = 41'h0;
      end
      16'h0018 : begin
        MatrixCol_Switch_1[23 : 0] = 24'hffffff;
        MatrixCol_Switch_1[63 : 24] = 40'h0;
      end
      16'h0019 : begin
        MatrixCol_Switch_1[24 : 0] = 25'h1ffffff;
        MatrixCol_Switch_1[63 : 25] = 39'h0;
      end
      16'h001a : begin
        MatrixCol_Switch_1[25 : 0] = 26'h3ffffff;
        MatrixCol_Switch_1[63 : 26] = 38'h0;
      end
      16'h001b : begin
        MatrixCol_Switch_1[26 : 0] = 27'h7ffffff;
        MatrixCol_Switch_1[63 : 27] = 37'h0;
      end
      16'h001c : begin
        MatrixCol_Switch_1[27 : 0] = 28'hfffffff;
        MatrixCol_Switch_1[63 : 28] = 36'h0;
      end
      16'h001d : begin
        MatrixCol_Switch_1[28 : 0] = 29'h1fffffff;
        MatrixCol_Switch_1[63 : 29] = 35'h0;
      end
      16'h001e : begin
        MatrixCol_Switch_1[29 : 0] = 30'h3fffffff;
        MatrixCol_Switch_1[63 : 30] = 34'h0;
      end
      16'h001f : begin
        MatrixCol_Switch_1[30 : 0] = 31'h7fffffff;
        MatrixCol_Switch_1[63 : 31] = 33'h0;
      end
      16'h0020 : begin
        MatrixCol_Switch_1[31 : 0] = 32'hffffffff;
        MatrixCol_Switch_1[63 : 32] = 32'h0;
      end
      16'h0021 : begin
        MatrixCol_Switch_1[32 : 0] = 33'h1ffffffff;
        MatrixCol_Switch_1[63 : 33] = 31'h0;
      end
      16'h0022 : begin
        MatrixCol_Switch_1[33 : 0] = 34'h3ffffffff;
        MatrixCol_Switch_1[63 : 34] = 30'h0;
      end
      16'h0023 : begin
        MatrixCol_Switch_1[34 : 0] = 35'h7ffffffff;
        MatrixCol_Switch_1[63 : 35] = 29'h0;
      end
      16'h0024 : begin
        MatrixCol_Switch_1[35 : 0] = 36'hfffffffff;
        MatrixCol_Switch_1[63 : 36] = 28'h0;
      end
      16'h0025 : begin
        MatrixCol_Switch_1[36 : 0] = 37'h1fffffffff;
        MatrixCol_Switch_1[63 : 37] = 27'h0;
      end
      16'h0026 : begin
        MatrixCol_Switch_1[37 : 0] = 38'h3fffffffff;
        MatrixCol_Switch_1[63 : 38] = 26'h0;
      end
      16'h0027 : begin
        MatrixCol_Switch_1[38 : 0] = 39'h7fffffffff;
        MatrixCol_Switch_1[63 : 39] = 25'h0;
      end
      16'h0028 : begin
        MatrixCol_Switch_1[39 : 0] = 40'hffffffffff;
        MatrixCol_Switch_1[63 : 40] = 24'h0;
      end
      16'h0029 : begin
        MatrixCol_Switch_1[40 : 0] = 41'h1ffffffffff;
        MatrixCol_Switch_1[63 : 41] = 23'h0;
      end
      16'h002a : begin
        MatrixCol_Switch_1[41 : 0] = 42'h3ffffffffff;
        MatrixCol_Switch_1[63 : 42] = 22'h0;
      end
      16'h002b : begin
        MatrixCol_Switch_1[42 : 0] = 43'h7ffffffffff;
        MatrixCol_Switch_1[63 : 43] = 21'h0;
      end
      16'h002c : begin
        MatrixCol_Switch_1[43 : 0] = 44'hfffffffffff;
        MatrixCol_Switch_1[63 : 44] = 20'h0;
      end
      16'h002d : begin
        MatrixCol_Switch_1[44 : 0] = 45'h1fffffffffff;
        MatrixCol_Switch_1[63 : 45] = 19'h0;
      end
      16'h002e : begin
        MatrixCol_Switch_1[45 : 0] = 46'h3fffffffffff;
        MatrixCol_Switch_1[63 : 46] = 18'h0;
      end
      16'h002f : begin
        MatrixCol_Switch_1[46 : 0] = 47'h7fffffffffff;
        MatrixCol_Switch_1[63 : 47] = 17'h0;
      end
      16'h0030 : begin
        MatrixCol_Switch_1[47 : 0] = 48'hffffffffffff;
        MatrixCol_Switch_1[63 : 48] = 16'h0;
      end
      16'h0031 : begin
        MatrixCol_Switch_1[48 : 0] = 49'h1ffffffffffff;
        MatrixCol_Switch_1[63 : 49] = 15'h0;
      end
      16'h0032 : begin
        MatrixCol_Switch_1[49 : 0] = 50'h3ffffffffffff;
        MatrixCol_Switch_1[63 : 50] = 14'h0;
      end
      16'h0033 : begin
        MatrixCol_Switch_1[50 : 0] = 51'h7ffffffffffff;
        MatrixCol_Switch_1[63 : 51] = 13'h0;
      end
      16'h0034 : begin
        MatrixCol_Switch_1[51 : 0] = 52'hfffffffffffff;
        MatrixCol_Switch_1[63 : 52] = 12'h0;
      end
      16'h0035 : begin
        MatrixCol_Switch_1[52 : 0] = 53'h1fffffffffffff;
        MatrixCol_Switch_1[63 : 53] = 11'h0;
      end
      16'h0036 : begin
        MatrixCol_Switch_1[53 : 0] = 54'h3fffffffffffff;
        MatrixCol_Switch_1[63 : 54] = 10'h0;
      end
      16'h0037 : begin
        MatrixCol_Switch_1[54 : 0] = 55'h7fffffffffffff;
        MatrixCol_Switch_1[63 : 55] = 9'h0;
      end
      16'h0038 : begin
        MatrixCol_Switch_1[55 : 0] = 56'hffffffffffffff;
        MatrixCol_Switch_1[63 : 56] = 8'h0;
      end
      16'h0039 : begin
        MatrixCol_Switch_1[56 : 0] = 57'h1ffffffffffffff;
        MatrixCol_Switch_1[63 : 57] = 7'h0;
      end
      16'h003a : begin
        MatrixCol_Switch_1[57 : 0] = 58'h3ffffffffffffff;
        MatrixCol_Switch_1[63 : 58] = 6'h0;
      end
      16'h003b : begin
        MatrixCol_Switch_1[58 : 0] = 59'h7ffffffffffffff;
        MatrixCol_Switch_1[63 : 59] = 5'h0;
      end
      16'h003c : begin
        MatrixCol_Switch_1[59 : 0] = 60'hfffffffffffffff;
        MatrixCol_Switch_1[63 : 60] = 4'b0000;
      end
      16'h003d : begin
        MatrixCol_Switch_1[60 : 0] = 61'h1fffffffffffffff;
        MatrixCol_Switch_1[63 : 61] = 3'b000;
      end
      16'h003e : begin
        MatrixCol_Switch_1[61 : 0] = 62'h3fffffffffffffff;
        MatrixCol_Switch_1[63 : 62] = 2'b00;
      end
      16'h003f : begin
        MatrixCol_Switch_1[62 : 0] = 63'h7fffffffffffffff;
        MatrixCol_Switch_1[63 : 63] = 1'b0;
      end
      default : begin
        MatrixCol_Switch_1 = 64'hffffffffffffffff;
      end
    endcase
  end

  assign MatrixCol_Switch = MatrixCol_Switch_1_regNext;
  always @(posedge clk) begin
    start_regNext <= start;
    if(OutRow_Cnt_valid) begin
      if(OutCol_Cnt_valid) begin
        OutCol_Cnt_count <= Matrix_Col;
      end else begin
        OutCol_Cnt_count <= (OutCol_Cnt_count - _zz_OutCol_Cnt_count_1);
      end
    end
    if(start) begin
      OutCol_Cnt_count <= Matrix_Col;
    end
    MatrixCol_Switch_1_regNext <= MatrixCol_Switch_1;
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= WEIGHT_CACHE_STATUS_IDLE;
      Init_Count_count <= 3'b000;
      InData_Switch <= 64'h0000000000000001;
      In_Row_Cnt_count <= 16'h0;
      In_Col_Cnt_count <= 16'h0;
      Read_Row_Base_Addr <= 16'h0;
      Write_Row_Base_Addr <= 16'h0;
      OutRow_Cnt_count <= 16'h0;
      Col_In_8_Cnt_count <= 6'h0;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l19) begin
        Init_Count_count <= (Init_Count_count + 3'b001);
        if(Init_Count_valid) begin
          Init_Count_count <= 3'b000;
        end
      end
      if(sData_fire) begin
        if(In_Row_Cnt_valid) begin
          In_Row_Cnt_count <= 16'h0;
        end else begin
          In_Row_Cnt_count <= (In_Row_Cnt_count + 16'h0001);
        end
      end
      if(In_Row_Cnt_valid) begin
        if(In_Col_Cnt_valid) begin
          In_Col_Cnt_count <= 16'h0;
        end else begin
          In_Col_Cnt_count <= (In_Col_Cnt_count + 16'h0001);
        end
      end
      if(when_WaCounter_l40) begin
        if(OutRow_Cnt_valid) begin
          OutRow_Cnt_count <= 16'h0;
        end else begin
          OutRow_Cnt_count <= (OutRow_Cnt_count + 16'h0001);
        end
      end
      if(In_Row_Cnt_valid) begin
        if(Col_In_8_Cnt_valid) begin
          Col_In_8_Cnt_count <= 6'h0;
        end else begin
          Col_In_8_Cnt_count <= (Col_In_8_Cnt_count + 6'h01);
        end
      end
      if(OutCol_Cnt_valid) begin
        Col_In_8_Cnt_count <= 6'h0;
        Read_Row_Base_Addr <= 16'h0;
      end else begin
        if(OutRow_Cnt_valid) begin
          Read_Row_Base_Addr <= (Read_Row_Base_Addr + Matrix_Row);
        end
      end
      if(when_SA3D_WeightCache_l131) begin
        InData_Switch <= 64'h0000000000000001;
      end else begin
        if(In_Row_Cnt_valid) begin
          InData_Switch <= {InData_Switch[62 : 0],InData_Switch[63 : 63]};
        end
      end
      if(when_SA3D_WeightCache_l136) begin
        Write_Row_Base_Addr <= 16'h0;
      end else begin
        if(Col_In_8_Cnt_valid) begin
          Write_Row_Base_Addr <= (Write_Row_Base_Addr + _zz_Write_Row_Base_Addr);
        end
      end
    end
  end


endmodule

module SA_2D (
  input      [7:0]    io_MatrixA_0,
  input      [7:0]    io_MatrixA_1,
  input      [7:0]    io_MatrixA_2,
  input      [7:0]    io_MatrixA_3,
  input      [7:0]    io_MatrixA_4,
  input      [7:0]    io_MatrixA_5,
  input      [7:0]    io_MatrixA_6,
  input      [7:0]    io_MatrixA_7,
  input      [7:0]    io_MatrixB_0,
  input      [7:0]    io_MatrixB_1,
  input      [7:0]    io_MatrixB_2,
  input      [7:0]    io_MatrixB_3,
  input      [7:0]    io_MatrixB_4,
  input      [7:0]    io_MatrixB_5,
  input      [7:0]    io_MatrixB_6,
  input      [7:0]    io_MatrixB_7,
  input      [7:0]    io_MatrixB_8,
  input      [7:0]    io_MatrixB_9,
  input      [7:0]    io_MatrixB_10,
  input      [7:0]    io_MatrixB_11,
  input      [7:0]    io_MatrixB_12,
  input      [7:0]    io_MatrixB_13,
  input      [7:0]    io_MatrixB_14,
  input      [7:0]    io_MatrixB_15,
  input      [7:0]    io_MatrixB_16,
  input      [7:0]    io_MatrixB_17,
  input      [7:0]    io_MatrixB_18,
  input      [7:0]    io_MatrixB_19,
  input      [7:0]    io_MatrixB_20,
  input      [7:0]    io_MatrixB_21,
  input      [7:0]    io_MatrixB_22,
  input      [7:0]    io_MatrixB_23,
  input      [7:0]    io_MatrixB_24,
  input      [7:0]    io_MatrixB_25,
  input      [7:0]    io_MatrixB_26,
  input      [7:0]    io_MatrixB_27,
  input      [7:0]    io_MatrixB_28,
  input      [7:0]    io_MatrixB_29,
  input      [7:0]    io_MatrixB_30,
  input      [7:0]    io_MatrixB_31,
  input      [7:0]    io_MatrixB_32,
  input      [7:0]    io_MatrixB_33,
  input      [7:0]    io_MatrixB_34,
  input      [7:0]    io_MatrixB_35,
  input      [7:0]    io_MatrixB_36,
  input      [7:0]    io_MatrixB_37,
  input      [7:0]    io_MatrixB_38,
  input      [7:0]    io_MatrixB_39,
  input      [7:0]    io_MatrixB_40,
  input      [7:0]    io_MatrixB_41,
  input      [7:0]    io_MatrixB_42,
  input      [7:0]    io_MatrixB_43,
  input      [7:0]    io_MatrixB_44,
  input      [7:0]    io_MatrixB_45,
  input      [7:0]    io_MatrixB_46,
  input      [7:0]    io_MatrixB_47,
  input      [7:0]    io_MatrixB_48,
  input      [7:0]    io_MatrixB_49,
  input      [7:0]    io_MatrixB_50,
  input      [7:0]    io_MatrixB_51,
  input      [7:0]    io_MatrixB_52,
  input      [7:0]    io_MatrixB_53,
  input      [7:0]    io_MatrixB_54,
  input      [7:0]    io_MatrixB_55,
  input      [7:0]    io_MatrixB_56,
  input      [7:0]    io_MatrixB_57,
  input      [7:0]    io_MatrixB_58,
  input      [7:0]    io_MatrixB_59,
  input      [7:0]    io_MatrixB_60,
  input      [7:0]    io_MatrixB_61,
  input      [7:0]    io_MatrixB_62,
  input      [7:0]    io_MatrixB_63,
  input               io_A_Valid_0,
  input               io_A_Valid_1,
  input               io_A_Valid_2,
  input               io_A_Valid_3,
  input               io_A_Valid_4,
  input               io_A_Valid_5,
  input               io_A_Valid_6,
  input               io_A_Valid_7,
  input               io_B_Valid_0,
  input               io_B_Valid_1,
  input               io_B_Valid_2,
  input               io_B_Valid_3,
  input               io_B_Valid_4,
  input               io_B_Valid_5,
  input               io_B_Valid_6,
  input               io_B_Valid_7,
  input               io_B_Valid_8,
  input               io_B_Valid_9,
  input               io_B_Valid_10,
  input               io_B_Valid_11,
  input               io_B_Valid_12,
  input               io_B_Valid_13,
  input               io_B_Valid_14,
  input               io_B_Valid_15,
  input               io_B_Valid_16,
  input               io_B_Valid_17,
  input               io_B_Valid_18,
  input               io_B_Valid_19,
  input               io_B_Valid_20,
  input               io_B_Valid_21,
  input               io_B_Valid_22,
  input               io_B_Valid_23,
  input               io_B_Valid_24,
  input               io_B_Valid_25,
  input               io_B_Valid_26,
  input               io_B_Valid_27,
  input               io_B_Valid_28,
  input               io_B_Valid_29,
  input               io_B_Valid_30,
  input               io_B_Valid_31,
  input               io_B_Valid_32,
  input               io_B_Valid_33,
  input               io_B_Valid_34,
  input               io_B_Valid_35,
  input               io_B_Valid_36,
  input               io_B_Valid_37,
  input               io_B_Valid_38,
  input               io_B_Valid_39,
  input               io_B_Valid_40,
  input               io_B_Valid_41,
  input               io_B_Valid_42,
  input               io_B_Valid_43,
  input               io_B_Valid_44,
  input               io_B_Valid_45,
  input               io_B_Valid_46,
  input               io_B_Valid_47,
  input               io_B_Valid_48,
  input               io_B_Valid_49,
  input               io_B_Valid_50,
  input               io_B_Valid_51,
  input               io_B_Valid_52,
  input               io_B_Valid_53,
  input               io_B_Valid_54,
  input               io_B_Valid_55,
  input               io_B_Valid_56,
  input               io_B_Valid_57,
  input               io_B_Valid_58,
  input               io_B_Valid_59,
  input               io_B_Valid_60,
  input               io_B_Valid_61,
  input               io_B_Valid_62,
  input               io_B_Valid_63,
  input      [15:0]   io_signCount,
  output reg [31:0]   MatrixC_0,
  output reg [31:0]   MatrixC_1,
  output reg [31:0]   MatrixC_2,
  output reg [31:0]   MatrixC_3,
  output reg [31:0]   MatrixC_4,
  output reg [31:0]   MatrixC_5,
  output reg [31:0]   MatrixC_6,
  output reg [31:0]   MatrixC_7,
  output              C_Valid_0,
  output              C_Valid_1,
  output              C_Valid_2,
  output              C_Valid_3,
  output              C_Valid_4,
  output              C_Valid_5,
  output              C_Valid_6,
  output              C_Valid_7,
  input               start,
  input               clk,
  input               reset
);

  wire                PE00_valid;
  wire                PE01_valid;
  wire                PE02_valid;
  wire                PE03_valid;
  wire                PE04_valid;
  wire                PE05_valid;
  wire                PE06_valid;
  wire                PE07_valid;
  wire                PE08_valid;
  wire                PE09_valid;
  wire                PE010_valid;
  wire                PE011_valid;
  wire                PE012_valid;
  wire                PE013_valid;
  wire                PE014_valid;
  wire                PE015_valid;
  wire                PE016_valid;
  wire                PE017_valid;
  wire                PE018_valid;
  wire                PE019_valid;
  wire                PE020_valid;
  wire                PE021_valid;
  wire                PE022_valid;
  wire                PE023_valid;
  wire                PE024_valid;
  wire                PE025_valid;
  wire                PE026_valid;
  wire                PE027_valid;
  wire                PE028_valid;
  wire                PE029_valid;
  wire                PE030_valid;
  wire                PE031_valid;
  wire                PE032_valid;
  wire                PE033_valid;
  wire                PE034_valid;
  wire                PE035_valid;
  wire                PE036_valid;
  wire                PE037_valid;
  wire                PE038_valid;
  wire                PE039_valid;
  wire                PE040_valid;
  wire                PE041_valid;
  wire                PE042_valid;
  wire                PE043_valid;
  wire                PE044_valid;
  wire                PE045_valid;
  wire                PE046_valid;
  wire                PE047_valid;
  wire                PE048_valid;
  wire                PE049_valid;
  wire                PE050_valid;
  wire                PE051_valid;
  wire                PE052_valid;
  wire                PE053_valid;
  wire                PE054_valid;
  wire                PE055_valid;
  wire                PE056_valid;
  wire                PE057_valid;
  wire                PE058_valid;
  wire                PE059_valid;
  wire                PE060_valid;
  wire                PE061_valid;
  wire                PE062_valid;
  wire                PE063_valid;
  wire                PE10_valid;
  wire                PE11_valid;
  wire                PE12_valid;
  wire                PE13_valid;
  wire                PE14_valid;
  wire                PE15_valid;
  wire                PE16_valid;
  wire                PE17_valid;
  wire                PE18_valid;
  wire                PE19_valid;
  wire                PE110_valid;
  wire                PE111_valid;
  wire                PE112_valid;
  wire                PE113_valid;
  wire                PE114_valid;
  wire                PE115_valid;
  wire                PE116_valid;
  wire                PE117_valid;
  wire                PE118_valid;
  wire                PE119_valid;
  wire                PE120_valid;
  wire                PE121_valid;
  wire                PE122_valid;
  wire                PE123_valid;
  wire                PE124_valid;
  wire                PE125_valid;
  wire                PE126_valid;
  wire                PE127_valid;
  wire                PE128_valid;
  wire                PE129_valid;
  wire                PE130_valid;
  wire                PE131_valid;
  wire                PE132_valid;
  wire                PE133_valid;
  wire                PE134_valid;
  wire                PE135_valid;
  wire                PE136_valid;
  wire                PE137_valid;
  wire                PE138_valid;
  wire                PE139_valid;
  wire                PE140_valid;
  wire                PE141_valid;
  wire                PE142_valid;
  wire                PE143_valid;
  wire                PE144_valid;
  wire                PE145_valid;
  wire                PE146_valid;
  wire                PE147_valid;
  wire                PE148_valid;
  wire                PE149_valid;
  wire                PE150_valid;
  wire                PE151_valid;
  wire                PE152_valid;
  wire                PE153_valid;
  wire                PE154_valid;
  wire                PE155_valid;
  wire                PE156_valid;
  wire                PE157_valid;
  wire                PE158_valid;
  wire                PE159_valid;
  wire                PE160_valid;
  wire                PE161_valid;
  wire                PE162_valid;
  wire                PE163_valid;
  wire                PE20_valid;
  wire                PE21_valid;
  wire                PE22_valid;
  wire                PE23_valid;
  wire                PE24_valid;
  wire                PE25_valid;
  wire                PE26_valid;
  wire                PE27_valid;
  wire                PE28_valid;
  wire                PE29_valid;
  wire                PE210_valid;
  wire                PE211_valid;
  wire                PE212_valid;
  wire                PE213_valid;
  wire                PE214_valid;
  wire                PE215_valid;
  wire                PE216_valid;
  wire                PE217_valid;
  wire                PE218_valid;
  wire                PE219_valid;
  wire                PE220_valid;
  wire                PE221_valid;
  wire                PE222_valid;
  wire                PE223_valid;
  wire                PE224_valid;
  wire                PE225_valid;
  wire                PE226_valid;
  wire                PE227_valid;
  wire                PE228_valid;
  wire                PE229_valid;
  wire                PE230_valid;
  wire                PE231_valid;
  wire                PE232_valid;
  wire                PE233_valid;
  wire                PE234_valid;
  wire                PE235_valid;
  wire                PE236_valid;
  wire                PE237_valid;
  wire                PE238_valid;
  wire                PE239_valid;
  wire                PE240_valid;
  wire                PE241_valid;
  wire                PE242_valid;
  wire                PE243_valid;
  wire                PE244_valid;
  wire                PE245_valid;
  wire                PE246_valid;
  wire                PE247_valid;
  wire                PE248_valid;
  wire                PE249_valid;
  wire                PE250_valid;
  wire                PE251_valid;
  wire                PE252_valid;
  wire                PE253_valid;
  wire                PE254_valid;
  wire                PE255_valid;
  wire                PE256_valid;
  wire                PE257_valid;
  wire                PE258_valid;
  wire                PE259_valid;
  wire                PE260_valid;
  wire                PE261_valid;
  wire                PE262_valid;
  wire                PE263_valid;
  wire                PE30_valid;
  wire                PE31_valid;
  wire                PE32_valid;
  wire                PE33_valid;
  wire                PE34_valid;
  wire                PE35_valid;
  wire                PE36_valid;
  wire                PE37_valid;
  wire                PE38_valid;
  wire                PE39_valid;
  wire                PE310_valid;
  wire                PE311_valid;
  wire                PE312_valid;
  wire                PE313_valid;
  wire                PE314_valid;
  wire                PE315_valid;
  wire                PE316_valid;
  wire                PE317_valid;
  wire                PE318_valid;
  wire                PE319_valid;
  wire                PE320_valid;
  wire                PE321_valid;
  wire                PE322_valid;
  wire                PE323_valid;
  wire                PE324_valid;
  wire                PE325_valid;
  wire                PE326_valid;
  wire                PE327_valid;
  wire                PE328_valid;
  wire                PE329_valid;
  wire                PE330_valid;
  wire                PE331_valid;
  wire                PE332_valid;
  wire                PE333_valid;
  wire                PE334_valid;
  wire                PE335_valid;
  wire                PE336_valid;
  wire                PE337_valid;
  wire                PE338_valid;
  wire                PE339_valid;
  wire                PE340_valid;
  wire                PE341_valid;
  wire                PE342_valid;
  wire                PE343_valid;
  wire                PE344_valid;
  wire                PE345_valid;
  wire                PE346_valid;
  wire                PE347_valid;
  wire                PE348_valid;
  wire                PE349_valid;
  wire                PE350_valid;
  wire                PE351_valid;
  wire                PE352_valid;
  wire                PE353_valid;
  wire                PE354_valid;
  wire                PE355_valid;
  wire                PE356_valid;
  wire                PE357_valid;
  wire                PE358_valid;
  wire                PE359_valid;
  wire                PE360_valid;
  wire                PE361_valid;
  wire                PE362_valid;
  wire                PE363_valid;
  wire                PE40_valid;
  wire                PE41_valid;
  wire                PE42_valid;
  wire                PE43_valid;
  wire                PE44_valid;
  wire                PE45_valid;
  wire                PE46_valid;
  wire                PE47_valid;
  wire                PE48_valid;
  wire                PE49_valid;
  wire                PE410_valid;
  wire                PE411_valid;
  wire                PE412_valid;
  wire                PE413_valid;
  wire                PE414_valid;
  wire                PE415_valid;
  wire                PE416_valid;
  wire                PE417_valid;
  wire                PE418_valid;
  wire                PE419_valid;
  wire                PE420_valid;
  wire                PE421_valid;
  wire                PE422_valid;
  wire                PE423_valid;
  wire                PE424_valid;
  wire                PE425_valid;
  wire                PE426_valid;
  wire                PE427_valid;
  wire                PE428_valid;
  wire                PE429_valid;
  wire                PE430_valid;
  wire                PE431_valid;
  wire                PE432_valid;
  wire                PE433_valid;
  wire                PE434_valid;
  wire                PE435_valid;
  wire                PE436_valid;
  wire                PE437_valid;
  wire                PE438_valid;
  wire                PE439_valid;
  wire                PE440_valid;
  wire                PE441_valid;
  wire                PE442_valid;
  wire                PE443_valid;
  wire                PE444_valid;
  wire                PE445_valid;
  wire                PE446_valid;
  wire                PE447_valid;
  wire                PE448_valid;
  wire                PE449_valid;
  wire                PE450_valid;
  wire                PE451_valid;
  wire                PE452_valid;
  wire                PE453_valid;
  wire                PE454_valid;
  wire                PE455_valid;
  wire                PE456_valid;
  wire                PE457_valid;
  wire                PE458_valid;
  wire                PE459_valid;
  wire                PE460_valid;
  wire                PE461_valid;
  wire                PE462_valid;
  wire                PE463_valid;
  wire                PE50_valid;
  wire                PE51_valid;
  wire                PE52_valid;
  wire                PE53_valid;
  wire                PE54_valid;
  wire                PE55_valid;
  wire                PE56_valid;
  wire                PE57_valid;
  wire                PE58_valid;
  wire                PE59_valid;
  wire                PE510_valid;
  wire                PE511_valid;
  wire                PE512_valid;
  wire                PE513_valid;
  wire                PE514_valid;
  wire                PE515_valid;
  wire                PE516_valid;
  wire                PE517_valid;
  wire                PE518_valid;
  wire                PE519_valid;
  wire                PE520_valid;
  wire                PE521_valid;
  wire                PE522_valid;
  wire                PE523_valid;
  wire                PE524_valid;
  wire                PE525_valid;
  wire                PE526_valid;
  wire                PE527_valid;
  wire                PE528_valid;
  wire                PE529_valid;
  wire                PE530_valid;
  wire                PE531_valid;
  wire                PE532_valid;
  wire                PE533_valid;
  wire                PE534_valid;
  wire                PE535_valid;
  wire                PE536_valid;
  wire                PE537_valid;
  wire                PE538_valid;
  wire                PE539_valid;
  wire                PE540_valid;
  wire                PE541_valid;
  wire                PE542_valid;
  wire                PE543_valid;
  wire                PE544_valid;
  wire                PE545_valid;
  wire                PE546_valid;
  wire                PE547_valid;
  wire                PE548_valid;
  wire                PE549_valid;
  wire                PE550_valid;
  wire                PE551_valid;
  wire                PE552_valid;
  wire                PE553_valid;
  wire                PE554_valid;
  wire                PE555_valid;
  wire                PE556_valid;
  wire                PE557_valid;
  wire                PE558_valid;
  wire                PE559_valid;
  wire                PE560_valid;
  wire                PE561_valid;
  wire                PE562_valid;
  wire                PE563_valid;
  wire                PE60_valid;
  wire                PE61_valid;
  wire                PE62_valid;
  wire                PE63_valid;
  wire                PE64_valid;
  wire                PE65_valid;
  wire                PE66_valid;
  wire                PE67_valid;
  wire                PE68_valid;
  wire                PE69_valid;
  wire                PE610_valid;
  wire                PE611_valid;
  wire                PE612_valid;
  wire                PE613_valid;
  wire                PE614_valid;
  wire                PE615_valid;
  wire                PE616_valid;
  wire                PE617_valid;
  wire                PE618_valid;
  wire                PE619_valid;
  wire                PE620_valid;
  wire                PE621_valid;
  wire                PE622_valid;
  wire                PE623_valid;
  wire                PE624_valid;
  wire                PE625_valid;
  wire                PE626_valid;
  wire                PE627_valid;
  wire                PE628_valid;
  wire                PE629_valid;
  wire                PE630_valid;
  wire                PE631_valid;
  wire                PE632_valid;
  wire                PE633_valid;
  wire                PE634_valid;
  wire                PE635_valid;
  wire                PE636_valid;
  wire                PE637_valid;
  wire                PE638_valid;
  wire                PE639_valid;
  wire                PE640_valid;
  wire                PE641_valid;
  wire                PE642_valid;
  wire                PE643_valid;
  wire                PE644_valid;
  wire                PE645_valid;
  wire                PE646_valid;
  wire                PE647_valid;
  wire                PE648_valid;
  wire                PE649_valid;
  wire                PE650_valid;
  wire                PE651_valid;
  wire                PE652_valid;
  wire                PE653_valid;
  wire                PE654_valid;
  wire                PE655_valid;
  wire                PE656_valid;
  wire                PE657_valid;
  wire                PE658_valid;
  wire                PE659_valid;
  wire                PE660_valid;
  wire                PE661_valid;
  wire                PE662_valid;
  wire                PE663_valid;
  wire                PE70_valid;
  wire                PE71_valid;
  wire                PE72_valid;
  wire                PE73_valid;
  wire                PE74_valid;
  wire                PE75_valid;
  wire                PE76_valid;
  wire                PE77_valid;
  wire                PE78_valid;
  wire                PE79_valid;
  wire                PE710_valid;
  wire                PE711_valid;
  wire                PE712_valid;
  wire                PE713_valid;
  wire                PE714_valid;
  wire                PE715_valid;
  wire                PE716_valid;
  wire                PE717_valid;
  wire                PE718_valid;
  wire                PE719_valid;
  wire                PE720_valid;
  wire                PE721_valid;
  wire                PE722_valid;
  wire                PE723_valid;
  wire                PE724_valid;
  wire                PE725_valid;
  wire                PE726_valid;
  wire                PE727_valid;
  wire                PE728_valid;
  wire                PE729_valid;
  wire                PE730_valid;
  wire                PE731_valid;
  wire                PE732_valid;
  wire                PE733_valid;
  wire                PE734_valid;
  wire                PE735_valid;
  wire                PE736_valid;
  wire                PE737_valid;
  wire                PE738_valid;
  wire                PE739_valid;
  wire                PE740_valid;
  wire                PE741_valid;
  wire                PE742_valid;
  wire                PE743_valid;
  wire                PE744_valid;
  wire                PE745_valid;
  wire                PE746_valid;
  wire                PE747_valid;
  wire                PE748_valid;
  wire                PE749_valid;
  wire                PE750_valid;
  wire                PE751_valid;
  wire                PE752_valid;
  wire                PE753_valid;
  wire                PE754_valid;
  wire                PE755_valid;
  wire                PE756_valid;
  wire                PE757_valid;
  wire                PE758_valid;
  wire                PE759_valid;
  wire                PE760_valid;
  wire                PE761_valid;
  wire                PE762_valid;
  wire                PE763_valid;
  wire       [7:0]    PE00_acount;
  wire       [7:0]    PE00_bcount;
  wire       [31:0]   PE00_PE_OUT;
  wire                PE00_finish;
  wire       [7:0]    PE01_acount;
  wire       [7:0]    PE01_bcount;
  wire       [31:0]   PE01_PE_OUT;
  wire                PE01_finish;
  wire       [7:0]    PE02_acount;
  wire       [7:0]    PE02_bcount;
  wire       [31:0]   PE02_PE_OUT;
  wire                PE02_finish;
  wire       [7:0]    PE03_acount;
  wire       [7:0]    PE03_bcount;
  wire       [31:0]   PE03_PE_OUT;
  wire                PE03_finish;
  wire       [7:0]    PE04_acount;
  wire       [7:0]    PE04_bcount;
  wire       [31:0]   PE04_PE_OUT;
  wire                PE04_finish;
  wire       [7:0]    PE05_acount;
  wire       [7:0]    PE05_bcount;
  wire       [31:0]   PE05_PE_OUT;
  wire                PE05_finish;
  wire       [7:0]    PE06_acount;
  wire       [7:0]    PE06_bcount;
  wire       [31:0]   PE06_PE_OUT;
  wire                PE06_finish;
  wire       [7:0]    PE07_acount;
  wire       [7:0]    PE07_bcount;
  wire       [31:0]   PE07_PE_OUT;
  wire                PE07_finish;
  wire       [7:0]    PE08_acount;
  wire       [7:0]    PE08_bcount;
  wire       [31:0]   PE08_PE_OUT;
  wire                PE08_finish;
  wire       [7:0]    PE09_acount;
  wire       [7:0]    PE09_bcount;
  wire       [31:0]   PE09_PE_OUT;
  wire                PE09_finish;
  wire       [7:0]    PE010_acount;
  wire       [7:0]    PE010_bcount;
  wire       [31:0]   PE010_PE_OUT;
  wire                PE010_finish;
  wire       [7:0]    PE011_acount;
  wire       [7:0]    PE011_bcount;
  wire       [31:0]   PE011_PE_OUT;
  wire                PE011_finish;
  wire       [7:0]    PE012_acount;
  wire       [7:0]    PE012_bcount;
  wire       [31:0]   PE012_PE_OUT;
  wire                PE012_finish;
  wire       [7:0]    PE013_acount;
  wire       [7:0]    PE013_bcount;
  wire       [31:0]   PE013_PE_OUT;
  wire                PE013_finish;
  wire       [7:0]    PE014_acount;
  wire       [7:0]    PE014_bcount;
  wire       [31:0]   PE014_PE_OUT;
  wire                PE014_finish;
  wire       [7:0]    PE015_acount;
  wire       [7:0]    PE015_bcount;
  wire       [31:0]   PE015_PE_OUT;
  wire                PE015_finish;
  wire       [7:0]    PE016_acount;
  wire       [7:0]    PE016_bcount;
  wire       [31:0]   PE016_PE_OUT;
  wire                PE016_finish;
  wire       [7:0]    PE017_acount;
  wire       [7:0]    PE017_bcount;
  wire       [31:0]   PE017_PE_OUT;
  wire                PE017_finish;
  wire       [7:0]    PE018_acount;
  wire       [7:0]    PE018_bcount;
  wire       [31:0]   PE018_PE_OUT;
  wire                PE018_finish;
  wire       [7:0]    PE019_acount;
  wire       [7:0]    PE019_bcount;
  wire       [31:0]   PE019_PE_OUT;
  wire                PE019_finish;
  wire       [7:0]    PE020_acount;
  wire       [7:0]    PE020_bcount;
  wire       [31:0]   PE020_PE_OUT;
  wire                PE020_finish;
  wire       [7:0]    PE021_acount;
  wire       [7:0]    PE021_bcount;
  wire       [31:0]   PE021_PE_OUT;
  wire                PE021_finish;
  wire       [7:0]    PE022_acount;
  wire       [7:0]    PE022_bcount;
  wire       [31:0]   PE022_PE_OUT;
  wire                PE022_finish;
  wire       [7:0]    PE023_acount;
  wire       [7:0]    PE023_bcount;
  wire       [31:0]   PE023_PE_OUT;
  wire                PE023_finish;
  wire       [7:0]    PE024_acount;
  wire       [7:0]    PE024_bcount;
  wire       [31:0]   PE024_PE_OUT;
  wire                PE024_finish;
  wire       [7:0]    PE025_acount;
  wire       [7:0]    PE025_bcount;
  wire       [31:0]   PE025_PE_OUT;
  wire                PE025_finish;
  wire       [7:0]    PE026_acount;
  wire       [7:0]    PE026_bcount;
  wire       [31:0]   PE026_PE_OUT;
  wire                PE026_finish;
  wire       [7:0]    PE027_acount;
  wire       [7:0]    PE027_bcount;
  wire       [31:0]   PE027_PE_OUT;
  wire                PE027_finish;
  wire       [7:0]    PE028_acount;
  wire       [7:0]    PE028_bcount;
  wire       [31:0]   PE028_PE_OUT;
  wire                PE028_finish;
  wire       [7:0]    PE029_acount;
  wire       [7:0]    PE029_bcount;
  wire       [31:0]   PE029_PE_OUT;
  wire                PE029_finish;
  wire       [7:0]    PE030_acount;
  wire       [7:0]    PE030_bcount;
  wire       [31:0]   PE030_PE_OUT;
  wire                PE030_finish;
  wire       [7:0]    PE031_acount;
  wire       [7:0]    PE031_bcount;
  wire       [31:0]   PE031_PE_OUT;
  wire                PE031_finish;
  wire       [7:0]    PE032_acount;
  wire       [7:0]    PE032_bcount;
  wire       [31:0]   PE032_PE_OUT;
  wire                PE032_finish;
  wire       [7:0]    PE033_acount;
  wire       [7:0]    PE033_bcount;
  wire       [31:0]   PE033_PE_OUT;
  wire                PE033_finish;
  wire       [7:0]    PE034_acount;
  wire       [7:0]    PE034_bcount;
  wire       [31:0]   PE034_PE_OUT;
  wire                PE034_finish;
  wire       [7:0]    PE035_acount;
  wire       [7:0]    PE035_bcount;
  wire       [31:0]   PE035_PE_OUT;
  wire                PE035_finish;
  wire       [7:0]    PE036_acount;
  wire       [7:0]    PE036_bcount;
  wire       [31:0]   PE036_PE_OUT;
  wire                PE036_finish;
  wire       [7:0]    PE037_acount;
  wire       [7:0]    PE037_bcount;
  wire       [31:0]   PE037_PE_OUT;
  wire                PE037_finish;
  wire       [7:0]    PE038_acount;
  wire       [7:0]    PE038_bcount;
  wire       [31:0]   PE038_PE_OUT;
  wire                PE038_finish;
  wire       [7:0]    PE039_acount;
  wire       [7:0]    PE039_bcount;
  wire       [31:0]   PE039_PE_OUT;
  wire                PE039_finish;
  wire       [7:0]    PE040_acount;
  wire       [7:0]    PE040_bcount;
  wire       [31:0]   PE040_PE_OUT;
  wire                PE040_finish;
  wire       [7:0]    PE041_acount;
  wire       [7:0]    PE041_bcount;
  wire       [31:0]   PE041_PE_OUT;
  wire                PE041_finish;
  wire       [7:0]    PE042_acount;
  wire       [7:0]    PE042_bcount;
  wire       [31:0]   PE042_PE_OUT;
  wire                PE042_finish;
  wire       [7:0]    PE043_acount;
  wire       [7:0]    PE043_bcount;
  wire       [31:0]   PE043_PE_OUT;
  wire                PE043_finish;
  wire       [7:0]    PE044_acount;
  wire       [7:0]    PE044_bcount;
  wire       [31:0]   PE044_PE_OUT;
  wire                PE044_finish;
  wire       [7:0]    PE045_acount;
  wire       [7:0]    PE045_bcount;
  wire       [31:0]   PE045_PE_OUT;
  wire                PE045_finish;
  wire       [7:0]    PE046_acount;
  wire       [7:0]    PE046_bcount;
  wire       [31:0]   PE046_PE_OUT;
  wire                PE046_finish;
  wire       [7:0]    PE047_acount;
  wire       [7:0]    PE047_bcount;
  wire       [31:0]   PE047_PE_OUT;
  wire                PE047_finish;
  wire       [7:0]    PE048_acount;
  wire       [7:0]    PE048_bcount;
  wire       [31:0]   PE048_PE_OUT;
  wire                PE048_finish;
  wire       [7:0]    PE049_acount;
  wire       [7:0]    PE049_bcount;
  wire       [31:0]   PE049_PE_OUT;
  wire                PE049_finish;
  wire       [7:0]    PE050_acount;
  wire       [7:0]    PE050_bcount;
  wire       [31:0]   PE050_PE_OUT;
  wire                PE050_finish;
  wire       [7:0]    PE051_acount;
  wire       [7:0]    PE051_bcount;
  wire       [31:0]   PE051_PE_OUT;
  wire                PE051_finish;
  wire       [7:0]    PE052_acount;
  wire       [7:0]    PE052_bcount;
  wire       [31:0]   PE052_PE_OUT;
  wire                PE052_finish;
  wire       [7:0]    PE053_acount;
  wire       [7:0]    PE053_bcount;
  wire       [31:0]   PE053_PE_OUT;
  wire                PE053_finish;
  wire       [7:0]    PE054_acount;
  wire       [7:0]    PE054_bcount;
  wire       [31:0]   PE054_PE_OUT;
  wire                PE054_finish;
  wire       [7:0]    PE055_acount;
  wire       [7:0]    PE055_bcount;
  wire       [31:0]   PE055_PE_OUT;
  wire                PE055_finish;
  wire       [7:0]    PE056_acount;
  wire       [7:0]    PE056_bcount;
  wire       [31:0]   PE056_PE_OUT;
  wire                PE056_finish;
  wire       [7:0]    PE057_acount;
  wire       [7:0]    PE057_bcount;
  wire       [31:0]   PE057_PE_OUT;
  wire                PE057_finish;
  wire       [7:0]    PE058_acount;
  wire       [7:0]    PE058_bcount;
  wire       [31:0]   PE058_PE_OUT;
  wire                PE058_finish;
  wire       [7:0]    PE059_acount;
  wire       [7:0]    PE059_bcount;
  wire       [31:0]   PE059_PE_OUT;
  wire                PE059_finish;
  wire       [7:0]    PE060_acount;
  wire       [7:0]    PE060_bcount;
  wire       [31:0]   PE060_PE_OUT;
  wire                PE060_finish;
  wire       [7:0]    PE061_acount;
  wire       [7:0]    PE061_bcount;
  wire       [31:0]   PE061_PE_OUT;
  wire                PE061_finish;
  wire       [7:0]    PE062_acount;
  wire       [7:0]    PE062_bcount;
  wire       [31:0]   PE062_PE_OUT;
  wire                PE062_finish;
  wire       [7:0]    PE063_acount;
  wire       [7:0]    PE063_bcount;
  wire       [31:0]   PE063_PE_OUT;
  wire                PE063_finish;
  wire       [7:0]    PE10_acount;
  wire       [7:0]    PE10_bcount;
  wire       [31:0]   PE10_PE_OUT;
  wire                PE10_finish;
  wire       [7:0]    PE11_acount;
  wire       [7:0]    PE11_bcount;
  wire       [31:0]   PE11_PE_OUT;
  wire                PE11_finish;
  wire       [7:0]    PE12_acount;
  wire       [7:0]    PE12_bcount;
  wire       [31:0]   PE12_PE_OUT;
  wire                PE12_finish;
  wire       [7:0]    PE13_acount;
  wire       [7:0]    PE13_bcount;
  wire       [31:0]   PE13_PE_OUT;
  wire                PE13_finish;
  wire       [7:0]    PE14_acount;
  wire       [7:0]    PE14_bcount;
  wire       [31:0]   PE14_PE_OUT;
  wire                PE14_finish;
  wire       [7:0]    PE15_acount;
  wire       [7:0]    PE15_bcount;
  wire       [31:0]   PE15_PE_OUT;
  wire                PE15_finish;
  wire       [7:0]    PE16_acount;
  wire       [7:0]    PE16_bcount;
  wire       [31:0]   PE16_PE_OUT;
  wire                PE16_finish;
  wire       [7:0]    PE17_acount;
  wire       [7:0]    PE17_bcount;
  wire       [31:0]   PE17_PE_OUT;
  wire                PE17_finish;
  wire       [7:0]    PE18_acount;
  wire       [7:0]    PE18_bcount;
  wire       [31:0]   PE18_PE_OUT;
  wire                PE18_finish;
  wire       [7:0]    PE19_acount;
  wire       [7:0]    PE19_bcount;
  wire       [31:0]   PE19_PE_OUT;
  wire                PE19_finish;
  wire       [7:0]    PE110_acount;
  wire       [7:0]    PE110_bcount;
  wire       [31:0]   PE110_PE_OUT;
  wire                PE110_finish;
  wire       [7:0]    PE111_acount;
  wire       [7:0]    PE111_bcount;
  wire       [31:0]   PE111_PE_OUT;
  wire                PE111_finish;
  wire       [7:0]    PE112_acount;
  wire       [7:0]    PE112_bcount;
  wire       [31:0]   PE112_PE_OUT;
  wire                PE112_finish;
  wire       [7:0]    PE113_acount;
  wire       [7:0]    PE113_bcount;
  wire       [31:0]   PE113_PE_OUT;
  wire                PE113_finish;
  wire       [7:0]    PE114_acount;
  wire       [7:0]    PE114_bcount;
  wire       [31:0]   PE114_PE_OUT;
  wire                PE114_finish;
  wire       [7:0]    PE115_acount;
  wire       [7:0]    PE115_bcount;
  wire       [31:0]   PE115_PE_OUT;
  wire                PE115_finish;
  wire       [7:0]    PE116_acount;
  wire       [7:0]    PE116_bcount;
  wire       [31:0]   PE116_PE_OUT;
  wire                PE116_finish;
  wire       [7:0]    PE117_acount;
  wire       [7:0]    PE117_bcount;
  wire       [31:0]   PE117_PE_OUT;
  wire                PE117_finish;
  wire       [7:0]    PE118_acount;
  wire       [7:0]    PE118_bcount;
  wire       [31:0]   PE118_PE_OUT;
  wire                PE118_finish;
  wire       [7:0]    PE119_acount;
  wire       [7:0]    PE119_bcount;
  wire       [31:0]   PE119_PE_OUT;
  wire                PE119_finish;
  wire       [7:0]    PE120_acount;
  wire       [7:0]    PE120_bcount;
  wire       [31:0]   PE120_PE_OUT;
  wire                PE120_finish;
  wire       [7:0]    PE121_acount;
  wire       [7:0]    PE121_bcount;
  wire       [31:0]   PE121_PE_OUT;
  wire                PE121_finish;
  wire       [7:0]    PE122_acount;
  wire       [7:0]    PE122_bcount;
  wire       [31:0]   PE122_PE_OUT;
  wire                PE122_finish;
  wire       [7:0]    PE123_acount;
  wire       [7:0]    PE123_bcount;
  wire       [31:0]   PE123_PE_OUT;
  wire                PE123_finish;
  wire       [7:0]    PE124_acount;
  wire       [7:0]    PE124_bcount;
  wire       [31:0]   PE124_PE_OUT;
  wire                PE124_finish;
  wire       [7:0]    PE125_acount;
  wire       [7:0]    PE125_bcount;
  wire       [31:0]   PE125_PE_OUT;
  wire                PE125_finish;
  wire       [7:0]    PE126_acount;
  wire       [7:0]    PE126_bcount;
  wire       [31:0]   PE126_PE_OUT;
  wire                PE126_finish;
  wire       [7:0]    PE127_acount;
  wire       [7:0]    PE127_bcount;
  wire       [31:0]   PE127_PE_OUT;
  wire                PE127_finish;
  wire       [7:0]    PE128_acount;
  wire       [7:0]    PE128_bcount;
  wire       [31:0]   PE128_PE_OUT;
  wire                PE128_finish;
  wire       [7:0]    PE129_acount;
  wire       [7:0]    PE129_bcount;
  wire       [31:0]   PE129_PE_OUT;
  wire                PE129_finish;
  wire       [7:0]    PE130_acount;
  wire       [7:0]    PE130_bcount;
  wire       [31:0]   PE130_PE_OUT;
  wire                PE130_finish;
  wire       [7:0]    PE131_acount;
  wire       [7:0]    PE131_bcount;
  wire       [31:0]   PE131_PE_OUT;
  wire                PE131_finish;
  wire       [7:0]    PE132_acount;
  wire       [7:0]    PE132_bcount;
  wire       [31:0]   PE132_PE_OUT;
  wire                PE132_finish;
  wire       [7:0]    PE133_acount;
  wire       [7:0]    PE133_bcount;
  wire       [31:0]   PE133_PE_OUT;
  wire                PE133_finish;
  wire       [7:0]    PE134_acount;
  wire       [7:0]    PE134_bcount;
  wire       [31:0]   PE134_PE_OUT;
  wire                PE134_finish;
  wire       [7:0]    PE135_acount;
  wire       [7:0]    PE135_bcount;
  wire       [31:0]   PE135_PE_OUT;
  wire                PE135_finish;
  wire       [7:0]    PE136_acount;
  wire       [7:0]    PE136_bcount;
  wire       [31:0]   PE136_PE_OUT;
  wire                PE136_finish;
  wire       [7:0]    PE137_acount;
  wire       [7:0]    PE137_bcount;
  wire       [31:0]   PE137_PE_OUT;
  wire                PE137_finish;
  wire       [7:0]    PE138_acount;
  wire       [7:0]    PE138_bcount;
  wire       [31:0]   PE138_PE_OUT;
  wire                PE138_finish;
  wire       [7:0]    PE139_acount;
  wire       [7:0]    PE139_bcount;
  wire       [31:0]   PE139_PE_OUT;
  wire                PE139_finish;
  wire       [7:0]    PE140_acount;
  wire       [7:0]    PE140_bcount;
  wire       [31:0]   PE140_PE_OUT;
  wire                PE140_finish;
  wire       [7:0]    PE141_acount;
  wire       [7:0]    PE141_bcount;
  wire       [31:0]   PE141_PE_OUT;
  wire                PE141_finish;
  wire       [7:0]    PE142_acount;
  wire       [7:0]    PE142_bcount;
  wire       [31:0]   PE142_PE_OUT;
  wire                PE142_finish;
  wire       [7:0]    PE143_acount;
  wire       [7:0]    PE143_bcount;
  wire       [31:0]   PE143_PE_OUT;
  wire                PE143_finish;
  wire       [7:0]    PE144_acount;
  wire       [7:0]    PE144_bcount;
  wire       [31:0]   PE144_PE_OUT;
  wire                PE144_finish;
  wire       [7:0]    PE145_acount;
  wire       [7:0]    PE145_bcount;
  wire       [31:0]   PE145_PE_OUT;
  wire                PE145_finish;
  wire       [7:0]    PE146_acount;
  wire       [7:0]    PE146_bcount;
  wire       [31:0]   PE146_PE_OUT;
  wire                PE146_finish;
  wire       [7:0]    PE147_acount;
  wire       [7:0]    PE147_bcount;
  wire       [31:0]   PE147_PE_OUT;
  wire                PE147_finish;
  wire       [7:0]    PE148_acount;
  wire       [7:0]    PE148_bcount;
  wire       [31:0]   PE148_PE_OUT;
  wire                PE148_finish;
  wire       [7:0]    PE149_acount;
  wire       [7:0]    PE149_bcount;
  wire       [31:0]   PE149_PE_OUT;
  wire                PE149_finish;
  wire       [7:0]    PE150_acount;
  wire       [7:0]    PE150_bcount;
  wire       [31:0]   PE150_PE_OUT;
  wire                PE150_finish;
  wire       [7:0]    PE151_acount;
  wire       [7:0]    PE151_bcount;
  wire       [31:0]   PE151_PE_OUT;
  wire                PE151_finish;
  wire       [7:0]    PE152_acount;
  wire       [7:0]    PE152_bcount;
  wire       [31:0]   PE152_PE_OUT;
  wire                PE152_finish;
  wire       [7:0]    PE153_acount;
  wire       [7:0]    PE153_bcount;
  wire       [31:0]   PE153_PE_OUT;
  wire                PE153_finish;
  wire       [7:0]    PE154_acount;
  wire       [7:0]    PE154_bcount;
  wire       [31:0]   PE154_PE_OUT;
  wire                PE154_finish;
  wire       [7:0]    PE155_acount;
  wire       [7:0]    PE155_bcount;
  wire       [31:0]   PE155_PE_OUT;
  wire                PE155_finish;
  wire       [7:0]    PE156_acount;
  wire       [7:0]    PE156_bcount;
  wire       [31:0]   PE156_PE_OUT;
  wire                PE156_finish;
  wire       [7:0]    PE157_acount;
  wire       [7:0]    PE157_bcount;
  wire       [31:0]   PE157_PE_OUT;
  wire                PE157_finish;
  wire       [7:0]    PE158_acount;
  wire       [7:0]    PE158_bcount;
  wire       [31:0]   PE158_PE_OUT;
  wire                PE158_finish;
  wire       [7:0]    PE159_acount;
  wire       [7:0]    PE159_bcount;
  wire       [31:0]   PE159_PE_OUT;
  wire                PE159_finish;
  wire       [7:0]    PE160_acount;
  wire       [7:0]    PE160_bcount;
  wire       [31:0]   PE160_PE_OUT;
  wire                PE160_finish;
  wire       [7:0]    PE161_acount;
  wire       [7:0]    PE161_bcount;
  wire       [31:0]   PE161_PE_OUT;
  wire                PE161_finish;
  wire       [7:0]    PE162_acount;
  wire       [7:0]    PE162_bcount;
  wire       [31:0]   PE162_PE_OUT;
  wire                PE162_finish;
  wire       [7:0]    PE163_acount;
  wire       [7:0]    PE163_bcount;
  wire       [31:0]   PE163_PE_OUT;
  wire                PE163_finish;
  wire       [7:0]    PE20_acount;
  wire       [7:0]    PE20_bcount;
  wire       [31:0]   PE20_PE_OUT;
  wire                PE20_finish;
  wire       [7:0]    PE21_acount;
  wire       [7:0]    PE21_bcount;
  wire       [31:0]   PE21_PE_OUT;
  wire                PE21_finish;
  wire       [7:0]    PE22_acount;
  wire       [7:0]    PE22_bcount;
  wire       [31:0]   PE22_PE_OUT;
  wire                PE22_finish;
  wire       [7:0]    PE23_acount;
  wire       [7:0]    PE23_bcount;
  wire       [31:0]   PE23_PE_OUT;
  wire                PE23_finish;
  wire       [7:0]    PE24_acount;
  wire       [7:0]    PE24_bcount;
  wire       [31:0]   PE24_PE_OUT;
  wire                PE24_finish;
  wire       [7:0]    PE25_acount;
  wire       [7:0]    PE25_bcount;
  wire       [31:0]   PE25_PE_OUT;
  wire                PE25_finish;
  wire       [7:0]    PE26_acount;
  wire       [7:0]    PE26_bcount;
  wire       [31:0]   PE26_PE_OUT;
  wire                PE26_finish;
  wire       [7:0]    PE27_acount;
  wire       [7:0]    PE27_bcount;
  wire       [31:0]   PE27_PE_OUT;
  wire                PE27_finish;
  wire       [7:0]    PE28_acount;
  wire       [7:0]    PE28_bcount;
  wire       [31:0]   PE28_PE_OUT;
  wire                PE28_finish;
  wire       [7:0]    PE29_acount;
  wire       [7:0]    PE29_bcount;
  wire       [31:0]   PE29_PE_OUT;
  wire                PE29_finish;
  wire       [7:0]    PE210_acount;
  wire       [7:0]    PE210_bcount;
  wire       [31:0]   PE210_PE_OUT;
  wire                PE210_finish;
  wire       [7:0]    PE211_acount;
  wire       [7:0]    PE211_bcount;
  wire       [31:0]   PE211_PE_OUT;
  wire                PE211_finish;
  wire       [7:0]    PE212_acount;
  wire       [7:0]    PE212_bcount;
  wire       [31:0]   PE212_PE_OUT;
  wire                PE212_finish;
  wire       [7:0]    PE213_acount;
  wire       [7:0]    PE213_bcount;
  wire       [31:0]   PE213_PE_OUT;
  wire                PE213_finish;
  wire       [7:0]    PE214_acount;
  wire       [7:0]    PE214_bcount;
  wire       [31:0]   PE214_PE_OUT;
  wire                PE214_finish;
  wire       [7:0]    PE215_acount;
  wire       [7:0]    PE215_bcount;
  wire       [31:0]   PE215_PE_OUT;
  wire                PE215_finish;
  wire       [7:0]    PE216_acount;
  wire       [7:0]    PE216_bcount;
  wire       [31:0]   PE216_PE_OUT;
  wire                PE216_finish;
  wire       [7:0]    PE217_acount;
  wire       [7:0]    PE217_bcount;
  wire       [31:0]   PE217_PE_OUT;
  wire                PE217_finish;
  wire       [7:0]    PE218_acount;
  wire       [7:0]    PE218_bcount;
  wire       [31:0]   PE218_PE_OUT;
  wire                PE218_finish;
  wire       [7:0]    PE219_acount;
  wire       [7:0]    PE219_bcount;
  wire       [31:0]   PE219_PE_OUT;
  wire                PE219_finish;
  wire       [7:0]    PE220_acount;
  wire       [7:0]    PE220_bcount;
  wire       [31:0]   PE220_PE_OUT;
  wire                PE220_finish;
  wire       [7:0]    PE221_acount;
  wire       [7:0]    PE221_bcount;
  wire       [31:0]   PE221_PE_OUT;
  wire                PE221_finish;
  wire       [7:0]    PE222_acount;
  wire       [7:0]    PE222_bcount;
  wire       [31:0]   PE222_PE_OUT;
  wire                PE222_finish;
  wire       [7:0]    PE223_acount;
  wire       [7:0]    PE223_bcount;
  wire       [31:0]   PE223_PE_OUT;
  wire                PE223_finish;
  wire       [7:0]    PE224_acount;
  wire       [7:0]    PE224_bcount;
  wire       [31:0]   PE224_PE_OUT;
  wire                PE224_finish;
  wire       [7:0]    PE225_acount;
  wire       [7:0]    PE225_bcount;
  wire       [31:0]   PE225_PE_OUT;
  wire                PE225_finish;
  wire       [7:0]    PE226_acount;
  wire       [7:0]    PE226_bcount;
  wire       [31:0]   PE226_PE_OUT;
  wire                PE226_finish;
  wire       [7:0]    PE227_acount;
  wire       [7:0]    PE227_bcount;
  wire       [31:0]   PE227_PE_OUT;
  wire                PE227_finish;
  wire       [7:0]    PE228_acount;
  wire       [7:0]    PE228_bcount;
  wire       [31:0]   PE228_PE_OUT;
  wire                PE228_finish;
  wire       [7:0]    PE229_acount;
  wire       [7:0]    PE229_bcount;
  wire       [31:0]   PE229_PE_OUT;
  wire                PE229_finish;
  wire       [7:0]    PE230_acount;
  wire       [7:0]    PE230_bcount;
  wire       [31:0]   PE230_PE_OUT;
  wire                PE230_finish;
  wire       [7:0]    PE231_acount;
  wire       [7:0]    PE231_bcount;
  wire       [31:0]   PE231_PE_OUT;
  wire                PE231_finish;
  wire       [7:0]    PE232_acount;
  wire       [7:0]    PE232_bcount;
  wire       [31:0]   PE232_PE_OUT;
  wire                PE232_finish;
  wire       [7:0]    PE233_acount;
  wire       [7:0]    PE233_bcount;
  wire       [31:0]   PE233_PE_OUT;
  wire                PE233_finish;
  wire       [7:0]    PE234_acount;
  wire       [7:0]    PE234_bcount;
  wire       [31:0]   PE234_PE_OUT;
  wire                PE234_finish;
  wire       [7:0]    PE235_acount;
  wire       [7:0]    PE235_bcount;
  wire       [31:0]   PE235_PE_OUT;
  wire                PE235_finish;
  wire       [7:0]    PE236_acount;
  wire       [7:0]    PE236_bcount;
  wire       [31:0]   PE236_PE_OUT;
  wire                PE236_finish;
  wire       [7:0]    PE237_acount;
  wire       [7:0]    PE237_bcount;
  wire       [31:0]   PE237_PE_OUT;
  wire                PE237_finish;
  wire       [7:0]    PE238_acount;
  wire       [7:0]    PE238_bcount;
  wire       [31:0]   PE238_PE_OUT;
  wire                PE238_finish;
  wire       [7:0]    PE239_acount;
  wire       [7:0]    PE239_bcount;
  wire       [31:0]   PE239_PE_OUT;
  wire                PE239_finish;
  wire       [7:0]    PE240_acount;
  wire       [7:0]    PE240_bcount;
  wire       [31:0]   PE240_PE_OUT;
  wire                PE240_finish;
  wire       [7:0]    PE241_acount;
  wire       [7:0]    PE241_bcount;
  wire       [31:0]   PE241_PE_OUT;
  wire                PE241_finish;
  wire       [7:0]    PE242_acount;
  wire       [7:0]    PE242_bcount;
  wire       [31:0]   PE242_PE_OUT;
  wire                PE242_finish;
  wire       [7:0]    PE243_acount;
  wire       [7:0]    PE243_bcount;
  wire       [31:0]   PE243_PE_OUT;
  wire                PE243_finish;
  wire       [7:0]    PE244_acount;
  wire       [7:0]    PE244_bcount;
  wire       [31:0]   PE244_PE_OUT;
  wire                PE244_finish;
  wire       [7:0]    PE245_acount;
  wire       [7:0]    PE245_bcount;
  wire       [31:0]   PE245_PE_OUT;
  wire                PE245_finish;
  wire       [7:0]    PE246_acount;
  wire       [7:0]    PE246_bcount;
  wire       [31:0]   PE246_PE_OUT;
  wire                PE246_finish;
  wire       [7:0]    PE247_acount;
  wire       [7:0]    PE247_bcount;
  wire       [31:0]   PE247_PE_OUT;
  wire                PE247_finish;
  wire       [7:0]    PE248_acount;
  wire       [7:0]    PE248_bcount;
  wire       [31:0]   PE248_PE_OUT;
  wire                PE248_finish;
  wire       [7:0]    PE249_acount;
  wire       [7:0]    PE249_bcount;
  wire       [31:0]   PE249_PE_OUT;
  wire                PE249_finish;
  wire       [7:0]    PE250_acount;
  wire       [7:0]    PE250_bcount;
  wire       [31:0]   PE250_PE_OUT;
  wire                PE250_finish;
  wire       [7:0]    PE251_acount;
  wire       [7:0]    PE251_bcount;
  wire       [31:0]   PE251_PE_OUT;
  wire                PE251_finish;
  wire       [7:0]    PE252_acount;
  wire       [7:0]    PE252_bcount;
  wire       [31:0]   PE252_PE_OUT;
  wire                PE252_finish;
  wire       [7:0]    PE253_acount;
  wire       [7:0]    PE253_bcount;
  wire       [31:0]   PE253_PE_OUT;
  wire                PE253_finish;
  wire       [7:0]    PE254_acount;
  wire       [7:0]    PE254_bcount;
  wire       [31:0]   PE254_PE_OUT;
  wire                PE254_finish;
  wire       [7:0]    PE255_acount;
  wire       [7:0]    PE255_bcount;
  wire       [31:0]   PE255_PE_OUT;
  wire                PE255_finish;
  wire       [7:0]    PE256_acount;
  wire       [7:0]    PE256_bcount;
  wire       [31:0]   PE256_PE_OUT;
  wire                PE256_finish;
  wire       [7:0]    PE257_acount;
  wire       [7:0]    PE257_bcount;
  wire       [31:0]   PE257_PE_OUT;
  wire                PE257_finish;
  wire       [7:0]    PE258_acount;
  wire       [7:0]    PE258_bcount;
  wire       [31:0]   PE258_PE_OUT;
  wire                PE258_finish;
  wire       [7:0]    PE259_acount;
  wire       [7:0]    PE259_bcount;
  wire       [31:0]   PE259_PE_OUT;
  wire                PE259_finish;
  wire       [7:0]    PE260_acount;
  wire       [7:0]    PE260_bcount;
  wire       [31:0]   PE260_PE_OUT;
  wire                PE260_finish;
  wire       [7:0]    PE261_acount;
  wire       [7:0]    PE261_bcount;
  wire       [31:0]   PE261_PE_OUT;
  wire                PE261_finish;
  wire       [7:0]    PE262_acount;
  wire       [7:0]    PE262_bcount;
  wire       [31:0]   PE262_PE_OUT;
  wire                PE262_finish;
  wire       [7:0]    PE263_acount;
  wire       [7:0]    PE263_bcount;
  wire       [31:0]   PE263_PE_OUT;
  wire                PE263_finish;
  wire       [7:0]    PE30_acount;
  wire       [7:0]    PE30_bcount;
  wire       [31:0]   PE30_PE_OUT;
  wire                PE30_finish;
  wire       [7:0]    PE31_acount;
  wire       [7:0]    PE31_bcount;
  wire       [31:0]   PE31_PE_OUT;
  wire                PE31_finish;
  wire       [7:0]    PE32_acount;
  wire       [7:0]    PE32_bcount;
  wire       [31:0]   PE32_PE_OUT;
  wire                PE32_finish;
  wire       [7:0]    PE33_acount;
  wire       [7:0]    PE33_bcount;
  wire       [31:0]   PE33_PE_OUT;
  wire                PE33_finish;
  wire       [7:0]    PE34_acount;
  wire       [7:0]    PE34_bcount;
  wire       [31:0]   PE34_PE_OUT;
  wire                PE34_finish;
  wire       [7:0]    PE35_acount;
  wire       [7:0]    PE35_bcount;
  wire       [31:0]   PE35_PE_OUT;
  wire                PE35_finish;
  wire       [7:0]    PE36_acount;
  wire       [7:0]    PE36_bcount;
  wire       [31:0]   PE36_PE_OUT;
  wire                PE36_finish;
  wire       [7:0]    PE37_acount;
  wire       [7:0]    PE37_bcount;
  wire       [31:0]   PE37_PE_OUT;
  wire                PE37_finish;
  wire       [7:0]    PE38_acount;
  wire       [7:0]    PE38_bcount;
  wire       [31:0]   PE38_PE_OUT;
  wire                PE38_finish;
  wire       [7:0]    PE39_acount;
  wire       [7:0]    PE39_bcount;
  wire       [31:0]   PE39_PE_OUT;
  wire                PE39_finish;
  wire       [7:0]    PE310_acount;
  wire       [7:0]    PE310_bcount;
  wire       [31:0]   PE310_PE_OUT;
  wire                PE310_finish;
  wire       [7:0]    PE311_acount;
  wire       [7:0]    PE311_bcount;
  wire       [31:0]   PE311_PE_OUT;
  wire                PE311_finish;
  wire       [7:0]    PE312_acount;
  wire       [7:0]    PE312_bcount;
  wire       [31:0]   PE312_PE_OUT;
  wire                PE312_finish;
  wire       [7:0]    PE313_acount;
  wire       [7:0]    PE313_bcount;
  wire       [31:0]   PE313_PE_OUT;
  wire                PE313_finish;
  wire       [7:0]    PE314_acount;
  wire       [7:0]    PE314_bcount;
  wire       [31:0]   PE314_PE_OUT;
  wire                PE314_finish;
  wire       [7:0]    PE315_acount;
  wire       [7:0]    PE315_bcount;
  wire       [31:0]   PE315_PE_OUT;
  wire                PE315_finish;
  wire       [7:0]    PE316_acount;
  wire       [7:0]    PE316_bcount;
  wire       [31:0]   PE316_PE_OUT;
  wire                PE316_finish;
  wire       [7:0]    PE317_acount;
  wire       [7:0]    PE317_bcount;
  wire       [31:0]   PE317_PE_OUT;
  wire                PE317_finish;
  wire       [7:0]    PE318_acount;
  wire       [7:0]    PE318_bcount;
  wire       [31:0]   PE318_PE_OUT;
  wire                PE318_finish;
  wire       [7:0]    PE319_acount;
  wire       [7:0]    PE319_bcount;
  wire       [31:0]   PE319_PE_OUT;
  wire                PE319_finish;
  wire       [7:0]    PE320_acount;
  wire       [7:0]    PE320_bcount;
  wire       [31:0]   PE320_PE_OUT;
  wire                PE320_finish;
  wire       [7:0]    PE321_acount;
  wire       [7:0]    PE321_bcount;
  wire       [31:0]   PE321_PE_OUT;
  wire                PE321_finish;
  wire       [7:0]    PE322_acount;
  wire       [7:0]    PE322_bcount;
  wire       [31:0]   PE322_PE_OUT;
  wire                PE322_finish;
  wire       [7:0]    PE323_acount;
  wire       [7:0]    PE323_bcount;
  wire       [31:0]   PE323_PE_OUT;
  wire                PE323_finish;
  wire       [7:0]    PE324_acount;
  wire       [7:0]    PE324_bcount;
  wire       [31:0]   PE324_PE_OUT;
  wire                PE324_finish;
  wire       [7:0]    PE325_acount;
  wire       [7:0]    PE325_bcount;
  wire       [31:0]   PE325_PE_OUT;
  wire                PE325_finish;
  wire       [7:0]    PE326_acount;
  wire       [7:0]    PE326_bcount;
  wire       [31:0]   PE326_PE_OUT;
  wire                PE326_finish;
  wire       [7:0]    PE327_acount;
  wire       [7:0]    PE327_bcount;
  wire       [31:0]   PE327_PE_OUT;
  wire                PE327_finish;
  wire       [7:0]    PE328_acount;
  wire       [7:0]    PE328_bcount;
  wire       [31:0]   PE328_PE_OUT;
  wire                PE328_finish;
  wire       [7:0]    PE329_acount;
  wire       [7:0]    PE329_bcount;
  wire       [31:0]   PE329_PE_OUT;
  wire                PE329_finish;
  wire       [7:0]    PE330_acount;
  wire       [7:0]    PE330_bcount;
  wire       [31:0]   PE330_PE_OUT;
  wire                PE330_finish;
  wire       [7:0]    PE331_acount;
  wire       [7:0]    PE331_bcount;
  wire       [31:0]   PE331_PE_OUT;
  wire                PE331_finish;
  wire       [7:0]    PE332_acount;
  wire       [7:0]    PE332_bcount;
  wire       [31:0]   PE332_PE_OUT;
  wire                PE332_finish;
  wire       [7:0]    PE333_acount;
  wire       [7:0]    PE333_bcount;
  wire       [31:0]   PE333_PE_OUT;
  wire                PE333_finish;
  wire       [7:0]    PE334_acount;
  wire       [7:0]    PE334_bcount;
  wire       [31:0]   PE334_PE_OUT;
  wire                PE334_finish;
  wire       [7:0]    PE335_acount;
  wire       [7:0]    PE335_bcount;
  wire       [31:0]   PE335_PE_OUT;
  wire                PE335_finish;
  wire       [7:0]    PE336_acount;
  wire       [7:0]    PE336_bcount;
  wire       [31:0]   PE336_PE_OUT;
  wire                PE336_finish;
  wire       [7:0]    PE337_acount;
  wire       [7:0]    PE337_bcount;
  wire       [31:0]   PE337_PE_OUT;
  wire                PE337_finish;
  wire       [7:0]    PE338_acount;
  wire       [7:0]    PE338_bcount;
  wire       [31:0]   PE338_PE_OUT;
  wire                PE338_finish;
  wire       [7:0]    PE339_acount;
  wire       [7:0]    PE339_bcount;
  wire       [31:0]   PE339_PE_OUT;
  wire                PE339_finish;
  wire       [7:0]    PE340_acount;
  wire       [7:0]    PE340_bcount;
  wire       [31:0]   PE340_PE_OUT;
  wire                PE340_finish;
  wire       [7:0]    PE341_acount;
  wire       [7:0]    PE341_bcount;
  wire       [31:0]   PE341_PE_OUT;
  wire                PE341_finish;
  wire       [7:0]    PE342_acount;
  wire       [7:0]    PE342_bcount;
  wire       [31:0]   PE342_PE_OUT;
  wire                PE342_finish;
  wire       [7:0]    PE343_acount;
  wire       [7:0]    PE343_bcount;
  wire       [31:0]   PE343_PE_OUT;
  wire                PE343_finish;
  wire       [7:0]    PE344_acount;
  wire       [7:0]    PE344_bcount;
  wire       [31:0]   PE344_PE_OUT;
  wire                PE344_finish;
  wire       [7:0]    PE345_acount;
  wire       [7:0]    PE345_bcount;
  wire       [31:0]   PE345_PE_OUT;
  wire                PE345_finish;
  wire       [7:0]    PE346_acount;
  wire       [7:0]    PE346_bcount;
  wire       [31:0]   PE346_PE_OUT;
  wire                PE346_finish;
  wire       [7:0]    PE347_acount;
  wire       [7:0]    PE347_bcount;
  wire       [31:0]   PE347_PE_OUT;
  wire                PE347_finish;
  wire       [7:0]    PE348_acount;
  wire       [7:0]    PE348_bcount;
  wire       [31:0]   PE348_PE_OUT;
  wire                PE348_finish;
  wire       [7:0]    PE349_acount;
  wire       [7:0]    PE349_bcount;
  wire       [31:0]   PE349_PE_OUT;
  wire                PE349_finish;
  wire       [7:0]    PE350_acount;
  wire       [7:0]    PE350_bcount;
  wire       [31:0]   PE350_PE_OUT;
  wire                PE350_finish;
  wire       [7:0]    PE351_acount;
  wire       [7:0]    PE351_bcount;
  wire       [31:0]   PE351_PE_OUT;
  wire                PE351_finish;
  wire       [7:0]    PE352_acount;
  wire       [7:0]    PE352_bcount;
  wire       [31:0]   PE352_PE_OUT;
  wire                PE352_finish;
  wire       [7:0]    PE353_acount;
  wire       [7:0]    PE353_bcount;
  wire       [31:0]   PE353_PE_OUT;
  wire                PE353_finish;
  wire       [7:0]    PE354_acount;
  wire       [7:0]    PE354_bcount;
  wire       [31:0]   PE354_PE_OUT;
  wire                PE354_finish;
  wire       [7:0]    PE355_acount;
  wire       [7:0]    PE355_bcount;
  wire       [31:0]   PE355_PE_OUT;
  wire                PE355_finish;
  wire       [7:0]    PE356_acount;
  wire       [7:0]    PE356_bcount;
  wire       [31:0]   PE356_PE_OUT;
  wire                PE356_finish;
  wire       [7:0]    PE357_acount;
  wire       [7:0]    PE357_bcount;
  wire       [31:0]   PE357_PE_OUT;
  wire                PE357_finish;
  wire       [7:0]    PE358_acount;
  wire       [7:0]    PE358_bcount;
  wire       [31:0]   PE358_PE_OUT;
  wire                PE358_finish;
  wire       [7:0]    PE359_acount;
  wire       [7:0]    PE359_bcount;
  wire       [31:0]   PE359_PE_OUT;
  wire                PE359_finish;
  wire       [7:0]    PE360_acount;
  wire       [7:0]    PE360_bcount;
  wire       [31:0]   PE360_PE_OUT;
  wire                PE360_finish;
  wire       [7:0]    PE361_acount;
  wire       [7:0]    PE361_bcount;
  wire       [31:0]   PE361_PE_OUT;
  wire                PE361_finish;
  wire       [7:0]    PE362_acount;
  wire       [7:0]    PE362_bcount;
  wire       [31:0]   PE362_PE_OUT;
  wire                PE362_finish;
  wire       [7:0]    PE363_acount;
  wire       [7:0]    PE363_bcount;
  wire       [31:0]   PE363_PE_OUT;
  wire                PE363_finish;
  wire       [7:0]    PE40_acount;
  wire       [7:0]    PE40_bcount;
  wire       [31:0]   PE40_PE_OUT;
  wire                PE40_finish;
  wire       [7:0]    PE41_acount;
  wire       [7:0]    PE41_bcount;
  wire       [31:0]   PE41_PE_OUT;
  wire                PE41_finish;
  wire       [7:0]    PE42_acount;
  wire       [7:0]    PE42_bcount;
  wire       [31:0]   PE42_PE_OUT;
  wire                PE42_finish;
  wire       [7:0]    PE43_acount;
  wire       [7:0]    PE43_bcount;
  wire       [31:0]   PE43_PE_OUT;
  wire                PE43_finish;
  wire       [7:0]    PE44_acount;
  wire       [7:0]    PE44_bcount;
  wire       [31:0]   PE44_PE_OUT;
  wire                PE44_finish;
  wire       [7:0]    PE45_acount;
  wire       [7:0]    PE45_bcount;
  wire       [31:0]   PE45_PE_OUT;
  wire                PE45_finish;
  wire       [7:0]    PE46_acount;
  wire       [7:0]    PE46_bcount;
  wire       [31:0]   PE46_PE_OUT;
  wire                PE46_finish;
  wire       [7:0]    PE47_acount;
  wire       [7:0]    PE47_bcount;
  wire       [31:0]   PE47_PE_OUT;
  wire                PE47_finish;
  wire       [7:0]    PE48_acount;
  wire       [7:0]    PE48_bcount;
  wire       [31:0]   PE48_PE_OUT;
  wire                PE48_finish;
  wire       [7:0]    PE49_acount;
  wire       [7:0]    PE49_bcount;
  wire       [31:0]   PE49_PE_OUT;
  wire                PE49_finish;
  wire       [7:0]    PE410_acount;
  wire       [7:0]    PE410_bcount;
  wire       [31:0]   PE410_PE_OUT;
  wire                PE410_finish;
  wire       [7:0]    PE411_acount;
  wire       [7:0]    PE411_bcount;
  wire       [31:0]   PE411_PE_OUT;
  wire                PE411_finish;
  wire       [7:0]    PE412_acount;
  wire       [7:0]    PE412_bcount;
  wire       [31:0]   PE412_PE_OUT;
  wire                PE412_finish;
  wire       [7:0]    PE413_acount;
  wire       [7:0]    PE413_bcount;
  wire       [31:0]   PE413_PE_OUT;
  wire                PE413_finish;
  wire       [7:0]    PE414_acount;
  wire       [7:0]    PE414_bcount;
  wire       [31:0]   PE414_PE_OUT;
  wire                PE414_finish;
  wire       [7:0]    PE415_acount;
  wire       [7:0]    PE415_bcount;
  wire       [31:0]   PE415_PE_OUT;
  wire                PE415_finish;
  wire       [7:0]    PE416_acount;
  wire       [7:0]    PE416_bcount;
  wire       [31:0]   PE416_PE_OUT;
  wire                PE416_finish;
  wire       [7:0]    PE417_acount;
  wire       [7:0]    PE417_bcount;
  wire       [31:0]   PE417_PE_OUT;
  wire                PE417_finish;
  wire       [7:0]    PE418_acount;
  wire       [7:0]    PE418_bcount;
  wire       [31:0]   PE418_PE_OUT;
  wire                PE418_finish;
  wire       [7:0]    PE419_acount;
  wire       [7:0]    PE419_bcount;
  wire       [31:0]   PE419_PE_OUT;
  wire                PE419_finish;
  wire       [7:0]    PE420_acount;
  wire       [7:0]    PE420_bcount;
  wire       [31:0]   PE420_PE_OUT;
  wire                PE420_finish;
  wire       [7:0]    PE421_acount;
  wire       [7:0]    PE421_bcount;
  wire       [31:0]   PE421_PE_OUT;
  wire                PE421_finish;
  wire       [7:0]    PE422_acount;
  wire       [7:0]    PE422_bcount;
  wire       [31:0]   PE422_PE_OUT;
  wire                PE422_finish;
  wire       [7:0]    PE423_acount;
  wire       [7:0]    PE423_bcount;
  wire       [31:0]   PE423_PE_OUT;
  wire                PE423_finish;
  wire       [7:0]    PE424_acount;
  wire       [7:0]    PE424_bcount;
  wire       [31:0]   PE424_PE_OUT;
  wire                PE424_finish;
  wire       [7:0]    PE425_acount;
  wire       [7:0]    PE425_bcount;
  wire       [31:0]   PE425_PE_OUT;
  wire                PE425_finish;
  wire       [7:0]    PE426_acount;
  wire       [7:0]    PE426_bcount;
  wire       [31:0]   PE426_PE_OUT;
  wire                PE426_finish;
  wire       [7:0]    PE427_acount;
  wire       [7:0]    PE427_bcount;
  wire       [31:0]   PE427_PE_OUT;
  wire                PE427_finish;
  wire       [7:0]    PE428_acount;
  wire       [7:0]    PE428_bcount;
  wire       [31:0]   PE428_PE_OUT;
  wire                PE428_finish;
  wire       [7:0]    PE429_acount;
  wire       [7:0]    PE429_bcount;
  wire       [31:0]   PE429_PE_OUT;
  wire                PE429_finish;
  wire       [7:0]    PE430_acount;
  wire       [7:0]    PE430_bcount;
  wire       [31:0]   PE430_PE_OUT;
  wire                PE430_finish;
  wire       [7:0]    PE431_acount;
  wire       [7:0]    PE431_bcount;
  wire       [31:0]   PE431_PE_OUT;
  wire                PE431_finish;
  wire       [7:0]    PE432_acount;
  wire       [7:0]    PE432_bcount;
  wire       [31:0]   PE432_PE_OUT;
  wire                PE432_finish;
  wire       [7:0]    PE433_acount;
  wire       [7:0]    PE433_bcount;
  wire       [31:0]   PE433_PE_OUT;
  wire                PE433_finish;
  wire       [7:0]    PE434_acount;
  wire       [7:0]    PE434_bcount;
  wire       [31:0]   PE434_PE_OUT;
  wire                PE434_finish;
  wire       [7:0]    PE435_acount;
  wire       [7:0]    PE435_bcount;
  wire       [31:0]   PE435_PE_OUT;
  wire                PE435_finish;
  wire       [7:0]    PE436_acount;
  wire       [7:0]    PE436_bcount;
  wire       [31:0]   PE436_PE_OUT;
  wire                PE436_finish;
  wire       [7:0]    PE437_acount;
  wire       [7:0]    PE437_bcount;
  wire       [31:0]   PE437_PE_OUT;
  wire                PE437_finish;
  wire       [7:0]    PE438_acount;
  wire       [7:0]    PE438_bcount;
  wire       [31:0]   PE438_PE_OUT;
  wire                PE438_finish;
  wire       [7:0]    PE439_acount;
  wire       [7:0]    PE439_bcount;
  wire       [31:0]   PE439_PE_OUT;
  wire                PE439_finish;
  wire       [7:0]    PE440_acount;
  wire       [7:0]    PE440_bcount;
  wire       [31:0]   PE440_PE_OUT;
  wire                PE440_finish;
  wire       [7:0]    PE441_acount;
  wire       [7:0]    PE441_bcount;
  wire       [31:0]   PE441_PE_OUT;
  wire                PE441_finish;
  wire       [7:0]    PE442_acount;
  wire       [7:0]    PE442_bcount;
  wire       [31:0]   PE442_PE_OUT;
  wire                PE442_finish;
  wire       [7:0]    PE443_acount;
  wire       [7:0]    PE443_bcount;
  wire       [31:0]   PE443_PE_OUT;
  wire                PE443_finish;
  wire       [7:0]    PE444_acount;
  wire       [7:0]    PE444_bcount;
  wire       [31:0]   PE444_PE_OUT;
  wire                PE444_finish;
  wire       [7:0]    PE445_acount;
  wire       [7:0]    PE445_bcount;
  wire       [31:0]   PE445_PE_OUT;
  wire                PE445_finish;
  wire       [7:0]    PE446_acount;
  wire       [7:0]    PE446_bcount;
  wire       [31:0]   PE446_PE_OUT;
  wire                PE446_finish;
  wire       [7:0]    PE447_acount;
  wire       [7:0]    PE447_bcount;
  wire       [31:0]   PE447_PE_OUT;
  wire                PE447_finish;
  wire       [7:0]    PE448_acount;
  wire       [7:0]    PE448_bcount;
  wire       [31:0]   PE448_PE_OUT;
  wire                PE448_finish;
  wire       [7:0]    PE449_acount;
  wire       [7:0]    PE449_bcount;
  wire       [31:0]   PE449_PE_OUT;
  wire                PE449_finish;
  wire       [7:0]    PE450_acount;
  wire       [7:0]    PE450_bcount;
  wire       [31:0]   PE450_PE_OUT;
  wire                PE450_finish;
  wire       [7:0]    PE451_acount;
  wire       [7:0]    PE451_bcount;
  wire       [31:0]   PE451_PE_OUT;
  wire                PE451_finish;
  wire       [7:0]    PE452_acount;
  wire       [7:0]    PE452_bcount;
  wire       [31:0]   PE452_PE_OUT;
  wire                PE452_finish;
  wire       [7:0]    PE453_acount;
  wire       [7:0]    PE453_bcount;
  wire       [31:0]   PE453_PE_OUT;
  wire                PE453_finish;
  wire       [7:0]    PE454_acount;
  wire       [7:0]    PE454_bcount;
  wire       [31:0]   PE454_PE_OUT;
  wire                PE454_finish;
  wire       [7:0]    PE455_acount;
  wire       [7:0]    PE455_bcount;
  wire       [31:0]   PE455_PE_OUT;
  wire                PE455_finish;
  wire       [7:0]    PE456_acount;
  wire       [7:0]    PE456_bcount;
  wire       [31:0]   PE456_PE_OUT;
  wire                PE456_finish;
  wire       [7:0]    PE457_acount;
  wire       [7:0]    PE457_bcount;
  wire       [31:0]   PE457_PE_OUT;
  wire                PE457_finish;
  wire       [7:0]    PE458_acount;
  wire       [7:0]    PE458_bcount;
  wire       [31:0]   PE458_PE_OUT;
  wire                PE458_finish;
  wire       [7:0]    PE459_acount;
  wire       [7:0]    PE459_bcount;
  wire       [31:0]   PE459_PE_OUT;
  wire                PE459_finish;
  wire       [7:0]    PE460_acount;
  wire       [7:0]    PE460_bcount;
  wire       [31:0]   PE460_PE_OUT;
  wire                PE460_finish;
  wire       [7:0]    PE461_acount;
  wire       [7:0]    PE461_bcount;
  wire       [31:0]   PE461_PE_OUT;
  wire                PE461_finish;
  wire       [7:0]    PE462_acount;
  wire       [7:0]    PE462_bcount;
  wire       [31:0]   PE462_PE_OUT;
  wire                PE462_finish;
  wire       [7:0]    PE463_acount;
  wire       [7:0]    PE463_bcount;
  wire       [31:0]   PE463_PE_OUT;
  wire                PE463_finish;
  wire       [7:0]    PE50_acount;
  wire       [7:0]    PE50_bcount;
  wire       [31:0]   PE50_PE_OUT;
  wire                PE50_finish;
  wire       [7:0]    PE51_acount;
  wire       [7:0]    PE51_bcount;
  wire       [31:0]   PE51_PE_OUT;
  wire                PE51_finish;
  wire       [7:0]    PE52_acount;
  wire       [7:0]    PE52_bcount;
  wire       [31:0]   PE52_PE_OUT;
  wire                PE52_finish;
  wire       [7:0]    PE53_acount;
  wire       [7:0]    PE53_bcount;
  wire       [31:0]   PE53_PE_OUT;
  wire                PE53_finish;
  wire       [7:0]    PE54_acount;
  wire       [7:0]    PE54_bcount;
  wire       [31:0]   PE54_PE_OUT;
  wire                PE54_finish;
  wire       [7:0]    PE55_acount;
  wire       [7:0]    PE55_bcount;
  wire       [31:0]   PE55_PE_OUT;
  wire                PE55_finish;
  wire       [7:0]    PE56_acount;
  wire       [7:0]    PE56_bcount;
  wire       [31:0]   PE56_PE_OUT;
  wire                PE56_finish;
  wire       [7:0]    PE57_acount;
  wire       [7:0]    PE57_bcount;
  wire       [31:0]   PE57_PE_OUT;
  wire                PE57_finish;
  wire       [7:0]    PE58_acount;
  wire       [7:0]    PE58_bcount;
  wire       [31:0]   PE58_PE_OUT;
  wire                PE58_finish;
  wire       [7:0]    PE59_acount;
  wire       [7:0]    PE59_bcount;
  wire       [31:0]   PE59_PE_OUT;
  wire                PE59_finish;
  wire       [7:0]    PE510_acount;
  wire       [7:0]    PE510_bcount;
  wire       [31:0]   PE510_PE_OUT;
  wire                PE510_finish;
  wire       [7:0]    PE511_acount;
  wire       [7:0]    PE511_bcount;
  wire       [31:0]   PE511_PE_OUT;
  wire                PE511_finish;
  wire       [7:0]    PE512_acount;
  wire       [7:0]    PE512_bcount;
  wire       [31:0]   PE512_PE_OUT;
  wire                PE512_finish;
  wire       [7:0]    PE513_acount;
  wire       [7:0]    PE513_bcount;
  wire       [31:0]   PE513_PE_OUT;
  wire                PE513_finish;
  wire       [7:0]    PE514_acount;
  wire       [7:0]    PE514_bcount;
  wire       [31:0]   PE514_PE_OUT;
  wire                PE514_finish;
  wire       [7:0]    PE515_acount;
  wire       [7:0]    PE515_bcount;
  wire       [31:0]   PE515_PE_OUT;
  wire                PE515_finish;
  wire       [7:0]    PE516_acount;
  wire       [7:0]    PE516_bcount;
  wire       [31:0]   PE516_PE_OUT;
  wire                PE516_finish;
  wire       [7:0]    PE517_acount;
  wire       [7:0]    PE517_bcount;
  wire       [31:0]   PE517_PE_OUT;
  wire                PE517_finish;
  wire       [7:0]    PE518_acount;
  wire       [7:0]    PE518_bcount;
  wire       [31:0]   PE518_PE_OUT;
  wire                PE518_finish;
  wire       [7:0]    PE519_acount;
  wire       [7:0]    PE519_bcount;
  wire       [31:0]   PE519_PE_OUT;
  wire                PE519_finish;
  wire       [7:0]    PE520_acount;
  wire       [7:0]    PE520_bcount;
  wire       [31:0]   PE520_PE_OUT;
  wire                PE520_finish;
  wire       [7:0]    PE521_acount;
  wire       [7:0]    PE521_bcount;
  wire       [31:0]   PE521_PE_OUT;
  wire                PE521_finish;
  wire       [7:0]    PE522_acount;
  wire       [7:0]    PE522_bcount;
  wire       [31:0]   PE522_PE_OUT;
  wire                PE522_finish;
  wire       [7:0]    PE523_acount;
  wire       [7:0]    PE523_bcount;
  wire       [31:0]   PE523_PE_OUT;
  wire                PE523_finish;
  wire       [7:0]    PE524_acount;
  wire       [7:0]    PE524_bcount;
  wire       [31:0]   PE524_PE_OUT;
  wire                PE524_finish;
  wire       [7:0]    PE525_acount;
  wire       [7:0]    PE525_bcount;
  wire       [31:0]   PE525_PE_OUT;
  wire                PE525_finish;
  wire       [7:0]    PE526_acount;
  wire       [7:0]    PE526_bcount;
  wire       [31:0]   PE526_PE_OUT;
  wire                PE526_finish;
  wire       [7:0]    PE527_acount;
  wire       [7:0]    PE527_bcount;
  wire       [31:0]   PE527_PE_OUT;
  wire                PE527_finish;
  wire       [7:0]    PE528_acount;
  wire       [7:0]    PE528_bcount;
  wire       [31:0]   PE528_PE_OUT;
  wire                PE528_finish;
  wire       [7:0]    PE529_acount;
  wire       [7:0]    PE529_bcount;
  wire       [31:0]   PE529_PE_OUT;
  wire                PE529_finish;
  wire       [7:0]    PE530_acount;
  wire       [7:0]    PE530_bcount;
  wire       [31:0]   PE530_PE_OUT;
  wire                PE530_finish;
  wire       [7:0]    PE531_acount;
  wire       [7:0]    PE531_bcount;
  wire       [31:0]   PE531_PE_OUT;
  wire                PE531_finish;
  wire       [7:0]    PE532_acount;
  wire       [7:0]    PE532_bcount;
  wire       [31:0]   PE532_PE_OUT;
  wire                PE532_finish;
  wire       [7:0]    PE533_acount;
  wire       [7:0]    PE533_bcount;
  wire       [31:0]   PE533_PE_OUT;
  wire                PE533_finish;
  wire       [7:0]    PE534_acount;
  wire       [7:0]    PE534_bcount;
  wire       [31:0]   PE534_PE_OUT;
  wire                PE534_finish;
  wire       [7:0]    PE535_acount;
  wire       [7:0]    PE535_bcount;
  wire       [31:0]   PE535_PE_OUT;
  wire                PE535_finish;
  wire       [7:0]    PE536_acount;
  wire       [7:0]    PE536_bcount;
  wire       [31:0]   PE536_PE_OUT;
  wire                PE536_finish;
  wire       [7:0]    PE537_acount;
  wire       [7:0]    PE537_bcount;
  wire       [31:0]   PE537_PE_OUT;
  wire                PE537_finish;
  wire       [7:0]    PE538_acount;
  wire       [7:0]    PE538_bcount;
  wire       [31:0]   PE538_PE_OUT;
  wire                PE538_finish;
  wire       [7:0]    PE539_acount;
  wire       [7:0]    PE539_bcount;
  wire       [31:0]   PE539_PE_OUT;
  wire                PE539_finish;
  wire       [7:0]    PE540_acount;
  wire       [7:0]    PE540_bcount;
  wire       [31:0]   PE540_PE_OUT;
  wire                PE540_finish;
  wire       [7:0]    PE541_acount;
  wire       [7:0]    PE541_bcount;
  wire       [31:0]   PE541_PE_OUT;
  wire                PE541_finish;
  wire       [7:0]    PE542_acount;
  wire       [7:0]    PE542_bcount;
  wire       [31:0]   PE542_PE_OUT;
  wire                PE542_finish;
  wire       [7:0]    PE543_acount;
  wire       [7:0]    PE543_bcount;
  wire       [31:0]   PE543_PE_OUT;
  wire                PE543_finish;
  wire       [7:0]    PE544_acount;
  wire       [7:0]    PE544_bcount;
  wire       [31:0]   PE544_PE_OUT;
  wire                PE544_finish;
  wire       [7:0]    PE545_acount;
  wire       [7:0]    PE545_bcount;
  wire       [31:0]   PE545_PE_OUT;
  wire                PE545_finish;
  wire       [7:0]    PE546_acount;
  wire       [7:0]    PE546_bcount;
  wire       [31:0]   PE546_PE_OUT;
  wire                PE546_finish;
  wire       [7:0]    PE547_acount;
  wire       [7:0]    PE547_bcount;
  wire       [31:0]   PE547_PE_OUT;
  wire                PE547_finish;
  wire       [7:0]    PE548_acount;
  wire       [7:0]    PE548_bcount;
  wire       [31:0]   PE548_PE_OUT;
  wire                PE548_finish;
  wire       [7:0]    PE549_acount;
  wire       [7:0]    PE549_bcount;
  wire       [31:0]   PE549_PE_OUT;
  wire                PE549_finish;
  wire       [7:0]    PE550_acount;
  wire       [7:0]    PE550_bcount;
  wire       [31:0]   PE550_PE_OUT;
  wire                PE550_finish;
  wire       [7:0]    PE551_acount;
  wire       [7:0]    PE551_bcount;
  wire       [31:0]   PE551_PE_OUT;
  wire                PE551_finish;
  wire       [7:0]    PE552_acount;
  wire       [7:0]    PE552_bcount;
  wire       [31:0]   PE552_PE_OUT;
  wire                PE552_finish;
  wire       [7:0]    PE553_acount;
  wire       [7:0]    PE553_bcount;
  wire       [31:0]   PE553_PE_OUT;
  wire                PE553_finish;
  wire       [7:0]    PE554_acount;
  wire       [7:0]    PE554_bcount;
  wire       [31:0]   PE554_PE_OUT;
  wire                PE554_finish;
  wire       [7:0]    PE555_acount;
  wire       [7:0]    PE555_bcount;
  wire       [31:0]   PE555_PE_OUT;
  wire                PE555_finish;
  wire       [7:0]    PE556_acount;
  wire       [7:0]    PE556_bcount;
  wire       [31:0]   PE556_PE_OUT;
  wire                PE556_finish;
  wire       [7:0]    PE557_acount;
  wire       [7:0]    PE557_bcount;
  wire       [31:0]   PE557_PE_OUT;
  wire                PE557_finish;
  wire       [7:0]    PE558_acount;
  wire       [7:0]    PE558_bcount;
  wire       [31:0]   PE558_PE_OUT;
  wire                PE558_finish;
  wire       [7:0]    PE559_acount;
  wire       [7:0]    PE559_bcount;
  wire       [31:0]   PE559_PE_OUT;
  wire                PE559_finish;
  wire       [7:0]    PE560_acount;
  wire       [7:0]    PE560_bcount;
  wire       [31:0]   PE560_PE_OUT;
  wire                PE560_finish;
  wire       [7:0]    PE561_acount;
  wire       [7:0]    PE561_bcount;
  wire       [31:0]   PE561_PE_OUT;
  wire                PE561_finish;
  wire       [7:0]    PE562_acount;
  wire       [7:0]    PE562_bcount;
  wire       [31:0]   PE562_PE_OUT;
  wire                PE562_finish;
  wire       [7:0]    PE563_acount;
  wire       [7:0]    PE563_bcount;
  wire       [31:0]   PE563_PE_OUT;
  wire                PE563_finish;
  wire       [7:0]    PE60_acount;
  wire       [7:0]    PE60_bcount;
  wire       [31:0]   PE60_PE_OUT;
  wire                PE60_finish;
  wire       [7:0]    PE61_acount;
  wire       [7:0]    PE61_bcount;
  wire       [31:0]   PE61_PE_OUT;
  wire                PE61_finish;
  wire       [7:0]    PE62_acount;
  wire       [7:0]    PE62_bcount;
  wire       [31:0]   PE62_PE_OUT;
  wire                PE62_finish;
  wire       [7:0]    PE63_acount;
  wire       [7:0]    PE63_bcount;
  wire       [31:0]   PE63_PE_OUT;
  wire                PE63_finish;
  wire       [7:0]    PE64_acount;
  wire       [7:0]    PE64_bcount;
  wire       [31:0]   PE64_PE_OUT;
  wire                PE64_finish;
  wire       [7:0]    PE65_acount;
  wire       [7:0]    PE65_bcount;
  wire       [31:0]   PE65_PE_OUT;
  wire                PE65_finish;
  wire       [7:0]    PE66_acount;
  wire       [7:0]    PE66_bcount;
  wire       [31:0]   PE66_PE_OUT;
  wire                PE66_finish;
  wire       [7:0]    PE67_acount;
  wire       [7:0]    PE67_bcount;
  wire       [31:0]   PE67_PE_OUT;
  wire                PE67_finish;
  wire       [7:0]    PE68_acount;
  wire       [7:0]    PE68_bcount;
  wire       [31:0]   PE68_PE_OUT;
  wire                PE68_finish;
  wire       [7:0]    PE69_acount;
  wire       [7:0]    PE69_bcount;
  wire       [31:0]   PE69_PE_OUT;
  wire                PE69_finish;
  wire       [7:0]    PE610_acount;
  wire       [7:0]    PE610_bcount;
  wire       [31:0]   PE610_PE_OUT;
  wire                PE610_finish;
  wire       [7:0]    PE611_acount;
  wire       [7:0]    PE611_bcount;
  wire       [31:0]   PE611_PE_OUT;
  wire                PE611_finish;
  wire       [7:0]    PE612_acount;
  wire       [7:0]    PE612_bcount;
  wire       [31:0]   PE612_PE_OUT;
  wire                PE612_finish;
  wire       [7:0]    PE613_acount;
  wire       [7:0]    PE613_bcount;
  wire       [31:0]   PE613_PE_OUT;
  wire                PE613_finish;
  wire       [7:0]    PE614_acount;
  wire       [7:0]    PE614_bcount;
  wire       [31:0]   PE614_PE_OUT;
  wire                PE614_finish;
  wire       [7:0]    PE615_acount;
  wire       [7:0]    PE615_bcount;
  wire       [31:0]   PE615_PE_OUT;
  wire                PE615_finish;
  wire       [7:0]    PE616_acount;
  wire       [7:0]    PE616_bcount;
  wire       [31:0]   PE616_PE_OUT;
  wire                PE616_finish;
  wire       [7:0]    PE617_acount;
  wire       [7:0]    PE617_bcount;
  wire       [31:0]   PE617_PE_OUT;
  wire                PE617_finish;
  wire       [7:0]    PE618_acount;
  wire       [7:0]    PE618_bcount;
  wire       [31:0]   PE618_PE_OUT;
  wire                PE618_finish;
  wire       [7:0]    PE619_acount;
  wire       [7:0]    PE619_bcount;
  wire       [31:0]   PE619_PE_OUT;
  wire                PE619_finish;
  wire       [7:0]    PE620_acount;
  wire       [7:0]    PE620_bcount;
  wire       [31:0]   PE620_PE_OUT;
  wire                PE620_finish;
  wire       [7:0]    PE621_acount;
  wire       [7:0]    PE621_bcount;
  wire       [31:0]   PE621_PE_OUT;
  wire                PE621_finish;
  wire       [7:0]    PE622_acount;
  wire       [7:0]    PE622_bcount;
  wire       [31:0]   PE622_PE_OUT;
  wire                PE622_finish;
  wire       [7:0]    PE623_acount;
  wire       [7:0]    PE623_bcount;
  wire       [31:0]   PE623_PE_OUT;
  wire                PE623_finish;
  wire       [7:0]    PE624_acount;
  wire       [7:0]    PE624_bcount;
  wire       [31:0]   PE624_PE_OUT;
  wire                PE624_finish;
  wire       [7:0]    PE625_acount;
  wire       [7:0]    PE625_bcount;
  wire       [31:0]   PE625_PE_OUT;
  wire                PE625_finish;
  wire       [7:0]    PE626_acount;
  wire       [7:0]    PE626_bcount;
  wire       [31:0]   PE626_PE_OUT;
  wire                PE626_finish;
  wire       [7:0]    PE627_acount;
  wire       [7:0]    PE627_bcount;
  wire       [31:0]   PE627_PE_OUT;
  wire                PE627_finish;
  wire       [7:0]    PE628_acount;
  wire       [7:0]    PE628_bcount;
  wire       [31:0]   PE628_PE_OUT;
  wire                PE628_finish;
  wire       [7:0]    PE629_acount;
  wire       [7:0]    PE629_bcount;
  wire       [31:0]   PE629_PE_OUT;
  wire                PE629_finish;
  wire       [7:0]    PE630_acount;
  wire       [7:0]    PE630_bcount;
  wire       [31:0]   PE630_PE_OUT;
  wire                PE630_finish;
  wire       [7:0]    PE631_acount;
  wire       [7:0]    PE631_bcount;
  wire       [31:0]   PE631_PE_OUT;
  wire                PE631_finish;
  wire       [7:0]    PE632_acount;
  wire       [7:0]    PE632_bcount;
  wire       [31:0]   PE632_PE_OUT;
  wire                PE632_finish;
  wire       [7:0]    PE633_acount;
  wire       [7:0]    PE633_bcount;
  wire       [31:0]   PE633_PE_OUT;
  wire                PE633_finish;
  wire       [7:0]    PE634_acount;
  wire       [7:0]    PE634_bcount;
  wire       [31:0]   PE634_PE_OUT;
  wire                PE634_finish;
  wire       [7:0]    PE635_acount;
  wire       [7:0]    PE635_bcount;
  wire       [31:0]   PE635_PE_OUT;
  wire                PE635_finish;
  wire       [7:0]    PE636_acount;
  wire       [7:0]    PE636_bcount;
  wire       [31:0]   PE636_PE_OUT;
  wire                PE636_finish;
  wire       [7:0]    PE637_acount;
  wire       [7:0]    PE637_bcount;
  wire       [31:0]   PE637_PE_OUT;
  wire                PE637_finish;
  wire       [7:0]    PE638_acount;
  wire       [7:0]    PE638_bcount;
  wire       [31:0]   PE638_PE_OUT;
  wire                PE638_finish;
  wire       [7:0]    PE639_acount;
  wire       [7:0]    PE639_bcount;
  wire       [31:0]   PE639_PE_OUT;
  wire                PE639_finish;
  wire       [7:0]    PE640_acount;
  wire       [7:0]    PE640_bcount;
  wire       [31:0]   PE640_PE_OUT;
  wire                PE640_finish;
  wire       [7:0]    PE641_acount;
  wire       [7:0]    PE641_bcount;
  wire       [31:0]   PE641_PE_OUT;
  wire                PE641_finish;
  wire       [7:0]    PE642_acount;
  wire       [7:0]    PE642_bcount;
  wire       [31:0]   PE642_PE_OUT;
  wire                PE642_finish;
  wire       [7:0]    PE643_acount;
  wire       [7:0]    PE643_bcount;
  wire       [31:0]   PE643_PE_OUT;
  wire                PE643_finish;
  wire       [7:0]    PE644_acount;
  wire       [7:0]    PE644_bcount;
  wire       [31:0]   PE644_PE_OUT;
  wire                PE644_finish;
  wire       [7:0]    PE645_acount;
  wire       [7:0]    PE645_bcount;
  wire       [31:0]   PE645_PE_OUT;
  wire                PE645_finish;
  wire       [7:0]    PE646_acount;
  wire       [7:0]    PE646_bcount;
  wire       [31:0]   PE646_PE_OUT;
  wire                PE646_finish;
  wire       [7:0]    PE647_acount;
  wire       [7:0]    PE647_bcount;
  wire       [31:0]   PE647_PE_OUT;
  wire                PE647_finish;
  wire       [7:0]    PE648_acount;
  wire       [7:0]    PE648_bcount;
  wire       [31:0]   PE648_PE_OUT;
  wire                PE648_finish;
  wire       [7:0]    PE649_acount;
  wire       [7:0]    PE649_bcount;
  wire       [31:0]   PE649_PE_OUT;
  wire                PE649_finish;
  wire       [7:0]    PE650_acount;
  wire       [7:0]    PE650_bcount;
  wire       [31:0]   PE650_PE_OUT;
  wire                PE650_finish;
  wire       [7:0]    PE651_acount;
  wire       [7:0]    PE651_bcount;
  wire       [31:0]   PE651_PE_OUT;
  wire                PE651_finish;
  wire       [7:0]    PE652_acount;
  wire       [7:0]    PE652_bcount;
  wire       [31:0]   PE652_PE_OUT;
  wire                PE652_finish;
  wire       [7:0]    PE653_acount;
  wire       [7:0]    PE653_bcount;
  wire       [31:0]   PE653_PE_OUT;
  wire                PE653_finish;
  wire       [7:0]    PE654_acount;
  wire       [7:0]    PE654_bcount;
  wire       [31:0]   PE654_PE_OUT;
  wire                PE654_finish;
  wire       [7:0]    PE655_acount;
  wire       [7:0]    PE655_bcount;
  wire       [31:0]   PE655_PE_OUT;
  wire                PE655_finish;
  wire       [7:0]    PE656_acount;
  wire       [7:0]    PE656_bcount;
  wire       [31:0]   PE656_PE_OUT;
  wire                PE656_finish;
  wire       [7:0]    PE657_acount;
  wire       [7:0]    PE657_bcount;
  wire       [31:0]   PE657_PE_OUT;
  wire                PE657_finish;
  wire       [7:0]    PE658_acount;
  wire       [7:0]    PE658_bcount;
  wire       [31:0]   PE658_PE_OUT;
  wire                PE658_finish;
  wire       [7:0]    PE659_acount;
  wire       [7:0]    PE659_bcount;
  wire       [31:0]   PE659_PE_OUT;
  wire                PE659_finish;
  wire       [7:0]    PE660_acount;
  wire       [7:0]    PE660_bcount;
  wire       [31:0]   PE660_PE_OUT;
  wire                PE660_finish;
  wire       [7:0]    PE661_acount;
  wire       [7:0]    PE661_bcount;
  wire       [31:0]   PE661_PE_OUT;
  wire                PE661_finish;
  wire       [7:0]    PE662_acount;
  wire       [7:0]    PE662_bcount;
  wire       [31:0]   PE662_PE_OUT;
  wire                PE662_finish;
  wire       [7:0]    PE663_acount;
  wire       [7:0]    PE663_bcount;
  wire       [31:0]   PE663_PE_OUT;
  wire                PE663_finish;
  wire       [7:0]    PE70_acount;
  wire       [7:0]    PE70_bcount;
  wire       [31:0]   PE70_PE_OUT;
  wire                PE70_finish;
  wire       [7:0]    PE71_acount;
  wire       [7:0]    PE71_bcount;
  wire       [31:0]   PE71_PE_OUT;
  wire                PE71_finish;
  wire       [7:0]    PE72_acount;
  wire       [7:0]    PE72_bcount;
  wire       [31:0]   PE72_PE_OUT;
  wire                PE72_finish;
  wire       [7:0]    PE73_acount;
  wire       [7:0]    PE73_bcount;
  wire       [31:0]   PE73_PE_OUT;
  wire                PE73_finish;
  wire       [7:0]    PE74_acount;
  wire       [7:0]    PE74_bcount;
  wire       [31:0]   PE74_PE_OUT;
  wire                PE74_finish;
  wire       [7:0]    PE75_acount;
  wire       [7:0]    PE75_bcount;
  wire       [31:0]   PE75_PE_OUT;
  wire                PE75_finish;
  wire       [7:0]    PE76_acount;
  wire       [7:0]    PE76_bcount;
  wire       [31:0]   PE76_PE_OUT;
  wire                PE76_finish;
  wire       [7:0]    PE77_acount;
  wire       [7:0]    PE77_bcount;
  wire       [31:0]   PE77_PE_OUT;
  wire                PE77_finish;
  wire       [7:0]    PE78_acount;
  wire       [7:0]    PE78_bcount;
  wire       [31:0]   PE78_PE_OUT;
  wire                PE78_finish;
  wire       [7:0]    PE79_acount;
  wire       [7:0]    PE79_bcount;
  wire       [31:0]   PE79_PE_OUT;
  wire                PE79_finish;
  wire       [7:0]    PE710_acount;
  wire       [7:0]    PE710_bcount;
  wire       [31:0]   PE710_PE_OUT;
  wire                PE710_finish;
  wire       [7:0]    PE711_acount;
  wire       [7:0]    PE711_bcount;
  wire       [31:0]   PE711_PE_OUT;
  wire                PE711_finish;
  wire       [7:0]    PE712_acount;
  wire       [7:0]    PE712_bcount;
  wire       [31:0]   PE712_PE_OUT;
  wire                PE712_finish;
  wire       [7:0]    PE713_acount;
  wire       [7:0]    PE713_bcount;
  wire       [31:0]   PE713_PE_OUT;
  wire                PE713_finish;
  wire       [7:0]    PE714_acount;
  wire       [7:0]    PE714_bcount;
  wire       [31:0]   PE714_PE_OUT;
  wire                PE714_finish;
  wire       [7:0]    PE715_acount;
  wire       [7:0]    PE715_bcount;
  wire       [31:0]   PE715_PE_OUT;
  wire                PE715_finish;
  wire       [7:0]    PE716_acount;
  wire       [7:0]    PE716_bcount;
  wire       [31:0]   PE716_PE_OUT;
  wire                PE716_finish;
  wire       [7:0]    PE717_acount;
  wire       [7:0]    PE717_bcount;
  wire       [31:0]   PE717_PE_OUT;
  wire                PE717_finish;
  wire       [7:0]    PE718_acount;
  wire       [7:0]    PE718_bcount;
  wire       [31:0]   PE718_PE_OUT;
  wire                PE718_finish;
  wire       [7:0]    PE719_acount;
  wire       [7:0]    PE719_bcount;
  wire       [31:0]   PE719_PE_OUT;
  wire                PE719_finish;
  wire       [7:0]    PE720_acount;
  wire       [7:0]    PE720_bcount;
  wire       [31:0]   PE720_PE_OUT;
  wire                PE720_finish;
  wire       [7:0]    PE721_acount;
  wire       [7:0]    PE721_bcount;
  wire       [31:0]   PE721_PE_OUT;
  wire                PE721_finish;
  wire       [7:0]    PE722_acount;
  wire       [7:0]    PE722_bcount;
  wire       [31:0]   PE722_PE_OUT;
  wire                PE722_finish;
  wire       [7:0]    PE723_acount;
  wire       [7:0]    PE723_bcount;
  wire       [31:0]   PE723_PE_OUT;
  wire                PE723_finish;
  wire       [7:0]    PE724_acount;
  wire       [7:0]    PE724_bcount;
  wire       [31:0]   PE724_PE_OUT;
  wire                PE724_finish;
  wire       [7:0]    PE725_acount;
  wire       [7:0]    PE725_bcount;
  wire       [31:0]   PE725_PE_OUT;
  wire                PE725_finish;
  wire       [7:0]    PE726_acount;
  wire       [7:0]    PE726_bcount;
  wire       [31:0]   PE726_PE_OUT;
  wire                PE726_finish;
  wire       [7:0]    PE727_acount;
  wire       [7:0]    PE727_bcount;
  wire       [31:0]   PE727_PE_OUT;
  wire                PE727_finish;
  wire       [7:0]    PE728_acount;
  wire       [7:0]    PE728_bcount;
  wire       [31:0]   PE728_PE_OUT;
  wire                PE728_finish;
  wire       [7:0]    PE729_acount;
  wire       [7:0]    PE729_bcount;
  wire       [31:0]   PE729_PE_OUT;
  wire                PE729_finish;
  wire       [7:0]    PE730_acount;
  wire       [7:0]    PE730_bcount;
  wire       [31:0]   PE730_PE_OUT;
  wire                PE730_finish;
  wire       [7:0]    PE731_acount;
  wire       [7:0]    PE731_bcount;
  wire       [31:0]   PE731_PE_OUT;
  wire                PE731_finish;
  wire       [7:0]    PE732_acount;
  wire       [7:0]    PE732_bcount;
  wire       [31:0]   PE732_PE_OUT;
  wire                PE732_finish;
  wire       [7:0]    PE733_acount;
  wire       [7:0]    PE733_bcount;
  wire       [31:0]   PE733_PE_OUT;
  wire                PE733_finish;
  wire       [7:0]    PE734_acount;
  wire       [7:0]    PE734_bcount;
  wire       [31:0]   PE734_PE_OUT;
  wire                PE734_finish;
  wire       [7:0]    PE735_acount;
  wire       [7:0]    PE735_bcount;
  wire       [31:0]   PE735_PE_OUT;
  wire                PE735_finish;
  wire       [7:0]    PE736_acount;
  wire       [7:0]    PE736_bcount;
  wire       [31:0]   PE736_PE_OUT;
  wire                PE736_finish;
  wire       [7:0]    PE737_acount;
  wire       [7:0]    PE737_bcount;
  wire       [31:0]   PE737_PE_OUT;
  wire                PE737_finish;
  wire       [7:0]    PE738_acount;
  wire       [7:0]    PE738_bcount;
  wire       [31:0]   PE738_PE_OUT;
  wire                PE738_finish;
  wire       [7:0]    PE739_acount;
  wire       [7:0]    PE739_bcount;
  wire       [31:0]   PE739_PE_OUT;
  wire                PE739_finish;
  wire       [7:0]    PE740_acount;
  wire       [7:0]    PE740_bcount;
  wire       [31:0]   PE740_PE_OUT;
  wire                PE740_finish;
  wire       [7:0]    PE741_acount;
  wire       [7:0]    PE741_bcount;
  wire       [31:0]   PE741_PE_OUT;
  wire                PE741_finish;
  wire       [7:0]    PE742_acount;
  wire       [7:0]    PE742_bcount;
  wire       [31:0]   PE742_PE_OUT;
  wire                PE742_finish;
  wire       [7:0]    PE743_acount;
  wire       [7:0]    PE743_bcount;
  wire       [31:0]   PE743_PE_OUT;
  wire                PE743_finish;
  wire       [7:0]    PE744_acount;
  wire       [7:0]    PE744_bcount;
  wire       [31:0]   PE744_PE_OUT;
  wire                PE744_finish;
  wire       [7:0]    PE745_acount;
  wire       [7:0]    PE745_bcount;
  wire       [31:0]   PE745_PE_OUT;
  wire                PE745_finish;
  wire       [7:0]    PE746_acount;
  wire       [7:0]    PE746_bcount;
  wire       [31:0]   PE746_PE_OUT;
  wire                PE746_finish;
  wire       [7:0]    PE747_acount;
  wire       [7:0]    PE747_bcount;
  wire       [31:0]   PE747_PE_OUT;
  wire                PE747_finish;
  wire       [7:0]    PE748_acount;
  wire       [7:0]    PE748_bcount;
  wire       [31:0]   PE748_PE_OUT;
  wire                PE748_finish;
  wire       [7:0]    PE749_acount;
  wire       [7:0]    PE749_bcount;
  wire       [31:0]   PE749_PE_OUT;
  wire                PE749_finish;
  wire       [7:0]    PE750_acount;
  wire       [7:0]    PE750_bcount;
  wire       [31:0]   PE750_PE_OUT;
  wire                PE750_finish;
  wire       [7:0]    PE751_acount;
  wire       [7:0]    PE751_bcount;
  wire       [31:0]   PE751_PE_OUT;
  wire                PE751_finish;
  wire       [7:0]    PE752_acount;
  wire       [7:0]    PE752_bcount;
  wire       [31:0]   PE752_PE_OUT;
  wire                PE752_finish;
  wire       [7:0]    PE753_acount;
  wire       [7:0]    PE753_bcount;
  wire       [31:0]   PE753_PE_OUT;
  wire                PE753_finish;
  wire       [7:0]    PE754_acount;
  wire       [7:0]    PE754_bcount;
  wire       [31:0]   PE754_PE_OUT;
  wire                PE754_finish;
  wire       [7:0]    PE755_acount;
  wire       [7:0]    PE755_bcount;
  wire       [31:0]   PE755_PE_OUT;
  wire                PE755_finish;
  wire       [7:0]    PE756_acount;
  wire       [7:0]    PE756_bcount;
  wire       [31:0]   PE756_PE_OUT;
  wire                PE756_finish;
  wire       [7:0]    PE757_acount;
  wire       [7:0]    PE757_bcount;
  wire       [31:0]   PE757_PE_OUT;
  wire                PE757_finish;
  wire       [7:0]    PE758_acount;
  wire       [7:0]    PE758_bcount;
  wire       [31:0]   PE758_PE_OUT;
  wire                PE758_finish;
  wire       [7:0]    PE759_acount;
  wire       [7:0]    PE759_bcount;
  wire       [31:0]   PE759_PE_OUT;
  wire                PE759_finish;
  wire       [7:0]    PE760_acount;
  wire       [7:0]    PE760_bcount;
  wire       [31:0]   PE760_PE_OUT;
  wire                PE760_finish;
  wire       [7:0]    PE761_acount;
  wire       [7:0]    PE761_bcount;
  wire       [31:0]   PE761_PE_OUT;
  wire                PE761_finish;
  wire       [7:0]    PE762_acount;
  wire       [7:0]    PE762_bcount;
  wire       [31:0]   PE762_PE_OUT;
  wire                PE762_finish;
  wire       [7:0]    PE763_acount;
  wire       [7:0]    PE763_bcount;
  wire       [31:0]   PE763_PE_OUT;
  wire                PE763_finish;
  reg        [63:0]   _zz_C_Valid_0;
  reg        [63:0]   _zz_C_Valid_1;
  reg        [63:0]   _zz_C_Valid_2;
  reg        [63:0]   _zz_C_Valid_3;
  reg        [63:0]   _zz_C_Valid_4;
  reg        [63:0]   _zz_C_Valid_5;
  reg        [63:0]   _zz_C_Valid_6;
  reg        [63:0]   _zz_C_Valid_7;
  reg        [15:0]   io_signCount_regNextWhen;
  reg                 io_A_Valid_0_delay_1;
  reg                 io_A_Valid_0_delay_1_1;
  reg                 io_A_Valid_0_delay_2;
  reg                 io_A_Valid_0_delay_1_2;
  reg                 io_A_Valid_0_delay_2_1;
  reg                 io_A_Valid_0_delay_3;
  reg                 io_A_Valid_0_delay_1_3;
  reg                 io_A_Valid_0_delay_2_2;
  reg                 io_A_Valid_0_delay_3_1;
  reg                 io_A_Valid_0_delay_4;
  reg                 io_A_Valid_0_delay_1_4;
  reg                 io_A_Valid_0_delay_2_3;
  reg                 io_A_Valid_0_delay_3_2;
  reg                 io_A_Valid_0_delay_4_1;
  reg                 io_A_Valid_0_delay_5;
  reg                 io_A_Valid_0_delay_1_5;
  reg                 io_A_Valid_0_delay_2_4;
  reg                 io_A_Valid_0_delay_3_3;
  reg                 io_A_Valid_0_delay_4_2;
  reg                 io_A_Valid_0_delay_5_1;
  reg                 io_A_Valid_0_delay_6;
  reg                 io_A_Valid_0_delay_1_6;
  reg                 io_A_Valid_0_delay_2_5;
  reg                 io_A_Valid_0_delay_3_4;
  reg                 io_A_Valid_0_delay_4_3;
  reg                 io_A_Valid_0_delay_5_2;
  reg                 io_A_Valid_0_delay_6_1;
  reg                 io_A_Valid_0_delay_7;
  reg                 io_A_Valid_0_delay_1_7;
  reg                 io_A_Valid_0_delay_2_6;
  reg                 io_A_Valid_0_delay_3_5;
  reg                 io_A_Valid_0_delay_4_4;
  reg                 io_A_Valid_0_delay_5_3;
  reg                 io_A_Valid_0_delay_6_2;
  reg                 io_A_Valid_0_delay_7_1;
  reg                 io_A_Valid_0_delay_8;
  reg                 io_A_Valid_0_delay_1_8;
  reg                 io_A_Valid_0_delay_2_7;
  reg                 io_A_Valid_0_delay_3_6;
  reg                 io_A_Valid_0_delay_4_5;
  reg                 io_A_Valid_0_delay_5_4;
  reg                 io_A_Valid_0_delay_6_3;
  reg                 io_A_Valid_0_delay_7_2;
  reg                 io_A_Valid_0_delay_8_1;
  reg                 io_A_Valid_0_delay_9;
  reg                 io_A_Valid_0_delay_1_9;
  reg                 io_A_Valid_0_delay_2_8;
  reg                 io_A_Valid_0_delay_3_7;
  reg                 io_A_Valid_0_delay_4_6;
  reg                 io_A_Valid_0_delay_5_5;
  reg                 io_A_Valid_0_delay_6_4;
  reg                 io_A_Valid_0_delay_7_3;
  reg                 io_A_Valid_0_delay_8_2;
  reg                 io_A_Valid_0_delay_9_1;
  reg                 io_A_Valid_0_delay_10;
  reg                 io_A_Valid_0_delay_1_10;
  reg                 io_A_Valid_0_delay_2_9;
  reg                 io_A_Valid_0_delay_3_8;
  reg                 io_A_Valid_0_delay_4_7;
  reg                 io_A_Valid_0_delay_5_6;
  reg                 io_A_Valid_0_delay_6_5;
  reg                 io_A_Valid_0_delay_7_4;
  reg                 io_A_Valid_0_delay_8_3;
  reg                 io_A_Valid_0_delay_9_2;
  reg                 io_A_Valid_0_delay_10_1;
  reg                 io_A_Valid_0_delay_11;
  reg                 io_A_Valid_0_delay_1_11;
  reg                 io_A_Valid_0_delay_2_10;
  reg                 io_A_Valid_0_delay_3_9;
  reg                 io_A_Valid_0_delay_4_8;
  reg                 io_A_Valid_0_delay_5_7;
  reg                 io_A_Valid_0_delay_6_6;
  reg                 io_A_Valid_0_delay_7_5;
  reg                 io_A_Valid_0_delay_8_4;
  reg                 io_A_Valid_0_delay_9_3;
  reg                 io_A_Valid_0_delay_10_2;
  reg                 io_A_Valid_0_delay_11_1;
  reg                 io_A_Valid_0_delay_12;
  reg                 io_A_Valid_0_delay_1_12;
  reg                 io_A_Valid_0_delay_2_11;
  reg                 io_A_Valid_0_delay_3_10;
  reg                 io_A_Valid_0_delay_4_9;
  reg                 io_A_Valid_0_delay_5_8;
  reg                 io_A_Valid_0_delay_6_7;
  reg                 io_A_Valid_0_delay_7_6;
  reg                 io_A_Valid_0_delay_8_5;
  reg                 io_A_Valid_0_delay_9_4;
  reg                 io_A_Valid_0_delay_10_3;
  reg                 io_A_Valid_0_delay_11_2;
  reg                 io_A_Valid_0_delay_12_1;
  reg                 io_A_Valid_0_delay_13;
  reg                 io_A_Valid_0_delay_1_13;
  reg                 io_A_Valid_0_delay_2_12;
  reg                 io_A_Valid_0_delay_3_11;
  reg                 io_A_Valid_0_delay_4_10;
  reg                 io_A_Valid_0_delay_5_9;
  reg                 io_A_Valid_0_delay_6_8;
  reg                 io_A_Valid_0_delay_7_7;
  reg                 io_A_Valid_0_delay_8_6;
  reg                 io_A_Valid_0_delay_9_5;
  reg                 io_A_Valid_0_delay_10_4;
  reg                 io_A_Valid_0_delay_11_3;
  reg                 io_A_Valid_0_delay_12_2;
  reg                 io_A_Valid_0_delay_13_1;
  reg                 io_A_Valid_0_delay_14;
  reg                 io_A_Valid_0_delay_1_14;
  reg                 io_A_Valid_0_delay_2_13;
  reg                 io_A_Valid_0_delay_3_12;
  reg                 io_A_Valid_0_delay_4_11;
  reg                 io_A_Valid_0_delay_5_10;
  reg                 io_A_Valid_0_delay_6_9;
  reg                 io_A_Valid_0_delay_7_8;
  reg                 io_A_Valid_0_delay_8_7;
  reg                 io_A_Valid_0_delay_9_6;
  reg                 io_A_Valid_0_delay_10_5;
  reg                 io_A_Valid_0_delay_11_4;
  reg                 io_A_Valid_0_delay_12_3;
  reg                 io_A_Valid_0_delay_13_2;
  reg                 io_A_Valid_0_delay_14_1;
  reg                 io_A_Valid_0_delay_15;
  reg                 io_A_Valid_0_delay_1_15;
  reg                 io_A_Valid_0_delay_2_14;
  reg                 io_A_Valid_0_delay_3_13;
  reg                 io_A_Valid_0_delay_4_12;
  reg                 io_A_Valid_0_delay_5_11;
  reg                 io_A_Valid_0_delay_6_10;
  reg                 io_A_Valid_0_delay_7_9;
  reg                 io_A_Valid_0_delay_8_8;
  reg                 io_A_Valid_0_delay_9_7;
  reg                 io_A_Valid_0_delay_10_6;
  reg                 io_A_Valid_0_delay_11_5;
  reg                 io_A_Valid_0_delay_12_4;
  reg                 io_A_Valid_0_delay_13_3;
  reg                 io_A_Valid_0_delay_14_2;
  reg                 io_A_Valid_0_delay_15_1;
  reg                 io_A_Valid_0_delay_16;
  reg                 io_A_Valid_0_delay_1_16;
  reg                 io_A_Valid_0_delay_2_15;
  reg                 io_A_Valid_0_delay_3_14;
  reg                 io_A_Valid_0_delay_4_13;
  reg                 io_A_Valid_0_delay_5_12;
  reg                 io_A_Valid_0_delay_6_11;
  reg                 io_A_Valid_0_delay_7_10;
  reg                 io_A_Valid_0_delay_8_9;
  reg                 io_A_Valid_0_delay_9_8;
  reg                 io_A_Valid_0_delay_10_7;
  reg                 io_A_Valid_0_delay_11_6;
  reg                 io_A_Valid_0_delay_12_5;
  reg                 io_A_Valid_0_delay_13_4;
  reg                 io_A_Valid_0_delay_14_3;
  reg                 io_A_Valid_0_delay_15_2;
  reg                 io_A_Valid_0_delay_16_1;
  reg                 io_A_Valid_0_delay_17;
  reg                 io_A_Valid_0_delay_1_17;
  reg                 io_A_Valid_0_delay_2_16;
  reg                 io_A_Valid_0_delay_3_15;
  reg                 io_A_Valid_0_delay_4_14;
  reg                 io_A_Valid_0_delay_5_13;
  reg                 io_A_Valid_0_delay_6_12;
  reg                 io_A_Valid_0_delay_7_11;
  reg                 io_A_Valid_0_delay_8_10;
  reg                 io_A_Valid_0_delay_9_9;
  reg                 io_A_Valid_0_delay_10_8;
  reg                 io_A_Valid_0_delay_11_7;
  reg                 io_A_Valid_0_delay_12_6;
  reg                 io_A_Valid_0_delay_13_5;
  reg                 io_A_Valid_0_delay_14_4;
  reg                 io_A_Valid_0_delay_15_3;
  reg                 io_A_Valid_0_delay_16_2;
  reg                 io_A_Valid_0_delay_17_1;
  reg                 io_A_Valid_0_delay_18;
  reg                 io_A_Valid_0_delay_1_18;
  reg                 io_A_Valid_0_delay_2_17;
  reg                 io_A_Valid_0_delay_3_16;
  reg                 io_A_Valid_0_delay_4_15;
  reg                 io_A_Valid_0_delay_5_14;
  reg                 io_A_Valid_0_delay_6_13;
  reg                 io_A_Valid_0_delay_7_12;
  reg                 io_A_Valid_0_delay_8_11;
  reg                 io_A_Valid_0_delay_9_10;
  reg                 io_A_Valid_0_delay_10_9;
  reg                 io_A_Valid_0_delay_11_8;
  reg                 io_A_Valid_0_delay_12_7;
  reg                 io_A_Valid_0_delay_13_6;
  reg                 io_A_Valid_0_delay_14_5;
  reg                 io_A_Valid_0_delay_15_4;
  reg                 io_A_Valid_0_delay_16_3;
  reg                 io_A_Valid_0_delay_17_2;
  reg                 io_A_Valid_0_delay_18_1;
  reg                 io_A_Valid_0_delay_19;
  reg                 io_A_Valid_0_delay_1_19;
  reg                 io_A_Valid_0_delay_2_18;
  reg                 io_A_Valid_0_delay_3_17;
  reg                 io_A_Valid_0_delay_4_16;
  reg                 io_A_Valid_0_delay_5_15;
  reg                 io_A_Valid_0_delay_6_14;
  reg                 io_A_Valid_0_delay_7_13;
  reg                 io_A_Valid_0_delay_8_12;
  reg                 io_A_Valid_0_delay_9_11;
  reg                 io_A_Valid_0_delay_10_10;
  reg                 io_A_Valid_0_delay_11_9;
  reg                 io_A_Valid_0_delay_12_8;
  reg                 io_A_Valid_0_delay_13_7;
  reg                 io_A_Valid_0_delay_14_6;
  reg                 io_A_Valid_0_delay_15_5;
  reg                 io_A_Valid_0_delay_16_4;
  reg                 io_A_Valid_0_delay_17_3;
  reg                 io_A_Valid_0_delay_18_2;
  reg                 io_A_Valid_0_delay_19_1;
  reg                 io_A_Valid_0_delay_20;
  reg                 io_A_Valid_0_delay_1_20;
  reg                 io_A_Valid_0_delay_2_19;
  reg                 io_A_Valid_0_delay_3_18;
  reg                 io_A_Valid_0_delay_4_17;
  reg                 io_A_Valid_0_delay_5_16;
  reg                 io_A_Valid_0_delay_6_15;
  reg                 io_A_Valid_0_delay_7_14;
  reg                 io_A_Valid_0_delay_8_13;
  reg                 io_A_Valid_0_delay_9_12;
  reg                 io_A_Valid_0_delay_10_11;
  reg                 io_A_Valid_0_delay_11_10;
  reg                 io_A_Valid_0_delay_12_9;
  reg                 io_A_Valid_0_delay_13_8;
  reg                 io_A_Valid_0_delay_14_7;
  reg                 io_A_Valid_0_delay_15_6;
  reg                 io_A_Valid_0_delay_16_5;
  reg                 io_A_Valid_0_delay_17_4;
  reg                 io_A_Valid_0_delay_18_3;
  reg                 io_A_Valid_0_delay_19_2;
  reg                 io_A_Valid_0_delay_20_1;
  reg                 io_A_Valid_0_delay_21;
  reg                 io_A_Valid_0_delay_1_21;
  reg                 io_A_Valid_0_delay_2_20;
  reg                 io_A_Valid_0_delay_3_19;
  reg                 io_A_Valid_0_delay_4_18;
  reg                 io_A_Valid_0_delay_5_17;
  reg                 io_A_Valid_0_delay_6_16;
  reg                 io_A_Valid_0_delay_7_15;
  reg                 io_A_Valid_0_delay_8_14;
  reg                 io_A_Valid_0_delay_9_13;
  reg                 io_A_Valid_0_delay_10_12;
  reg                 io_A_Valid_0_delay_11_11;
  reg                 io_A_Valid_0_delay_12_10;
  reg                 io_A_Valid_0_delay_13_9;
  reg                 io_A_Valid_0_delay_14_8;
  reg                 io_A_Valid_0_delay_15_7;
  reg                 io_A_Valid_0_delay_16_6;
  reg                 io_A_Valid_0_delay_17_5;
  reg                 io_A_Valid_0_delay_18_4;
  reg                 io_A_Valid_0_delay_19_3;
  reg                 io_A_Valid_0_delay_20_2;
  reg                 io_A_Valid_0_delay_21_1;
  reg                 io_A_Valid_0_delay_22;
  reg                 io_A_Valid_0_delay_1_22;
  reg                 io_A_Valid_0_delay_2_21;
  reg                 io_A_Valid_0_delay_3_20;
  reg                 io_A_Valid_0_delay_4_19;
  reg                 io_A_Valid_0_delay_5_18;
  reg                 io_A_Valid_0_delay_6_17;
  reg                 io_A_Valid_0_delay_7_16;
  reg                 io_A_Valid_0_delay_8_15;
  reg                 io_A_Valid_0_delay_9_14;
  reg                 io_A_Valid_0_delay_10_13;
  reg                 io_A_Valid_0_delay_11_12;
  reg                 io_A_Valid_0_delay_12_11;
  reg                 io_A_Valid_0_delay_13_10;
  reg                 io_A_Valid_0_delay_14_9;
  reg                 io_A_Valid_0_delay_15_8;
  reg                 io_A_Valid_0_delay_16_7;
  reg                 io_A_Valid_0_delay_17_6;
  reg                 io_A_Valid_0_delay_18_5;
  reg                 io_A_Valid_0_delay_19_4;
  reg                 io_A_Valid_0_delay_20_3;
  reg                 io_A_Valid_0_delay_21_2;
  reg                 io_A_Valid_0_delay_22_1;
  reg                 io_A_Valid_0_delay_23;
  reg                 io_A_Valid_0_delay_1_23;
  reg                 io_A_Valid_0_delay_2_22;
  reg                 io_A_Valid_0_delay_3_21;
  reg                 io_A_Valid_0_delay_4_20;
  reg                 io_A_Valid_0_delay_5_19;
  reg                 io_A_Valid_0_delay_6_18;
  reg                 io_A_Valid_0_delay_7_17;
  reg                 io_A_Valid_0_delay_8_16;
  reg                 io_A_Valid_0_delay_9_15;
  reg                 io_A_Valid_0_delay_10_14;
  reg                 io_A_Valid_0_delay_11_13;
  reg                 io_A_Valid_0_delay_12_12;
  reg                 io_A_Valid_0_delay_13_11;
  reg                 io_A_Valid_0_delay_14_10;
  reg                 io_A_Valid_0_delay_15_9;
  reg                 io_A_Valid_0_delay_16_8;
  reg                 io_A_Valid_0_delay_17_7;
  reg                 io_A_Valid_0_delay_18_6;
  reg                 io_A_Valid_0_delay_19_5;
  reg                 io_A_Valid_0_delay_20_4;
  reg                 io_A_Valid_0_delay_21_3;
  reg                 io_A_Valid_0_delay_22_2;
  reg                 io_A_Valid_0_delay_23_1;
  reg                 io_A_Valid_0_delay_24;
  reg                 io_A_Valid_0_delay_1_24;
  reg                 io_A_Valid_0_delay_2_23;
  reg                 io_A_Valid_0_delay_3_22;
  reg                 io_A_Valid_0_delay_4_21;
  reg                 io_A_Valid_0_delay_5_20;
  reg                 io_A_Valid_0_delay_6_19;
  reg                 io_A_Valid_0_delay_7_18;
  reg                 io_A_Valid_0_delay_8_17;
  reg                 io_A_Valid_0_delay_9_16;
  reg                 io_A_Valid_0_delay_10_15;
  reg                 io_A_Valid_0_delay_11_14;
  reg                 io_A_Valid_0_delay_12_13;
  reg                 io_A_Valid_0_delay_13_12;
  reg                 io_A_Valid_0_delay_14_11;
  reg                 io_A_Valid_0_delay_15_10;
  reg                 io_A_Valid_0_delay_16_9;
  reg                 io_A_Valid_0_delay_17_8;
  reg                 io_A_Valid_0_delay_18_7;
  reg                 io_A_Valid_0_delay_19_6;
  reg                 io_A_Valid_0_delay_20_5;
  reg                 io_A_Valid_0_delay_21_4;
  reg                 io_A_Valid_0_delay_22_3;
  reg                 io_A_Valid_0_delay_23_2;
  reg                 io_A_Valid_0_delay_24_1;
  reg                 io_A_Valid_0_delay_25;
  reg                 io_A_Valid_0_delay_1_25;
  reg                 io_A_Valid_0_delay_2_24;
  reg                 io_A_Valid_0_delay_3_23;
  reg                 io_A_Valid_0_delay_4_22;
  reg                 io_A_Valid_0_delay_5_21;
  reg                 io_A_Valid_0_delay_6_20;
  reg                 io_A_Valid_0_delay_7_19;
  reg                 io_A_Valid_0_delay_8_18;
  reg                 io_A_Valid_0_delay_9_17;
  reg                 io_A_Valid_0_delay_10_16;
  reg                 io_A_Valid_0_delay_11_15;
  reg                 io_A_Valid_0_delay_12_14;
  reg                 io_A_Valid_0_delay_13_13;
  reg                 io_A_Valid_0_delay_14_12;
  reg                 io_A_Valid_0_delay_15_11;
  reg                 io_A_Valid_0_delay_16_10;
  reg                 io_A_Valid_0_delay_17_9;
  reg                 io_A_Valid_0_delay_18_8;
  reg                 io_A_Valid_0_delay_19_7;
  reg                 io_A_Valid_0_delay_20_6;
  reg                 io_A_Valid_0_delay_21_5;
  reg                 io_A_Valid_0_delay_22_4;
  reg                 io_A_Valid_0_delay_23_3;
  reg                 io_A_Valid_0_delay_24_2;
  reg                 io_A_Valid_0_delay_25_1;
  reg                 io_A_Valid_0_delay_26;
  reg                 io_A_Valid_0_delay_1_26;
  reg                 io_A_Valid_0_delay_2_25;
  reg                 io_A_Valid_0_delay_3_24;
  reg                 io_A_Valid_0_delay_4_23;
  reg                 io_A_Valid_0_delay_5_22;
  reg                 io_A_Valid_0_delay_6_21;
  reg                 io_A_Valid_0_delay_7_20;
  reg                 io_A_Valid_0_delay_8_19;
  reg                 io_A_Valid_0_delay_9_18;
  reg                 io_A_Valid_0_delay_10_17;
  reg                 io_A_Valid_0_delay_11_16;
  reg                 io_A_Valid_0_delay_12_15;
  reg                 io_A_Valid_0_delay_13_14;
  reg                 io_A_Valid_0_delay_14_13;
  reg                 io_A_Valid_0_delay_15_12;
  reg                 io_A_Valid_0_delay_16_11;
  reg                 io_A_Valid_0_delay_17_10;
  reg                 io_A_Valid_0_delay_18_9;
  reg                 io_A_Valid_0_delay_19_8;
  reg                 io_A_Valid_0_delay_20_7;
  reg                 io_A_Valid_0_delay_21_6;
  reg                 io_A_Valid_0_delay_22_5;
  reg                 io_A_Valid_0_delay_23_4;
  reg                 io_A_Valid_0_delay_24_3;
  reg                 io_A_Valid_0_delay_25_2;
  reg                 io_A_Valid_0_delay_26_1;
  reg                 io_A_Valid_0_delay_27;
  reg                 io_A_Valid_0_delay_1_27;
  reg                 io_A_Valid_0_delay_2_26;
  reg                 io_A_Valid_0_delay_3_25;
  reg                 io_A_Valid_0_delay_4_24;
  reg                 io_A_Valid_0_delay_5_23;
  reg                 io_A_Valid_0_delay_6_22;
  reg                 io_A_Valid_0_delay_7_21;
  reg                 io_A_Valid_0_delay_8_20;
  reg                 io_A_Valid_0_delay_9_19;
  reg                 io_A_Valid_0_delay_10_18;
  reg                 io_A_Valid_0_delay_11_17;
  reg                 io_A_Valid_0_delay_12_16;
  reg                 io_A_Valid_0_delay_13_15;
  reg                 io_A_Valid_0_delay_14_14;
  reg                 io_A_Valid_0_delay_15_13;
  reg                 io_A_Valid_0_delay_16_12;
  reg                 io_A_Valid_0_delay_17_11;
  reg                 io_A_Valid_0_delay_18_10;
  reg                 io_A_Valid_0_delay_19_9;
  reg                 io_A_Valid_0_delay_20_8;
  reg                 io_A_Valid_0_delay_21_7;
  reg                 io_A_Valid_0_delay_22_6;
  reg                 io_A_Valid_0_delay_23_5;
  reg                 io_A_Valid_0_delay_24_4;
  reg                 io_A_Valid_0_delay_25_3;
  reg                 io_A_Valid_0_delay_26_2;
  reg                 io_A_Valid_0_delay_27_1;
  reg                 io_A_Valid_0_delay_28;
  reg                 io_A_Valid_0_delay_1_28;
  reg                 io_A_Valid_0_delay_2_27;
  reg                 io_A_Valid_0_delay_3_26;
  reg                 io_A_Valid_0_delay_4_25;
  reg                 io_A_Valid_0_delay_5_24;
  reg                 io_A_Valid_0_delay_6_23;
  reg                 io_A_Valid_0_delay_7_22;
  reg                 io_A_Valid_0_delay_8_21;
  reg                 io_A_Valid_0_delay_9_20;
  reg                 io_A_Valid_0_delay_10_19;
  reg                 io_A_Valid_0_delay_11_18;
  reg                 io_A_Valid_0_delay_12_17;
  reg                 io_A_Valid_0_delay_13_16;
  reg                 io_A_Valid_0_delay_14_15;
  reg                 io_A_Valid_0_delay_15_14;
  reg                 io_A_Valid_0_delay_16_13;
  reg                 io_A_Valid_0_delay_17_12;
  reg                 io_A_Valid_0_delay_18_11;
  reg                 io_A_Valid_0_delay_19_10;
  reg                 io_A_Valid_0_delay_20_9;
  reg                 io_A_Valid_0_delay_21_8;
  reg                 io_A_Valid_0_delay_22_7;
  reg                 io_A_Valid_0_delay_23_6;
  reg                 io_A_Valid_0_delay_24_5;
  reg                 io_A_Valid_0_delay_25_4;
  reg                 io_A_Valid_0_delay_26_3;
  reg                 io_A_Valid_0_delay_27_2;
  reg                 io_A_Valid_0_delay_28_1;
  reg                 io_A_Valid_0_delay_29;
  reg                 io_A_Valid_0_delay_1_29;
  reg                 io_A_Valid_0_delay_2_28;
  reg                 io_A_Valid_0_delay_3_27;
  reg                 io_A_Valid_0_delay_4_26;
  reg                 io_A_Valid_0_delay_5_25;
  reg                 io_A_Valid_0_delay_6_24;
  reg                 io_A_Valid_0_delay_7_23;
  reg                 io_A_Valid_0_delay_8_22;
  reg                 io_A_Valid_0_delay_9_21;
  reg                 io_A_Valid_0_delay_10_20;
  reg                 io_A_Valid_0_delay_11_19;
  reg                 io_A_Valid_0_delay_12_18;
  reg                 io_A_Valid_0_delay_13_17;
  reg                 io_A_Valid_0_delay_14_16;
  reg                 io_A_Valid_0_delay_15_15;
  reg                 io_A_Valid_0_delay_16_14;
  reg                 io_A_Valid_0_delay_17_13;
  reg                 io_A_Valid_0_delay_18_12;
  reg                 io_A_Valid_0_delay_19_11;
  reg                 io_A_Valid_0_delay_20_10;
  reg                 io_A_Valid_0_delay_21_9;
  reg                 io_A_Valid_0_delay_22_8;
  reg                 io_A_Valid_0_delay_23_7;
  reg                 io_A_Valid_0_delay_24_6;
  reg                 io_A_Valid_0_delay_25_5;
  reg                 io_A_Valid_0_delay_26_4;
  reg                 io_A_Valid_0_delay_27_3;
  reg                 io_A_Valid_0_delay_28_2;
  reg                 io_A_Valid_0_delay_29_1;
  reg                 io_A_Valid_0_delay_30;
  reg                 io_A_Valid_0_delay_1_30;
  reg                 io_A_Valid_0_delay_2_29;
  reg                 io_A_Valid_0_delay_3_28;
  reg                 io_A_Valid_0_delay_4_27;
  reg                 io_A_Valid_0_delay_5_26;
  reg                 io_A_Valid_0_delay_6_25;
  reg                 io_A_Valid_0_delay_7_24;
  reg                 io_A_Valid_0_delay_8_23;
  reg                 io_A_Valid_0_delay_9_22;
  reg                 io_A_Valid_0_delay_10_21;
  reg                 io_A_Valid_0_delay_11_20;
  reg                 io_A_Valid_0_delay_12_19;
  reg                 io_A_Valid_0_delay_13_18;
  reg                 io_A_Valid_0_delay_14_17;
  reg                 io_A_Valid_0_delay_15_16;
  reg                 io_A_Valid_0_delay_16_15;
  reg                 io_A_Valid_0_delay_17_14;
  reg                 io_A_Valid_0_delay_18_13;
  reg                 io_A_Valid_0_delay_19_12;
  reg                 io_A_Valid_0_delay_20_11;
  reg                 io_A_Valid_0_delay_21_10;
  reg                 io_A_Valid_0_delay_22_9;
  reg                 io_A_Valid_0_delay_23_8;
  reg                 io_A_Valid_0_delay_24_7;
  reg                 io_A_Valid_0_delay_25_6;
  reg                 io_A_Valid_0_delay_26_5;
  reg                 io_A_Valid_0_delay_27_4;
  reg                 io_A_Valid_0_delay_28_3;
  reg                 io_A_Valid_0_delay_29_2;
  reg                 io_A_Valid_0_delay_30_1;
  reg                 io_A_Valid_0_delay_31;
  reg                 io_A_Valid_0_delay_1_31;
  reg                 io_A_Valid_0_delay_2_30;
  reg                 io_A_Valid_0_delay_3_29;
  reg                 io_A_Valid_0_delay_4_28;
  reg                 io_A_Valid_0_delay_5_27;
  reg                 io_A_Valid_0_delay_6_26;
  reg                 io_A_Valid_0_delay_7_25;
  reg                 io_A_Valid_0_delay_8_24;
  reg                 io_A_Valid_0_delay_9_23;
  reg                 io_A_Valid_0_delay_10_22;
  reg                 io_A_Valid_0_delay_11_21;
  reg                 io_A_Valid_0_delay_12_20;
  reg                 io_A_Valid_0_delay_13_19;
  reg                 io_A_Valid_0_delay_14_18;
  reg                 io_A_Valid_0_delay_15_17;
  reg                 io_A_Valid_0_delay_16_16;
  reg                 io_A_Valid_0_delay_17_15;
  reg                 io_A_Valid_0_delay_18_14;
  reg                 io_A_Valid_0_delay_19_13;
  reg                 io_A_Valid_0_delay_20_12;
  reg                 io_A_Valid_0_delay_21_11;
  reg                 io_A_Valid_0_delay_22_10;
  reg                 io_A_Valid_0_delay_23_9;
  reg                 io_A_Valid_0_delay_24_8;
  reg                 io_A_Valid_0_delay_25_7;
  reg                 io_A_Valid_0_delay_26_6;
  reg                 io_A_Valid_0_delay_27_5;
  reg                 io_A_Valid_0_delay_28_4;
  reg                 io_A_Valid_0_delay_29_3;
  reg                 io_A_Valid_0_delay_30_2;
  reg                 io_A_Valid_0_delay_31_1;
  reg                 io_A_Valid_0_delay_32;
  reg                 io_A_Valid_0_delay_1_32;
  reg                 io_A_Valid_0_delay_2_31;
  reg                 io_A_Valid_0_delay_3_30;
  reg                 io_A_Valid_0_delay_4_29;
  reg                 io_A_Valid_0_delay_5_28;
  reg                 io_A_Valid_0_delay_6_27;
  reg                 io_A_Valid_0_delay_7_26;
  reg                 io_A_Valid_0_delay_8_25;
  reg                 io_A_Valid_0_delay_9_24;
  reg                 io_A_Valid_0_delay_10_23;
  reg                 io_A_Valid_0_delay_11_22;
  reg                 io_A_Valid_0_delay_12_21;
  reg                 io_A_Valid_0_delay_13_20;
  reg                 io_A_Valid_0_delay_14_19;
  reg                 io_A_Valid_0_delay_15_18;
  reg                 io_A_Valid_0_delay_16_17;
  reg                 io_A_Valid_0_delay_17_16;
  reg                 io_A_Valid_0_delay_18_15;
  reg                 io_A_Valid_0_delay_19_14;
  reg                 io_A_Valid_0_delay_20_13;
  reg                 io_A_Valid_0_delay_21_12;
  reg                 io_A_Valid_0_delay_22_11;
  reg                 io_A_Valid_0_delay_23_10;
  reg                 io_A_Valid_0_delay_24_9;
  reg                 io_A_Valid_0_delay_25_8;
  reg                 io_A_Valid_0_delay_26_7;
  reg                 io_A_Valid_0_delay_27_6;
  reg                 io_A_Valid_0_delay_28_5;
  reg                 io_A_Valid_0_delay_29_4;
  reg                 io_A_Valid_0_delay_30_3;
  reg                 io_A_Valid_0_delay_31_2;
  reg                 io_A_Valid_0_delay_32_1;
  reg                 io_A_Valid_0_delay_33;
  reg                 io_A_Valid_0_delay_1_33;
  reg                 io_A_Valid_0_delay_2_32;
  reg                 io_A_Valid_0_delay_3_31;
  reg                 io_A_Valid_0_delay_4_30;
  reg                 io_A_Valid_0_delay_5_29;
  reg                 io_A_Valid_0_delay_6_28;
  reg                 io_A_Valid_0_delay_7_27;
  reg                 io_A_Valid_0_delay_8_26;
  reg                 io_A_Valid_0_delay_9_25;
  reg                 io_A_Valid_0_delay_10_24;
  reg                 io_A_Valid_0_delay_11_23;
  reg                 io_A_Valid_0_delay_12_22;
  reg                 io_A_Valid_0_delay_13_21;
  reg                 io_A_Valid_0_delay_14_20;
  reg                 io_A_Valid_0_delay_15_19;
  reg                 io_A_Valid_0_delay_16_18;
  reg                 io_A_Valid_0_delay_17_17;
  reg                 io_A_Valid_0_delay_18_16;
  reg                 io_A_Valid_0_delay_19_15;
  reg                 io_A_Valid_0_delay_20_14;
  reg                 io_A_Valid_0_delay_21_13;
  reg                 io_A_Valid_0_delay_22_12;
  reg                 io_A_Valid_0_delay_23_11;
  reg                 io_A_Valid_0_delay_24_10;
  reg                 io_A_Valid_0_delay_25_9;
  reg                 io_A_Valid_0_delay_26_8;
  reg                 io_A_Valid_0_delay_27_7;
  reg                 io_A_Valid_0_delay_28_6;
  reg                 io_A_Valid_0_delay_29_5;
  reg                 io_A_Valid_0_delay_30_4;
  reg                 io_A_Valid_0_delay_31_3;
  reg                 io_A_Valid_0_delay_32_2;
  reg                 io_A_Valid_0_delay_33_1;
  reg                 io_A_Valid_0_delay_34;
  reg                 io_A_Valid_0_delay_1_34;
  reg                 io_A_Valid_0_delay_2_33;
  reg                 io_A_Valid_0_delay_3_32;
  reg                 io_A_Valid_0_delay_4_31;
  reg                 io_A_Valid_0_delay_5_30;
  reg                 io_A_Valid_0_delay_6_29;
  reg                 io_A_Valid_0_delay_7_28;
  reg                 io_A_Valid_0_delay_8_27;
  reg                 io_A_Valid_0_delay_9_26;
  reg                 io_A_Valid_0_delay_10_25;
  reg                 io_A_Valid_0_delay_11_24;
  reg                 io_A_Valid_0_delay_12_23;
  reg                 io_A_Valid_0_delay_13_22;
  reg                 io_A_Valid_0_delay_14_21;
  reg                 io_A_Valid_0_delay_15_20;
  reg                 io_A_Valid_0_delay_16_19;
  reg                 io_A_Valid_0_delay_17_18;
  reg                 io_A_Valid_0_delay_18_17;
  reg                 io_A_Valid_0_delay_19_16;
  reg                 io_A_Valid_0_delay_20_15;
  reg                 io_A_Valid_0_delay_21_14;
  reg                 io_A_Valid_0_delay_22_13;
  reg                 io_A_Valid_0_delay_23_12;
  reg                 io_A_Valid_0_delay_24_11;
  reg                 io_A_Valid_0_delay_25_10;
  reg                 io_A_Valid_0_delay_26_9;
  reg                 io_A_Valid_0_delay_27_8;
  reg                 io_A_Valid_0_delay_28_7;
  reg                 io_A_Valid_0_delay_29_6;
  reg                 io_A_Valid_0_delay_30_5;
  reg                 io_A_Valid_0_delay_31_4;
  reg                 io_A_Valid_0_delay_32_3;
  reg                 io_A_Valid_0_delay_33_2;
  reg                 io_A_Valid_0_delay_34_1;
  reg                 io_A_Valid_0_delay_35;
  reg                 io_A_Valid_0_delay_1_35;
  reg                 io_A_Valid_0_delay_2_34;
  reg                 io_A_Valid_0_delay_3_33;
  reg                 io_A_Valid_0_delay_4_32;
  reg                 io_A_Valid_0_delay_5_31;
  reg                 io_A_Valid_0_delay_6_30;
  reg                 io_A_Valid_0_delay_7_29;
  reg                 io_A_Valid_0_delay_8_28;
  reg                 io_A_Valid_0_delay_9_27;
  reg                 io_A_Valid_0_delay_10_26;
  reg                 io_A_Valid_0_delay_11_25;
  reg                 io_A_Valid_0_delay_12_24;
  reg                 io_A_Valid_0_delay_13_23;
  reg                 io_A_Valid_0_delay_14_22;
  reg                 io_A_Valid_0_delay_15_21;
  reg                 io_A_Valid_0_delay_16_20;
  reg                 io_A_Valid_0_delay_17_19;
  reg                 io_A_Valid_0_delay_18_18;
  reg                 io_A_Valid_0_delay_19_17;
  reg                 io_A_Valid_0_delay_20_16;
  reg                 io_A_Valid_0_delay_21_15;
  reg                 io_A_Valid_0_delay_22_14;
  reg                 io_A_Valid_0_delay_23_13;
  reg                 io_A_Valid_0_delay_24_12;
  reg                 io_A_Valid_0_delay_25_11;
  reg                 io_A_Valid_0_delay_26_10;
  reg                 io_A_Valid_0_delay_27_9;
  reg                 io_A_Valid_0_delay_28_8;
  reg                 io_A_Valid_0_delay_29_7;
  reg                 io_A_Valid_0_delay_30_6;
  reg                 io_A_Valid_0_delay_31_5;
  reg                 io_A_Valid_0_delay_32_4;
  reg                 io_A_Valid_0_delay_33_3;
  reg                 io_A_Valid_0_delay_34_2;
  reg                 io_A_Valid_0_delay_35_1;
  reg                 io_A_Valid_0_delay_36;
  reg                 io_A_Valid_0_delay_1_36;
  reg                 io_A_Valid_0_delay_2_35;
  reg                 io_A_Valid_0_delay_3_34;
  reg                 io_A_Valid_0_delay_4_33;
  reg                 io_A_Valid_0_delay_5_32;
  reg                 io_A_Valid_0_delay_6_31;
  reg                 io_A_Valid_0_delay_7_30;
  reg                 io_A_Valid_0_delay_8_29;
  reg                 io_A_Valid_0_delay_9_28;
  reg                 io_A_Valid_0_delay_10_27;
  reg                 io_A_Valid_0_delay_11_26;
  reg                 io_A_Valid_0_delay_12_25;
  reg                 io_A_Valid_0_delay_13_24;
  reg                 io_A_Valid_0_delay_14_23;
  reg                 io_A_Valid_0_delay_15_22;
  reg                 io_A_Valid_0_delay_16_21;
  reg                 io_A_Valid_0_delay_17_20;
  reg                 io_A_Valid_0_delay_18_19;
  reg                 io_A_Valid_0_delay_19_18;
  reg                 io_A_Valid_0_delay_20_17;
  reg                 io_A_Valid_0_delay_21_16;
  reg                 io_A_Valid_0_delay_22_15;
  reg                 io_A_Valid_0_delay_23_14;
  reg                 io_A_Valid_0_delay_24_13;
  reg                 io_A_Valid_0_delay_25_12;
  reg                 io_A_Valid_0_delay_26_11;
  reg                 io_A_Valid_0_delay_27_10;
  reg                 io_A_Valid_0_delay_28_9;
  reg                 io_A_Valid_0_delay_29_8;
  reg                 io_A_Valid_0_delay_30_7;
  reg                 io_A_Valid_0_delay_31_6;
  reg                 io_A_Valid_0_delay_32_5;
  reg                 io_A_Valid_0_delay_33_4;
  reg                 io_A_Valid_0_delay_34_3;
  reg                 io_A_Valid_0_delay_35_2;
  reg                 io_A_Valid_0_delay_36_1;
  reg                 io_A_Valid_0_delay_37;
  reg                 io_A_Valid_0_delay_1_37;
  reg                 io_A_Valid_0_delay_2_36;
  reg                 io_A_Valid_0_delay_3_35;
  reg                 io_A_Valid_0_delay_4_34;
  reg                 io_A_Valid_0_delay_5_33;
  reg                 io_A_Valid_0_delay_6_32;
  reg                 io_A_Valid_0_delay_7_31;
  reg                 io_A_Valid_0_delay_8_30;
  reg                 io_A_Valid_0_delay_9_29;
  reg                 io_A_Valid_0_delay_10_28;
  reg                 io_A_Valid_0_delay_11_27;
  reg                 io_A_Valid_0_delay_12_26;
  reg                 io_A_Valid_0_delay_13_25;
  reg                 io_A_Valid_0_delay_14_24;
  reg                 io_A_Valid_0_delay_15_23;
  reg                 io_A_Valid_0_delay_16_22;
  reg                 io_A_Valid_0_delay_17_21;
  reg                 io_A_Valid_0_delay_18_20;
  reg                 io_A_Valid_0_delay_19_19;
  reg                 io_A_Valid_0_delay_20_18;
  reg                 io_A_Valid_0_delay_21_17;
  reg                 io_A_Valid_0_delay_22_16;
  reg                 io_A_Valid_0_delay_23_15;
  reg                 io_A_Valid_0_delay_24_14;
  reg                 io_A_Valid_0_delay_25_13;
  reg                 io_A_Valid_0_delay_26_12;
  reg                 io_A_Valid_0_delay_27_11;
  reg                 io_A_Valid_0_delay_28_10;
  reg                 io_A_Valid_0_delay_29_9;
  reg                 io_A_Valid_0_delay_30_8;
  reg                 io_A_Valid_0_delay_31_7;
  reg                 io_A_Valid_0_delay_32_6;
  reg                 io_A_Valid_0_delay_33_5;
  reg                 io_A_Valid_0_delay_34_4;
  reg                 io_A_Valid_0_delay_35_3;
  reg                 io_A_Valid_0_delay_36_2;
  reg                 io_A_Valid_0_delay_37_1;
  reg                 io_A_Valid_0_delay_38;
  reg                 io_A_Valid_0_delay_1_38;
  reg                 io_A_Valid_0_delay_2_37;
  reg                 io_A_Valid_0_delay_3_36;
  reg                 io_A_Valid_0_delay_4_35;
  reg                 io_A_Valid_0_delay_5_34;
  reg                 io_A_Valid_0_delay_6_33;
  reg                 io_A_Valid_0_delay_7_32;
  reg                 io_A_Valid_0_delay_8_31;
  reg                 io_A_Valid_0_delay_9_30;
  reg                 io_A_Valid_0_delay_10_29;
  reg                 io_A_Valid_0_delay_11_28;
  reg                 io_A_Valid_0_delay_12_27;
  reg                 io_A_Valid_0_delay_13_26;
  reg                 io_A_Valid_0_delay_14_25;
  reg                 io_A_Valid_0_delay_15_24;
  reg                 io_A_Valid_0_delay_16_23;
  reg                 io_A_Valid_0_delay_17_22;
  reg                 io_A_Valid_0_delay_18_21;
  reg                 io_A_Valid_0_delay_19_20;
  reg                 io_A_Valid_0_delay_20_19;
  reg                 io_A_Valid_0_delay_21_18;
  reg                 io_A_Valid_0_delay_22_17;
  reg                 io_A_Valid_0_delay_23_16;
  reg                 io_A_Valid_0_delay_24_15;
  reg                 io_A_Valid_0_delay_25_14;
  reg                 io_A_Valid_0_delay_26_13;
  reg                 io_A_Valid_0_delay_27_12;
  reg                 io_A_Valid_0_delay_28_11;
  reg                 io_A_Valid_0_delay_29_10;
  reg                 io_A_Valid_0_delay_30_9;
  reg                 io_A_Valid_0_delay_31_8;
  reg                 io_A_Valid_0_delay_32_7;
  reg                 io_A_Valid_0_delay_33_6;
  reg                 io_A_Valid_0_delay_34_5;
  reg                 io_A_Valid_0_delay_35_4;
  reg                 io_A_Valid_0_delay_36_3;
  reg                 io_A_Valid_0_delay_37_2;
  reg                 io_A_Valid_0_delay_38_1;
  reg                 io_A_Valid_0_delay_39;
  reg                 io_A_Valid_0_delay_1_39;
  reg                 io_A_Valid_0_delay_2_38;
  reg                 io_A_Valid_0_delay_3_37;
  reg                 io_A_Valid_0_delay_4_36;
  reg                 io_A_Valid_0_delay_5_35;
  reg                 io_A_Valid_0_delay_6_34;
  reg                 io_A_Valid_0_delay_7_33;
  reg                 io_A_Valid_0_delay_8_32;
  reg                 io_A_Valid_0_delay_9_31;
  reg                 io_A_Valid_0_delay_10_30;
  reg                 io_A_Valid_0_delay_11_29;
  reg                 io_A_Valid_0_delay_12_28;
  reg                 io_A_Valid_0_delay_13_27;
  reg                 io_A_Valid_0_delay_14_26;
  reg                 io_A_Valid_0_delay_15_25;
  reg                 io_A_Valid_0_delay_16_24;
  reg                 io_A_Valid_0_delay_17_23;
  reg                 io_A_Valid_0_delay_18_22;
  reg                 io_A_Valid_0_delay_19_21;
  reg                 io_A_Valid_0_delay_20_20;
  reg                 io_A_Valid_0_delay_21_19;
  reg                 io_A_Valid_0_delay_22_18;
  reg                 io_A_Valid_0_delay_23_17;
  reg                 io_A_Valid_0_delay_24_16;
  reg                 io_A_Valid_0_delay_25_15;
  reg                 io_A_Valid_0_delay_26_14;
  reg                 io_A_Valid_0_delay_27_13;
  reg                 io_A_Valid_0_delay_28_12;
  reg                 io_A_Valid_0_delay_29_11;
  reg                 io_A_Valid_0_delay_30_10;
  reg                 io_A_Valid_0_delay_31_9;
  reg                 io_A_Valid_0_delay_32_8;
  reg                 io_A_Valid_0_delay_33_7;
  reg                 io_A_Valid_0_delay_34_6;
  reg                 io_A_Valid_0_delay_35_5;
  reg                 io_A_Valid_0_delay_36_4;
  reg                 io_A_Valid_0_delay_37_3;
  reg                 io_A_Valid_0_delay_38_2;
  reg                 io_A_Valid_0_delay_39_1;
  reg                 io_A_Valid_0_delay_40;
  reg                 io_A_Valid_0_delay_1_40;
  reg                 io_A_Valid_0_delay_2_39;
  reg                 io_A_Valid_0_delay_3_38;
  reg                 io_A_Valid_0_delay_4_37;
  reg                 io_A_Valid_0_delay_5_36;
  reg                 io_A_Valid_0_delay_6_35;
  reg                 io_A_Valid_0_delay_7_34;
  reg                 io_A_Valid_0_delay_8_33;
  reg                 io_A_Valid_0_delay_9_32;
  reg                 io_A_Valid_0_delay_10_31;
  reg                 io_A_Valid_0_delay_11_30;
  reg                 io_A_Valid_0_delay_12_29;
  reg                 io_A_Valid_0_delay_13_28;
  reg                 io_A_Valid_0_delay_14_27;
  reg                 io_A_Valid_0_delay_15_26;
  reg                 io_A_Valid_0_delay_16_25;
  reg                 io_A_Valid_0_delay_17_24;
  reg                 io_A_Valid_0_delay_18_23;
  reg                 io_A_Valid_0_delay_19_22;
  reg                 io_A_Valid_0_delay_20_21;
  reg                 io_A_Valid_0_delay_21_20;
  reg                 io_A_Valid_0_delay_22_19;
  reg                 io_A_Valid_0_delay_23_18;
  reg                 io_A_Valid_0_delay_24_17;
  reg                 io_A_Valid_0_delay_25_16;
  reg                 io_A_Valid_0_delay_26_15;
  reg                 io_A_Valid_0_delay_27_14;
  reg                 io_A_Valid_0_delay_28_13;
  reg                 io_A_Valid_0_delay_29_12;
  reg                 io_A_Valid_0_delay_30_11;
  reg                 io_A_Valid_0_delay_31_10;
  reg                 io_A_Valid_0_delay_32_9;
  reg                 io_A_Valid_0_delay_33_8;
  reg                 io_A_Valid_0_delay_34_7;
  reg                 io_A_Valid_0_delay_35_6;
  reg                 io_A_Valid_0_delay_36_5;
  reg                 io_A_Valid_0_delay_37_4;
  reg                 io_A_Valid_0_delay_38_3;
  reg                 io_A_Valid_0_delay_39_2;
  reg                 io_A_Valid_0_delay_40_1;
  reg                 io_A_Valid_0_delay_41;
  reg                 io_A_Valid_0_delay_1_41;
  reg                 io_A_Valid_0_delay_2_40;
  reg                 io_A_Valid_0_delay_3_39;
  reg                 io_A_Valid_0_delay_4_38;
  reg                 io_A_Valid_0_delay_5_37;
  reg                 io_A_Valid_0_delay_6_36;
  reg                 io_A_Valid_0_delay_7_35;
  reg                 io_A_Valid_0_delay_8_34;
  reg                 io_A_Valid_0_delay_9_33;
  reg                 io_A_Valid_0_delay_10_32;
  reg                 io_A_Valid_0_delay_11_31;
  reg                 io_A_Valid_0_delay_12_30;
  reg                 io_A_Valid_0_delay_13_29;
  reg                 io_A_Valid_0_delay_14_28;
  reg                 io_A_Valid_0_delay_15_27;
  reg                 io_A_Valid_0_delay_16_26;
  reg                 io_A_Valid_0_delay_17_25;
  reg                 io_A_Valid_0_delay_18_24;
  reg                 io_A_Valid_0_delay_19_23;
  reg                 io_A_Valid_0_delay_20_22;
  reg                 io_A_Valid_0_delay_21_21;
  reg                 io_A_Valid_0_delay_22_20;
  reg                 io_A_Valid_0_delay_23_19;
  reg                 io_A_Valid_0_delay_24_18;
  reg                 io_A_Valid_0_delay_25_17;
  reg                 io_A_Valid_0_delay_26_16;
  reg                 io_A_Valid_0_delay_27_15;
  reg                 io_A_Valid_0_delay_28_14;
  reg                 io_A_Valid_0_delay_29_13;
  reg                 io_A_Valid_0_delay_30_12;
  reg                 io_A_Valid_0_delay_31_11;
  reg                 io_A_Valid_0_delay_32_10;
  reg                 io_A_Valid_0_delay_33_9;
  reg                 io_A_Valid_0_delay_34_8;
  reg                 io_A_Valid_0_delay_35_7;
  reg                 io_A_Valid_0_delay_36_6;
  reg                 io_A_Valid_0_delay_37_5;
  reg                 io_A_Valid_0_delay_38_4;
  reg                 io_A_Valid_0_delay_39_3;
  reg                 io_A_Valid_0_delay_40_2;
  reg                 io_A_Valid_0_delay_41_1;
  reg                 io_A_Valid_0_delay_42;
  reg                 io_A_Valid_0_delay_1_42;
  reg                 io_A_Valid_0_delay_2_41;
  reg                 io_A_Valid_0_delay_3_40;
  reg                 io_A_Valid_0_delay_4_39;
  reg                 io_A_Valid_0_delay_5_38;
  reg                 io_A_Valid_0_delay_6_37;
  reg                 io_A_Valid_0_delay_7_36;
  reg                 io_A_Valid_0_delay_8_35;
  reg                 io_A_Valid_0_delay_9_34;
  reg                 io_A_Valid_0_delay_10_33;
  reg                 io_A_Valid_0_delay_11_32;
  reg                 io_A_Valid_0_delay_12_31;
  reg                 io_A_Valid_0_delay_13_30;
  reg                 io_A_Valid_0_delay_14_29;
  reg                 io_A_Valid_0_delay_15_28;
  reg                 io_A_Valid_0_delay_16_27;
  reg                 io_A_Valid_0_delay_17_26;
  reg                 io_A_Valid_0_delay_18_25;
  reg                 io_A_Valid_0_delay_19_24;
  reg                 io_A_Valid_0_delay_20_23;
  reg                 io_A_Valid_0_delay_21_22;
  reg                 io_A_Valid_0_delay_22_21;
  reg                 io_A_Valid_0_delay_23_20;
  reg                 io_A_Valid_0_delay_24_19;
  reg                 io_A_Valid_0_delay_25_18;
  reg                 io_A_Valid_0_delay_26_17;
  reg                 io_A_Valid_0_delay_27_16;
  reg                 io_A_Valid_0_delay_28_15;
  reg                 io_A_Valid_0_delay_29_14;
  reg                 io_A_Valid_0_delay_30_13;
  reg                 io_A_Valid_0_delay_31_12;
  reg                 io_A_Valid_0_delay_32_11;
  reg                 io_A_Valid_0_delay_33_10;
  reg                 io_A_Valid_0_delay_34_9;
  reg                 io_A_Valid_0_delay_35_8;
  reg                 io_A_Valid_0_delay_36_7;
  reg                 io_A_Valid_0_delay_37_6;
  reg                 io_A_Valid_0_delay_38_5;
  reg                 io_A_Valid_0_delay_39_4;
  reg                 io_A_Valid_0_delay_40_3;
  reg                 io_A_Valid_0_delay_41_2;
  reg                 io_A_Valid_0_delay_42_1;
  reg                 io_A_Valid_0_delay_43;
  reg                 io_A_Valid_0_delay_1_43;
  reg                 io_A_Valid_0_delay_2_42;
  reg                 io_A_Valid_0_delay_3_41;
  reg                 io_A_Valid_0_delay_4_40;
  reg                 io_A_Valid_0_delay_5_39;
  reg                 io_A_Valid_0_delay_6_38;
  reg                 io_A_Valid_0_delay_7_37;
  reg                 io_A_Valid_0_delay_8_36;
  reg                 io_A_Valid_0_delay_9_35;
  reg                 io_A_Valid_0_delay_10_34;
  reg                 io_A_Valid_0_delay_11_33;
  reg                 io_A_Valid_0_delay_12_32;
  reg                 io_A_Valid_0_delay_13_31;
  reg                 io_A_Valid_0_delay_14_30;
  reg                 io_A_Valid_0_delay_15_29;
  reg                 io_A_Valid_0_delay_16_28;
  reg                 io_A_Valid_0_delay_17_27;
  reg                 io_A_Valid_0_delay_18_26;
  reg                 io_A_Valid_0_delay_19_25;
  reg                 io_A_Valid_0_delay_20_24;
  reg                 io_A_Valid_0_delay_21_23;
  reg                 io_A_Valid_0_delay_22_22;
  reg                 io_A_Valid_0_delay_23_21;
  reg                 io_A_Valid_0_delay_24_20;
  reg                 io_A_Valid_0_delay_25_19;
  reg                 io_A_Valid_0_delay_26_18;
  reg                 io_A_Valid_0_delay_27_17;
  reg                 io_A_Valid_0_delay_28_16;
  reg                 io_A_Valid_0_delay_29_15;
  reg                 io_A_Valid_0_delay_30_14;
  reg                 io_A_Valid_0_delay_31_13;
  reg                 io_A_Valid_0_delay_32_12;
  reg                 io_A_Valid_0_delay_33_11;
  reg                 io_A_Valid_0_delay_34_10;
  reg                 io_A_Valid_0_delay_35_9;
  reg                 io_A_Valid_0_delay_36_8;
  reg                 io_A_Valid_0_delay_37_7;
  reg                 io_A_Valid_0_delay_38_6;
  reg                 io_A_Valid_0_delay_39_5;
  reg                 io_A_Valid_0_delay_40_4;
  reg                 io_A_Valid_0_delay_41_3;
  reg                 io_A_Valid_0_delay_42_2;
  reg                 io_A_Valid_0_delay_43_1;
  reg                 io_A_Valid_0_delay_44;
  reg                 io_A_Valid_0_delay_1_44;
  reg                 io_A_Valid_0_delay_2_43;
  reg                 io_A_Valid_0_delay_3_42;
  reg                 io_A_Valid_0_delay_4_41;
  reg                 io_A_Valid_0_delay_5_40;
  reg                 io_A_Valid_0_delay_6_39;
  reg                 io_A_Valid_0_delay_7_38;
  reg                 io_A_Valid_0_delay_8_37;
  reg                 io_A_Valid_0_delay_9_36;
  reg                 io_A_Valid_0_delay_10_35;
  reg                 io_A_Valid_0_delay_11_34;
  reg                 io_A_Valid_0_delay_12_33;
  reg                 io_A_Valid_0_delay_13_32;
  reg                 io_A_Valid_0_delay_14_31;
  reg                 io_A_Valid_0_delay_15_30;
  reg                 io_A_Valid_0_delay_16_29;
  reg                 io_A_Valid_0_delay_17_28;
  reg                 io_A_Valid_0_delay_18_27;
  reg                 io_A_Valid_0_delay_19_26;
  reg                 io_A_Valid_0_delay_20_25;
  reg                 io_A_Valid_0_delay_21_24;
  reg                 io_A_Valid_0_delay_22_23;
  reg                 io_A_Valid_0_delay_23_22;
  reg                 io_A_Valid_0_delay_24_21;
  reg                 io_A_Valid_0_delay_25_20;
  reg                 io_A_Valid_0_delay_26_19;
  reg                 io_A_Valid_0_delay_27_18;
  reg                 io_A_Valid_0_delay_28_17;
  reg                 io_A_Valid_0_delay_29_16;
  reg                 io_A_Valid_0_delay_30_15;
  reg                 io_A_Valid_0_delay_31_14;
  reg                 io_A_Valid_0_delay_32_13;
  reg                 io_A_Valid_0_delay_33_12;
  reg                 io_A_Valid_0_delay_34_11;
  reg                 io_A_Valid_0_delay_35_10;
  reg                 io_A_Valid_0_delay_36_9;
  reg                 io_A_Valid_0_delay_37_8;
  reg                 io_A_Valid_0_delay_38_7;
  reg                 io_A_Valid_0_delay_39_6;
  reg                 io_A_Valid_0_delay_40_5;
  reg                 io_A_Valid_0_delay_41_4;
  reg                 io_A_Valid_0_delay_42_3;
  reg                 io_A_Valid_0_delay_43_2;
  reg                 io_A_Valid_0_delay_44_1;
  reg                 io_A_Valid_0_delay_45;
  reg                 io_A_Valid_0_delay_1_45;
  reg                 io_A_Valid_0_delay_2_44;
  reg                 io_A_Valid_0_delay_3_43;
  reg                 io_A_Valid_0_delay_4_42;
  reg                 io_A_Valid_0_delay_5_41;
  reg                 io_A_Valid_0_delay_6_40;
  reg                 io_A_Valid_0_delay_7_39;
  reg                 io_A_Valid_0_delay_8_38;
  reg                 io_A_Valid_0_delay_9_37;
  reg                 io_A_Valid_0_delay_10_36;
  reg                 io_A_Valid_0_delay_11_35;
  reg                 io_A_Valid_0_delay_12_34;
  reg                 io_A_Valid_0_delay_13_33;
  reg                 io_A_Valid_0_delay_14_32;
  reg                 io_A_Valid_0_delay_15_31;
  reg                 io_A_Valid_0_delay_16_30;
  reg                 io_A_Valid_0_delay_17_29;
  reg                 io_A_Valid_0_delay_18_28;
  reg                 io_A_Valid_0_delay_19_27;
  reg                 io_A_Valid_0_delay_20_26;
  reg                 io_A_Valid_0_delay_21_25;
  reg                 io_A_Valid_0_delay_22_24;
  reg                 io_A_Valid_0_delay_23_23;
  reg                 io_A_Valid_0_delay_24_22;
  reg                 io_A_Valid_0_delay_25_21;
  reg                 io_A_Valid_0_delay_26_20;
  reg                 io_A_Valid_0_delay_27_19;
  reg                 io_A_Valid_0_delay_28_18;
  reg                 io_A_Valid_0_delay_29_17;
  reg                 io_A_Valid_0_delay_30_16;
  reg                 io_A_Valid_0_delay_31_15;
  reg                 io_A_Valid_0_delay_32_14;
  reg                 io_A_Valid_0_delay_33_13;
  reg                 io_A_Valid_0_delay_34_12;
  reg                 io_A_Valid_0_delay_35_11;
  reg                 io_A_Valid_0_delay_36_10;
  reg                 io_A_Valid_0_delay_37_9;
  reg                 io_A_Valid_0_delay_38_8;
  reg                 io_A_Valid_0_delay_39_7;
  reg                 io_A_Valid_0_delay_40_6;
  reg                 io_A_Valid_0_delay_41_5;
  reg                 io_A_Valid_0_delay_42_4;
  reg                 io_A_Valid_0_delay_43_3;
  reg                 io_A_Valid_0_delay_44_2;
  reg                 io_A_Valid_0_delay_45_1;
  reg                 io_A_Valid_0_delay_46;
  reg                 io_A_Valid_0_delay_1_46;
  reg                 io_A_Valid_0_delay_2_45;
  reg                 io_A_Valid_0_delay_3_44;
  reg                 io_A_Valid_0_delay_4_43;
  reg                 io_A_Valid_0_delay_5_42;
  reg                 io_A_Valid_0_delay_6_41;
  reg                 io_A_Valid_0_delay_7_40;
  reg                 io_A_Valid_0_delay_8_39;
  reg                 io_A_Valid_0_delay_9_38;
  reg                 io_A_Valid_0_delay_10_37;
  reg                 io_A_Valid_0_delay_11_36;
  reg                 io_A_Valid_0_delay_12_35;
  reg                 io_A_Valid_0_delay_13_34;
  reg                 io_A_Valid_0_delay_14_33;
  reg                 io_A_Valid_0_delay_15_32;
  reg                 io_A_Valid_0_delay_16_31;
  reg                 io_A_Valid_0_delay_17_30;
  reg                 io_A_Valid_0_delay_18_29;
  reg                 io_A_Valid_0_delay_19_28;
  reg                 io_A_Valid_0_delay_20_27;
  reg                 io_A_Valid_0_delay_21_26;
  reg                 io_A_Valid_0_delay_22_25;
  reg                 io_A_Valid_0_delay_23_24;
  reg                 io_A_Valid_0_delay_24_23;
  reg                 io_A_Valid_0_delay_25_22;
  reg                 io_A_Valid_0_delay_26_21;
  reg                 io_A_Valid_0_delay_27_20;
  reg                 io_A_Valid_0_delay_28_19;
  reg                 io_A_Valid_0_delay_29_18;
  reg                 io_A_Valid_0_delay_30_17;
  reg                 io_A_Valid_0_delay_31_16;
  reg                 io_A_Valid_0_delay_32_15;
  reg                 io_A_Valid_0_delay_33_14;
  reg                 io_A_Valid_0_delay_34_13;
  reg                 io_A_Valid_0_delay_35_12;
  reg                 io_A_Valid_0_delay_36_11;
  reg                 io_A_Valid_0_delay_37_10;
  reg                 io_A_Valid_0_delay_38_9;
  reg                 io_A_Valid_0_delay_39_8;
  reg                 io_A_Valid_0_delay_40_7;
  reg                 io_A_Valid_0_delay_41_6;
  reg                 io_A_Valid_0_delay_42_5;
  reg                 io_A_Valid_0_delay_43_4;
  reg                 io_A_Valid_0_delay_44_3;
  reg                 io_A_Valid_0_delay_45_2;
  reg                 io_A_Valid_0_delay_46_1;
  reg                 io_A_Valid_0_delay_47;
  reg                 io_A_Valid_0_delay_1_47;
  reg                 io_A_Valid_0_delay_2_46;
  reg                 io_A_Valid_0_delay_3_45;
  reg                 io_A_Valid_0_delay_4_44;
  reg                 io_A_Valid_0_delay_5_43;
  reg                 io_A_Valid_0_delay_6_42;
  reg                 io_A_Valid_0_delay_7_41;
  reg                 io_A_Valid_0_delay_8_40;
  reg                 io_A_Valid_0_delay_9_39;
  reg                 io_A_Valid_0_delay_10_38;
  reg                 io_A_Valid_0_delay_11_37;
  reg                 io_A_Valid_0_delay_12_36;
  reg                 io_A_Valid_0_delay_13_35;
  reg                 io_A_Valid_0_delay_14_34;
  reg                 io_A_Valid_0_delay_15_33;
  reg                 io_A_Valid_0_delay_16_32;
  reg                 io_A_Valid_0_delay_17_31;
  reg                 io_A_Valid_0_delay_18_30;
  reg                 io_A_Valid_0_delay_19_29;
  reg                 io_A_Valid_0_delay_20_28;
  reg                 io_A_Valid_0_delay_21_27;
  reg                 io_A_Valid_0_delay_22_26;
  reg                 io_A_Valid_0_delay_23_25;
  reg                 io_A_Valid_0_delay_24_24;
  reg                 io_A_Valid_0_delay_25_23;
  reg                 io_A_Valid_0_delay_26_22;
  reg                 io_A_Valid_0_delay_27_21;
  reg                 io_A_Valid_0_delay_28_20;
  reg                 io_A_Valid_0_delay_29_19;
  reg                 io_A_Valid_0_delay_30_18;
  reg                 io_A_Valid_0_delay_31_17;
  reg                 io_A_Valid_0_delay_32_16;
  reg                 io_A_Valid_0_delay_33_15;
  reg                 io_A_Valid_0_delay_34_14;
  reg                 io_A_Valid_0_delay_35_13;
  reg                 io_A_Valid_0_delay_36_12;
  reg                 io_A_Valid_0_delay_37_11;
  reg                 io_A_Valid_0_delay_38_10;
  reg                 io_A_Valid_0_delay_39_9;
  reg                 io_A_Valid_0_delay_40_8;
  reg                 io_A_Valid_0_delay_41_7;
  reg                 io_A_Valid_0_delay_42_6;
  reg                 io_A_Valid_0_delay_43_5;
  reg                 io_A_Valid_0_delay_44_4;
  reg                 io_A_Valid_0_delay_45_3;
  reg                 io_A_Valid_0_delay_46_2;
  reg                 io_A_Valid_0_delay_47_1;
  reg                 io_A_Valid_0_delay_48;
  reg                 io_A_Valid_0_delay_1_48;
  reg                 io_A_Valid_0_delay_2_47;
  reg                 io_A_Valid_0_delay_3_46;
  reg                 io_A_Valid_0_delay_4_45;
  reg                 io_A_Valid_0_delay_5_44;
  reg                 io_A_Valid_0_delay_6_43;
  reg                 io_A_Valid_0_delay_7_42;
  reg                 io_A_Valid_0_delay_8_41;
  reg                 io_A_Valid_0_delay_9_40;
  reg                 io_A_Valid_0_delay_10_39;
  reg                 io_A_Valid_0_delay_11_38;
  reg                 io_A_Valid_0_delay_12_37;
  reg                 io_A_Valid_0_delay_13_36;
  reg                 io_A_Valid_0_delay_14_35;
  reg                 io_A_Valid_0_delay_15_34;
  reg                 io_A_Valid_0_delay_16_33;
  reg                 io_A_Valid_0_delay_17_32;
  reg                 io_A_Valid_0_delay_18_31;
  reg                 io_A_Valid_0_delay_19_30;
  reg                 io_A_Valid_0_delay_20_29;
  reg                 io_A_Valid_0_delay_21_28;
  reg                 io_A_Valid_0_delay_22_27;
  reg                 io_A_Valid_0_delay_23_26;
  reg                 io_A_Valid_0_delay_24_25;
  reg                 io_A_Valid_0_delay_25_24;
  reg                 io_A_Valid_0_delay_26_23;
  reg                 io_A_Valid_0_delay_27_22;
  reg                 io_A_Valid_0_delay_28_21;
  reg                 io_A_Valid_0_delay_29_20;
  reg                 io_A_Valid_0_delay_30_19;
  reg                 io_A_Valid_0_delay_31_18;
  reg                 io_A_Valid_0_delay_32_17;
  reg                 io_A_Valid_0_delay_33_16;
  reg                 io_A_Valid_0_delay_34_15;
  reg                 io_A_Valid_0_delay_35_14;
  reg                 io_A_Valid_0_delay_36_13;
  reg                 io_A_Valid_0_delay_37_12;
  reg                 io_A_Valid_0_delay_38_11;
  reg                 io_A_Valid_0_delay_39_10;
  reg                 io_A_Valid_0_delay_40_9;
  reg                 io_A_Valid_0_delay_41_8;
  reg                 io_A_Valid_0_delay_42_7;
  reg                 io_A_Valid_0_delay_43_6;
  reg                 io_A_Valid_0_delay_44_5;
  reg                 io_A_Valid_0_delay_45_4;
  reg                 io_A_Valid_0_delay_46_3;
  reg                 io_A_Valid_0_delay_47_2;
  reg                 io_A_Valid_0_delay_48_1;
  reg                 io_A_Valid_0_delay_49;
  reg                 io_A_Valid_0_delay_1_49;
  reg                 io_A_Valid_0_delay_2_48;
  reg                 io_A_Valid_0_delay_3_47;
  reg                 io_A_Valid_0_delay_4_46;
  reg                 io_A_Valid_0_delay_5_45;
  reg                 io_A_Valid_0_delay_6_44;
  reg                 io_A_Valid_0_delay_7_43;
  reg                 io_A_Valid_0_delay_8_42;
  reg                 io_A_Valid_0_delay_9_41;
  reg                 io_A_Valid_0_delay_10_40;
  reg                 io_A_Valid_0_delay_11_39;
  reg                 io_A_Valid_0_delay_12_38;
  reg                 io_A_Valid_0_delay_13_37;
  reg                 io_A_Valid_0_delay_14_36;
  reg                 io_A_Valid_0_delay_15_35;
  reg                 io_A_Valid_0_delay_16_34;
  reg                 io_A_Valid_0_delay_17_33;
  reg                 io_A_Valid_0_delay_18_32;
  reg                 io_A_Valid_0_delay_19_31;
  reg                 io_A_Valid_0_delay_20_30;
  reg                 io_A_Valid_0_delay_21_29;
  reg                 io_A_Valid_0_delay_22_28;
  reg                 io_A_Valid_0_delay_23_27;
  reg                 io_A_Valid_0_delay_24_26;
  reg                 io_A_Valid_0_delay_25_25;
  reg                 io_A_Valid_0_delay_26_24;
  reg                 io_A_Valid_0_delay_27_23;
  reg                 io_A_Valid_0_delay_28_22;
  reg                 io_A_Valid_0_delay_29_21;
  reg                 io_A_Valid_0_delay_30_20;
  reg                 io_A_Valid_0_delay_31_19;
  reg                 io_A_Valid_0_delay_32_18;
  reg                 io_A_Valid_0_delay_33_17;
  reg                 io_A_Valid_0_delay_34_16;
  reg                 io_A_Valid_0_delay_35_15;
  reg                 io_A_Valid_0_delay_36_14;
  reg                 io_A_Valid_0_delay_37_13;
  reg                 io_A_Valid_0_delay_38_12;
  reg                 io_A_Valid_0_delay_39_11;
  reg                 io_A_Valid_0_delay_40_10;
  reg                 io_A_Valid_0_delay_41_9;
  reg                 io_A_Valid_0_delay_42_8;
  reg                 io_A_Valid_0_delay_43_7;
  reg                 io_A_Valid_0_delay_44_6;
  reg                 io_A_Valid_0_delay_45_5;
  reg                 io_A_Valid_0_delay_46_4;
  reg                 io_A_Valid_0_delay_47_3;
  reg                 io_A_Valid_0_delay_48_2;
  reg                 io_A_Valid_0_delay_49_1;
  reg                 io_A_Valid_0_delay_50;
  reg                 io_A_Valid_0_delay_1_50;
  reg                 io_A_Valid_0_delay_2_49;
  reg                 io_A_Valid_0_delay_3_48;
  reg                 io_A_Valid_0_delay_4_47;
  reg                 io_A_Valid_0_delay_5_46;
  reg                 io_A_Valid_0_delay_6_45;
  reg                 io_A_Valid_0_delay_7_44;
  reg                 io_A_Valid_0_delay_8_43;
  reg                 io_A_Valid_0_delay_9_42;
  reg                 io_A_Valid_0_delay_10_41;
  reg                 io_A_Valid_0_delay_11_40;
  reg                 io_A_Valid_0_delay_12_39;
  reg                 io_A_Valid_0_delay_13_38;
  reg                 io_A_Valid_0_delay_14_37;
  reg                 io_A_Valid_0_delay_15_36;
  reg                 io_A_Valid_0_delay_16_35;
  reg                 io_A_Valid_0_delay_17_34;
  reg                 io_A_Valid_0_delay_18_33;
  reg                 io_A_Valid_0_delay_19_32;
  reg                 io_A_Valid_0_delay_20_31;
  reg                 io_A_Valid_0_delay_21_30;
  reg                 io_A_Valid_0_delay_22_29;
  reg                 io_A_Valid_0_delay_23_28;
  reg                 io_A_Valid_0_delay_24_27;
  reg                 io_A_Valid_0_delay_25_26;
  reg                 io_A_Valid_0_delay_26_25;
  reg                 io_A_Valid_0_delay_27_24;
  reg                 io_A_Valid_0_delay_28_23;
  reg                 io_A_Valid_0_delay_29_22;
  reg                 io_A_Valid_0_delay_30_21;
  reg                 io_A_Valid_0_delay_31_20;
  reg                 io_A_Valid_0_delay_32_19;
  reg                 io_A_Valid_0_delay_33_18;
  reg                 io_A_Valid_0_delay_34_17;
  reg                 io_A_Valid_0_delay_35_16;
  reg                 io_A_Valid_0_delay_36_15;
  reg                 io_A_Valid_0_delay_37_14;
  reg                 io_A_Valid_0_delay_38_13;
  reg                 io_A_Valid_0_delay_39_12;
  reg                 io_A_Valid_0_delay_40_11;
  reg                 io_A_Valid_0_delay_41_10;
  reg                 io_A_Valid_0_delay_42_9;
  reg                 io_A_Valid_0_delay_43_8;
  reg                 io_A_Valid_0_delay_44_7;
  reg                 io_A_Valid_0_delay_45_6;
  reg                 io_A_Valid_0_delay_46_5;
  reg                 io_A_Valid_0_delay_47_4;
  reg                 io_A_Valid_0_delay_48_3;
  reg                 io_A_Valid_0_delay_49_2;
  reg                 io_A_Valid_0_delay_50_1;
  reg                 io_A_Valid_0_delay_51;
  reg                 io_A_Valid_0_delay_1_51;
  reg                 io_A_Valid_0_delay_2_50;
  reg                 io_A_Valid_0_delay_3_49;
  reg                 io_A_Valid_0_delay_4_48;
  reg                 io_A_Valid_0_delay_5_47;
  reg                 io_A_Valid_0_delay_6_46;
  reg                 io_A_Valid_0_delay_7_45;
  reg                 io_A_Valid_0_delay_8_44;
  reg                 io_A_Valid_0_delay_9_43;
  reg                 io_A_Valid_0_delay_10_42;
  reg                 io_A_Valid_0_delay_11_41;
  reg                 io_A_Valid_0_delay_12_40;
  reg                 io_A_Valid_0_delay_13_39;
  reg                 io_A_Valid_0_delay_14_38;
  reg                 io_A_Valid_0_delay_15_37;
  reg                 io_A_Valid_0_delay_16_36;
  reg                 io_A_Valid_0_delay_17_35;
  reg                 io_A_Valid_0_delay_18_34;
  reg                 io_A_Valid_0_delay_19_33;
  reg                 io_A_Valid_0_delay_20_32;
  reg                 io_A_Valid_0_delay_21_31;
  reg                 io_A_Valid_0_delay_22_30;
  reg                 io_A_Valid_0_delay_23_29;
  reg                 io_A_Valid_0_delay_24_28;
  reg                 io_A_Valid_0_delay_25_27;
  reg                 io_A_Valid_0_delay_26_26;
  reg                 io_A_Valid_0_delay_27_25;
  reg                 io_A_Valid_0_delay_28_24;
  reg                 io_A_Valid_0_delay_29_23;
  reg                 io_A_Valid_0_delay_30_22;
  reg                 io_A_Valid_0_delay_31_21;
  reg                 io_A_Valid_0_delay_32_20;
  reg                 io_A_Valid_0_delay_33_19;
  reg                 io_A_Valid_0_delay_34_18;
  reg                 io_A_Valid_0_delay_35_17;
  reg                 io_A_Valid_0_delay_36_16;
  reg                 io_A_Valid_0_delay_37_15;
  reg                 io_A_Valid_0_delay_38_14;
  reg                 io_A_Valid_0_delay_39_13;
  reg                 io_A_Valid_0_delay_40_12;
  reg                 io_A_Valid_0_delay_41_11;
  reg                 io_A_Valid_0_delay_42_10;
  reg                 io_A_Valid_0_delay_43_9;
  reg                 io_A_Valid_0_delay_44_8;
  reg                 io_A_Valid_0_delay_45_7;
  reg                 io_A_Valid_0_delay_46_6;
  reg                 io_A_Valid_0_delay_47_5;
  reg                 io_A_Valid_0_delay_48_4;
  reg                 io_A_Valid_0_delay_49_3;
  reg                 io_A_Valid_0_delay_50_2;
  reg                 io_A_Valid_0_delay_51_1;
  reg                 io_A_Valid_0_delay_52;
  reg                 io_A_Valid_0_delay_1_52;
  reg                 io_A_Valid_0_delay_2_51;
  reg                 io_A_Valid_0_delay_3_50;
  reg                 io_A_Valid_0_delay_4_49;
  reg                 io_A_Valid_0_delay_5_48;
  reg                 io_A_Valid_0_delay_6_47;
  reg                 io_A_Valid_0_delay_7_46;
  reg                 io_A_Valid_0_delay_8_45;
  reg                 io_A_Valid_0_delay_9_44;
  reg                 io_A_Valid_0_delay_10_43;
  reg                 io_A_Valid_0_delay_11_42;
  reg                 io_A_Valid_0_delay_12_41;
  reg                 io_A_Valid_0_delay_13_40;
  reg                 io_A_Valid_0_delay_14_39;
  reg                 io_A_Valid_0_delay_15_38;
  reg                 io_A_Valid_0_delay_16_37;
  reg                 io_A_Valid_0_delay_17_36;
  reg                 io_A_Valid_0_delay_18_35;
  reg                 io_A_Valid_0_delay_19_34;
  reg                 io_A_Valid_0_delay_20_33;
  reg                 io_A_Valid_0_delay_21_32;
  reg                 io_A_Valid_0_delay_22_31;
  reg                 io_A_Valid_0_delay_23_30;
  reg                 io_A_Valid_0_delay_24_29;
  reg                 io_A_Valid_0_delay_25_28;
  reg                 io_A_Valid_0_delay_26_27;
  reg                 io_A_Valid_0_delay_27_26;
  reg                 io_A_Valid_0_delay_28_25;
  reg                 io_A_Valid_0_delay_29_24;
  reg                 io_A_Valid_0_delay_30_23;
  reg                 io_A_Valid_0_delay_31_22;
  reg                 io_A_Valid_0_delay_32_21;
  reg                 io_A_Valid_0_delay_33_20;
  reg                 io_A_Valid_0_delay_34_19;
  reg                 io_A_Valid_0_delay_35_18;
  reg                 io_A_Valid_0_delay_36_17;
  reg                 io_A_Valid_0_delay_37_16;
  reg                 io_A_Valid_0_delay_38_15;
  reg                 io_A_Valid_0_delay_39_14;
  reg                 io_A_Valid_0_delay_40_13;
  reg                 io_A_Valid_0_delay_41_12;
  reg                 io_A_Valid_0_delay_42_11;
  reg                 io_A_Valid_0_delay_43_10;
  reg                 io_A_Valid_0_delay_44_9;
  reg                 io_A_Valid_0_delay_45_8;
  reg                 io_A_Valid_0_delay_46_7;
  reg                 io_A_Valid_0_delay_47_6;
  reg                 io_A_Valid_0_delay_48_5;
  reg                 io_A_Valid_0_delay_49_4;
  reg                 io_A_Valid_0_delay_50_3;
  reg                 io_A_Valid_0_delay_51_2;
  reg                 io_A_Valid_0_delay_52_1;
  reg                 io_A_Valid_0_delay_53;
  reg                 io_A_Valid_0_delay_1_53;
  reg                 io_A_Valid_0_delay_2_52;
  reg                 io_A_Valid_0_delay_3_51;
  reg                 io_A_Valid_0_delay_4_50;
  reg                 io_A_Valid_0_delay_5_49;
  reg                 io_A_Valid_0_delay_6_48;
  reg                 io_A_Valid_0_delay_7_47;
  reg                 io_A_Valid_0_delay_8_46;
  reg                 io_A_Valid_0_delay_9_45;
  reg                 io_A_Valid_0_delay_10_44;
  reg                 io_A_Valid_0_delay_11_43;
  reg                 io_A_Valid_0_delay_12_42;
  reg                 io_A_Valid_0_delay_13_41;
  reg                 io_A_Valid_0_delay_14_40;
  reg                 io_A_Valid_0_delay_15_39;
  reg                 io_A_Valid_0_delay_16_38;
  reg                 io_A_Valid_0_delay_17_37;
  reg                 io_A_Valid_0_delay_18_36;
  reg                 io_A_Valid_0_delay_19_35;
  reg                 io_A_Valid_0_delay_20_34;
  reg                 io_A_Valid_0_delay_21_33;
  reg                 io_A_Valid_0_delay_22_32;
  reg                 io_A_Valid_0_delay_23_31;
  reg                 io_A_Valid_0_delay_24_30;
  reg                 io_A_Valid_0_delay_25_29;
  reg                 io_A_Valid_0_delay_26_28;
  reg                 io_A_Valid_0_delay_27_27;
  reg                 io_A_Valid_0_delay_28_26;
  reg                 io_A_Valid_0_delay_29_25;
  reg                 io_A_Valid_0_delay_30_24;
  reg                 io_A_Valid_0_delay_31_23;
  reg                 io_A_Valid_0_delay_32_22;
  reg                 io_A_Valid_0_delay_33_21;
  reg                 io_A_Valid_0_delay_34_20;
  reg                 io_A_Valid_0_delay_35_19;
  reg                 io_A_Valid_0_delay_36_18;
  reg                 io_A_Valid_0_delay_37_17;
  reg                 io_A_Valid_0_delay_38_16;
  reg                 io_A_Valid_0_delay_39_15;
  reg                 io_A_Valid_0_delay_40_14;
  reg                 io_A_Valid_0_delay_41_13;
  reg                 io_A_Valid_0_delay_42_12;
  reg                 io_A_Valid_0_delay_43_11;
  reg                 io_A_Valid_0_delay_44_10;
  reg                 io_A_Valid_0_delay_45_9;
  reg                 io_A_Valid_0_delay_46_8;
  reg                 io_A_Valid_0_delay_47_7;
  reg                 io_A_Valid_0_delay_48_6;
  reg                 io_A_Valid_0_delay_49_5;
  reg                 io_A_Valid_0_delay_50_4;
  reg                 io_A_Valid_0_delay_51_3;
  reg                 io_A_Valid_0_delay_52_2;
  reg                 io_A_Valid_0_delay_53_1;
  reg                 io_A_Valid_0_delay_54;
  reg                 io_A_Valid_0_delay_1_54;
  reg                 io_A_Valid_0_delay_2_53;
  reg                 io_A_Valid_0_delay_3_52;
  reg                 io_A_Valid_0_delay_4_51;
  reg                 io_A_Valid_0_delay_5_50;
  reg                 io_A_Valid_0_delay_6_49;
  reg                 io_A_Valid_0_delay_7_48;
  reg                 io_A_Valid_0_delay_8_47;
  reg                 io_A_Valid_0_delay_9_46;
  reg                 io_A_Valid_0_delay_10_45;
  reg                 io_A_Valid_0_delay_11_44;
  reg                 io_A_Valid_0_delay_12_43;
  reg                 io_A_Valid_0_delay_13_42;
  reg                 io_A_Valid_0_delay_14_41;
  reg                 io_A_Valid_0_delay_15_40;
  reg                 io_A_Valid_0_delay_16_39;
  reg                 io_A_Valid_0_delay_17_38;
  reg                 io_A_Valid_0_delay_18_37;
  reg                 io_A_Valid_0_delay_19_36;
  reg                 io_A_Valid_0_delay_20_35;
  reg                 io_A_Valid_0_delay_21_34;
  reg                 io_A_Valid_0_delay_22_33;
  reg                 io_A_Valid_0_delay_23_32;
  reg                 io_A_Valid_0_delay_24_31;
  reg                 io_A_Valid_0_delay_25_30;
  reg                 io_A_Valid_0_delay_26_29;
  reg                 io_A_Valid_0_delay_27_28;
  reg                 io_A_Valid_0_delay_28_27;
  reg                 io_A_Valid_0_delay_29_26;
  reg                 io_A_Valid_0_delay_30_25;
  reg                 io_A_Valid_0_delay_31_24;
  reg                 io_A_Valid_0_delay_32_23;
  reg                 io_A_Valid_0_delay_33_22;
  reg                 io_A_Valid_0_delay_34_21;
  reg                 io_A_Valid_0_delay_35_20;
  reg                 io_A_Valid_0_delay_36_19;
  reg                 io_A_Valid_0_delay_37_18;
  reg                 io_A_Valid_0_delay_38_17;
  reg                 io_A_Valid_0_delay_39_16;
  reg                 io_A_Valid_0_delay_40_15;
  reg                 io_A_Valid_0_delay_41_14;
  reg                 io_A_Valid_0_delay_42_13;
  reg                 io_A_Valid_0_delay_43_12;
  reg                 io_A_Valid_0_delay_44_11;
  reg                 io_A_Valid_0_delay_45_10;
  reg                 io_A_Valid_0_delay_46_9;
  reg                 io_A_Valid_0_delay_47_8;
  reg                 io_A_Valid_0_delay_48_7;
  reg                 io_A_Valid_0_delay_49_6;
  reg                 io_A_Valid_0_delay_50_5;
  reg                 io_A_Valid_0_delay_51_4;
  reg                 io_A_Valid_0_delay_52_3;
  reg                 io_A_Valid_0_delay_53_2;
  reg                 io_A_Valid_0_delay_54_1;
  reg                 io_A_Valid_0_delay_55;
  reg                 io_A_Valid_0_delay_1_55;
  reg                 io_A_Valid_0_delay_2_54;
  reg                 io_A_Valid_0_delay_3_53;
  reg                 io_A_Valid_0_delay_4_52;
  reg                 io_A_Valid_0_delay_5_51;
  reg                 io_A_Valid_0_delay_6_50;
  reg                 io_A_Valid_0_delay_7_49;
  reg                 io_A_Valid_0_delay_8_48;
  reg                 io_A_Valid_0_delay_9_47;
  reg                 io_A_Valid_0_delay_10_46;
  reg                 io_A_Valid_0_delay_11_45;
  reg                 io_A_Valid_0_delay_12_44;
  reg                 io_A_Valid_0_delay_13_43;
  reg                 io_A_Valid_0_delay_14_42;
  reg                 io_A_Valid_0_delay_15_41;
  reg                 io_A_Valid_0_delay_16_40;
  reg                 io_A_Valid_0_delay_17_39;
  reg                 io_A_Valid_0_delay_18_38;
  reg                 io_A_Valid_0_delay_19_37;
  reg                 io_A_Valid_0_delay_20_36;
  reg                 io_A_Valid_0_delay_21_35;
  reg                 io_A_Valid_0_delay_22_34;
  reg                 io_A_Valid_0_delay_23_33;
  reg                 io_A_Valid_0_delay_24_32;
  reg                 io_A_Valid_0_delay_25_31;
  reg                 io_A_Valid_0_delay_26_30;
  reg                 io_A_Valid_0_delay_27_29;
  reg                 io_A_Valid_0_delay_28_28;
  reg                 io_A_Valid_0_delay_29_27;
  reg                 io_A_Valid_0_delay_30_26;
  reg                 io_A_Valid_0_delay_31_25;
  reg                 io_A_Valid_0_delay_32_24;
  reg                 io_A_Valid_0_delay_33_23;
  reg                 io_A_Valid_0_delay_34_22;
  reg                 io_A_Valid_0_delay_35_21;
  reg                 io_A_Valid_0_delay_36_20;
  reg                 io_A_Valid_0_delay_37_19;
  reg                 io_A_Valid_0_delay_38_18;
  reg                 io_A_Valid_0_delay_39_17;
  reg                 io_A_Valid_0_delay_40_16;
  reg                 io_A_Valid_0_delay_41_15;
  reg                 io_A_Valid_0_delay_42_14;
  reg                 io_A_Valid_0_delay_43_13;
  reg                 io_A_Valid_0_delay_44_12;
  reg                 io_A_Valid_0_delay_45_11;
  reg                 io_A_Valid_0_delay_46_10;
  reg                 io_A_Valid_0_delay_47_9;
  reg                 io_A_Valid_0_delay_48_8;
  reg                 io_A_Valid_0_delay_49_7;
  reg                 io_A_Valid_0_delay_50_6;
  reg                 io_A_Valid_0_delay_51_5;
  reg                 io_A_Valid_0_delay_52_4;
  reg                 io_A_Valid_0_delay_53_3;
  reg                 io_A_Valid_0_delay_54_2;
  reg                 io_A_Valid_0_delay_55_1;
  reg                 io_A_Valid_0_delay_56;
  reg                 io_A_Valid_0_delay_1_56;
  reg                 io_A_Valid_0_delay_2_55;
  reg                 io_A_Valid_0_delay_3_54;
  reg                 io_A_Valid_0_delay_4_53;
  reg                 io_A_Valid_0_delay_5_52;
  reg                 io_A_Valid_0_delay_6_51;
  reg                 io_A_Valid_0_delay_7_50;
  reg                 io_A_Valid_0_delay_8_49;
  reg                 io_A_Valid_0_delay_9_48;
  reg                 io_A_Valid_0_delay_10_47;
  reg                 io_A_Valid_0_delay_11_46;
  reg                 io_A_Valid_0_delay_12_45;
  reg                 io_A_Valid_0_delay_13_44;
  reg                 io_A_Valid_0_delay_14_43;
  reg                 io_A_Valid_0_delay_15_42;
  reg                 io_A_Valid_0_delay_16_41;
  reg                 io_A_Valid_0_delay_17_40;
  reg                 io_A_Valid_0_delay_18_39;
  reg                 io_A_Valid_0_delay_19_38;
  reg                 io_A_Valid_0_delay_20_37;
  reg                 io_A_Valid_0_delay_21_36;
  reg                 io_A_Valid_0_delay_22_35;
  reg                 io_A_Valid_0_delay_23_34;
  reg                 io_A_Valid_0_delay_24_33;
  reg                 io_A_Valid_0_delay_25_32;
  reg                 io_A_Valid_0_delay_26_31;
  reg                 io_A_Valid_0_delay_27_30;
  reg                 io_A_Valid_0_delay_28_29;
  reg                 io_A_Valid_0_delay_29_28;
  reg                 io_A_Valid_0_delay_30_27;
  reg                 io_A_Valid_0_delay_31_26;
  reg                 io_A_Valid_0_delay_32_25;
  reg                 io_A_Valid_0_delay_33_24;
  reg                 io_A_Valid_0_delay_34_23;
  reg                 io_A_Valid_0_delay_35_22;
  reg                 io_A_Valid_0_delay_36_21;
  reg                 io_A_Valid_0_delay_37_20;
  reg                 io_A_Valid_0_delay_38_19;
  reg                 io_A_Valid_0_delay_39_18;
  reg                 io_A_Valid_0_delay_40_17;
  reg                 io_A_Valid_0_delay_41_16;
  reg                 io_A_Valid_0_delay_42_15;
  reg                 io_A_Valid_0_delay_43_14;
  reg                 io_A_Valid_0_delay_44_13;
  reg                 io_A_Valid_0_delay_45_12;
  reg                 io_A_Valid_0_delay_46_11;
  reg                 io_A_Valid_0_delay_47_10;
  reg                 io_A_Valid_0_delay_48_9;
  reg                 io_A_Valid_0_delay_49_8;
  reg                 io_A_Valid_0_delay_50_7;
  reg                 io_A_Valid_0_delay_51_6;
  reg                 io_A_Valid_0_delay_52_5;
  reg                 io_A_Valid_0_delay_53_4;
  reg                 io_A_Valid_0_delay_54_3;
  reg                 io_A_Valid_0_delay_55_2;
  reg                 io_A_Valid_0_delay_56_1;
  reg                 io_A_Valid_0_delay_57;
  reg                 io_A_Valid_0_delay_1_57;
  reg                 io_A_Valid_0_delay_2_56;
  reg                 io_A_Valid_0_delay_3_55;
  reg                 io_A_Valid_0_delay_4_54;
  reg                 io_A_Valid_0_delay_5_53;
  reg                 io_A_Valid_0_delay_6_52;
  reg                 io_A_Valid_0_delay_7_51;
  reg                 io_A_Valid_0_delay_8_50;
  reg                 io_A_Valid_0_delay_9_49;
  reg                 io_A_Valid_0_delay_10_48;
  reg                 io_A_Valid_0_delay_11_47;
  reg                 io_A_Valid_0_delay_12_46;
  reg                 io_A_Valid_0_delay_13_45;
  reg                 io_A_Valid_0_delay_14_44;
  reg                 io_A_Valid_0_delay_15_43;
  reg                 io_A_Valid_0_delay_16_42;
  reg                 io_A_Valid_0_delay_17_41;
  reg                 io_A_Valid_0_delay_18_40;
  reg                 io_A_Valid_0_delay_19_39;
  reg                 io_A_Valid_0_delay_20_38;
  reg                 io_A_Valid_0_delay_21_37;
  reg                 io_A_Valid_0_delay_22_36;
  reg                 io_A_Valid_0_delay_23_35;
  reg                 io_A_Valid_0_delay_24_34;
  reg                 io_A_Valid_0_delay_25_33;
  reg                 io_A_Valid_0_delay_26_32;
  reg                 io_A_Valid_0_delay_27_31;
  reg                 io_A_Valid_0_delay_28_30;
  reg                 io_A_Valid_0_delay_29_29;
  reg                 io_A_Valid_0_delay_30_28;
  reg                 io_A_Valid_0_delay_31_27;
  reg                 io_A_Valid_0_delay_32_26;
  reg                 io_A_Valid_0_delay_33_25;
  reg                 io_A_Valid_0_delay_34_24;
  reg                 io_A_Valid_0_delay_35_23;
  reg                 io_A_Valid_0_delay_36_22;
  reg                 io_A_Valid_0_delay_37_21;
  reg                 io_A_Valid_0_delay_38_20;
  reg                 io_A_Valid_0_delay_39_19;
  reg                 io_A_Valid_0_delay_40_18;
  reg                 io_A_Valid_0_delay_41_17;
  reg                 io_A_Valid_0_delay_42_16;
  reg                 io_A_Valid_0_delay_43_15;
  reg                 io_A_Valid_0_delay_44_14;
  reg                 io_A_Valid_0_delay_45_13;
  reg                 io_A_Valid_0_delay_46_12;
  reg                 io_A_Valid_0_delay_47_11;
  reg                 io_A_Valid_0_delay_48_10;
  reg                 io_A_Valid_0_delay_49_9;
  reg                 io_A_Valid_0_delay_50_8;
  reg                 io_A_Valid_0_delay_51_7;
  reg                 io_A_Valid_0_delay_52_6;
  reg                 io_A_Valid_0_delay_53_5;
  reg                 io_A_Valid_0_delay_54_4;
  reg                 io_A_Valid_0_delay_55_3;
  reg                 io_A_Valid_0_delay_56_2;
  reg                 io_A_Valid_0_delay_57_1;
  reg                 io_A_Valid_0_delay_58;
  reg                 io_A_Valid_0_delay_1_58;
  reg                 io_A_Valid_0_delay_2_57;
  reg                 io_A_Valid_0_delay_3_56;
  reg                 io_A_Valid_0_delay_4_55;
  reg                 io_A_Valid_0_delay_5_54;
  reg                 io_A_Valid_0_delay_6_53;
  reg                 io_A_Valid_0_delay_7_52;
  reg                 io_A_Valid_0_delay_8_51;
  reg                 io_A_Valid_0_delay_9_50;
  reg                 io_A_Valid_0_delay_10_49;
  reg                 io_A_Valid_0_delay_11_48;
  reg                 io_A_Valid_0_delay_12_47;
  reg                 io_A_Valid_0_delay_13_46;
  reg                 io_A_Valid_0_delay_14_45;
  reg                 io_A_Valid_0_delay_15_44;
  reg                 io_A_Valid_0_delay_16_43;
  reg                 io_A_Valid_0_delay_17_42;
  reg                 io_A_Valid_0_delay_18_41;
  reg                 io_A_Valid_0_delay_19_40;
  reg                 io_A_Valid_0_delay_20_39;
  reg                 io_A_Valid_0_delay_21_38;
  reg                 io_A_Valid_0_delay_22_37;
  reg                 io_A_Valid_0_delay_23_36;
  reg                 io_A_Valid_0_delay_24_35;
  reg                 io_A_Valid_0_delay_25_34;
  reg                 io_A_Valid_0_delay_26_33;
  reg                 io_A_Valid_0_delay_27_32;
  reg                 io_A_Valid_0_delay_28_31;
  reg                 io_A_Valid_0_delay_29_30;
  reg                 io_A_Valid_0_delay_30_29;
  reg                 io_A_Valid_0_delay_31_28;
  reg                 io_A_Valid_0_delay_32_27;
  reg                 io_A_Valid_0_delay_33_26;
  reg                 io_A_Valid_0_delay_34_25;
  reg                 io_A_Valid_0_delay_35_24;
  reg                 io_A_Valid_0_delay_36_23;
  reg                 io_A_Valid_0_delay_37_22;
  reg                 io_A_Valid_0_delay_38_21;
  reg                 io_A_Valid_0_delay_39_20;
  reg                 io_A_Valid_0_delay_40_19;
  reg                 io_A_Valid_0_delay_41_18;
  reg                 io_A_Valid_0_delay_42_17;
  reg                 io_A_Valid_0_delay_43_16;
  reg                 io_A_Valid_0_delay_44_15;
  reg                 io_A_Valid_0_delay_45_14;
  reg                 io_A_Valid_0_delay_46_13;
  reg                 io_A_Valid_0_delay_47_12;
  reg                 io_A_Valid_0_delay_48_11;
  reg                 io_A_Valid_0_delay_49_10;
  reg                 io_A_Valid_0_delay_50_9;
  reg                 io_A_Valid_0_delay_51_8;
  reg                 io_A_Valid_0_delay_52_7;
  reg                 io_A_Valid_0_delay_53_6;
  reg                 io_A_Valid_0_delay_54_5;
  reg                 io_A_Valid_0_delay_55_4;
  reg                 io_A_Valid_0_delay_56_3;
  reg                 io_A_Valid_0_delay_57_2;
  reg                 io_A_Valid_0_delay_58_1;
  reg                 io_A_Valid_0_delay_59;
  reg                 io_A_Valid_0_delay_1_59;
  reg                 io_A_Valid_0_delay_2_58;
  reg                 io_A_Valid_0_delay_3_57;
  reg                 io_A_Valid_0_delay_4_56;
  reg                 io_A_Valid_0_delay_5_55;
  reg                 io_A_Valid_0_delay_6_54;
  reg                 io_A_Valid_0_delay_7_53;
  reg                 io_A_Valid_0_delay_8_52;
  reg                 io_A_Valid_0_delay_9_51;
  reg                 io_A_Valid_0_delay_10_50;
  reg                 io_A_Valid_0_delay_11_49;
  reg                 io_A_Valid_0_delay_12_48;
  reg                 io_A_Valid_0_delay_13_47;
  reg                 io_A_Valid_0_delay_14_46;
  reg                 io_A_Valid_0_delay_15_45;
  reg                 io_A_Valid_0_delay_16_44;
  reg                 io_A_Valid_0_delay_17_43;
  reg                 io_A_Valid_0_delay_18_42;
  reg                 io_A_Valid_0_delay_19_41;
  reg                 io_A_Valid_0_delay_20_40;
  reg                 io_A_Valid_0_delay_21_39;
  reg                 io_A_Valid_0_delay_22_38;
  reg                 io_A_Valid_0_delay_23_37;
  reg                 io_A_Valid_0_delay_24_36;
  reg                 io_A_Valid_0_delay_25_35;
  reg                 io_A_Valid_0_delay_26_34;
  reg                 io_A_Valid_0_delay_27_33;
  reg                 io_A_Valid_0_delay_28_32;
  reg                 io_A_Valid_0_delay_29_31;
  reg                 io_A_Valid_0_delay_30_30;
  reg                 io_A_Valid_0_delay_31_29;
  reg                 io_A_Valid_0_delay_32_28;
  reg                 io_A_Valid_0_delay_33_27;
  reg                 io_A_Valid_0_delay_34_26;
  reg                 io_A_Valid_0_delay_35_25;
  reg                 io_A_Valid_0_delay_36_24;
  reg                 io_A_Valid_0_delay_37_23;
  reg                 io_A_Valid_0_delay_38_22;
  reg                 io_A_Valid_0_delay_39_21;
  reg                 io_A_Valid_0_delay_40_20;
  reg                 io_A_Valid_0_delay_41_19;
  reg                 io_A_Valid_0_delay_42_18;
  reg                 io_A_Valid_0_delay_43_17;
  reg                 io_A_Valid_0_delay_44_16;
  reg                 io_A_Valid_0_delay_45_15;
  reg                 io_A_Valid_0_delay_46_14;
  reg                 io_A_Valid_0_delay_47_13;
  reg                 io_A_Valid_0_delay_48_12;
  reg                 io_A_Valid_0_delay_49_11;
  reg                 io_A_Valid_0_delay_50_10;
  reg                 io_A_Valid_0_delay_51_9;
  reg                 io_A_Valid_0_delay_52_8;
  reg                 io_A_Valid_0_delay_53_7;
  reg                 io_A_Valid_0_delay_54_6;
  reg                 io_A_Valid_0_delay_55_5;
  reg                 io_A_Valid_0_delay_56_4;
  reg                 io_A_Valid_0_delay_57_3;
  reg                 io_A_Valid_0_delay_58_2;
  reg                 io_A_Valid_0_delay_59_1;
  reg                 io_A_Valid_0_delay_60;
  reg                 io_A_Valid_0_delay_1_60;
  reg                 io_A_Valid_0_delay_2_59;
  reg                 io_A_Valid_0_delay_3_58;
  reg                 io_A_Valid_0_delay_4_57;
  reg                 io_A_Valid_0_delay_5_56;
  reg                 io_A_Valid_0_delay_6_55;
  reg                 io_A_Valid_0_delay_7_54;
  reg                 io_A_Valid_0_delay_8_53;
  reg                 io_A_Valid_0_delay_9_52;
  reg                 io_A_Valid_0_delay_10_51;
  reg                 io_A_Valid_0_delay_11_50;
  reg                 io_A_Valid_0_delay_12_49;
  reg                 io_A_Valid_0_delay_13_48;
  reg                 io_A_Valid_0_delay_14_47;
  reg                 io_A_Valid_0_delay_15_46;
  reg                 io_A_Valid_0_delay_16_45;
  reg                 io_A_Valid_0_delay_17_44;
  reg                 io_A_Valid_0_delay_18_43;
  reg                 io_A_Valid_0_delay_19_42;
  reg                 io_A_Valid_0_delay_20_41;
  reg                 io_A_Valid_0_delay_21_40;
  reg                 io_A_Valid_0_delay_22_39;
  reg                 io_A_Valid_0_delay_23_38;
  reg                 io_A_Valid_0_delay_24_37;
  reg                 io_A_Valid_0_delay_25_36;
  reg                 io_A_Valid_0_delay_26_35;
  reg                 io_A_Valid_0_delay_27_34;
  reg                 io_A_Valid_0_delay_28_33;
  reg                 io_A_Valid_0_delay_29_32;
  reg                 io_A_Valid_0_delay_30_31;
  reg                 io_A_Valid_0_delay_31_30;
  reg                 io_A_Valid_0_delay_32_29;
  reg                 io_A_Valid_0_delay_33_28;
  reg                 io_A_Valid_0_delay_34_27;
  reg                 io_A_Valid_0_delay_35_26;
  reg                 io_A_Valid_0_delay_36_25;
  reg                 io_A_Valid_0_delay_37_24;
  reg                 io_A_Valid_0_delay_38_23;
  reg                 io_A_Valid_0_delay_39_22;
  reg                 io_A_Valid_0_delay_40_21;
  reg                 io_A_Valid_0_delay_41_20;
  reg                 io_A_Valid_0_delay_42_19;
  reg                 io_A_Valid_0_delay_43_18;
  reg                 io_A_Valid_0_delay_44_17;
  reg                 io_A_Valid_0_delay_45_16;
  reg                 io_A_Valid_0_delay_46_15;
  reg                 io_A_Valid_0_delay_47_14;
  reg                 io_A_Valid_0_delay_48_13;
  reg                 io_A_Valid_0_delay_49_12;
  reg                 io_A_Valid_0_delay_50_11;
  reg                 io_A_Valid_0_delay_51_10;
  reg                 io_A_Valid_0_delay_52_9;
  reg                 io_A_Valid_0_delay_53_8;
  reg                 io_A_Valid_0_delay_54_7;
  reg                 io_A_Valid_0_delay_55_6;
  reg                 io_A_Valid_0_delay_56_5;
  reg                 io_A_Valid_0_delay_57_4;
  reg                 io_A_Valid_0_delay_58_3;
  reg                 io_A_Valid_0_delay_59_2;
  reg                 io_A_Valid_0_delay_60_1;
  reg                 io_A_Valid_0_delay_61;
  reg                 io_A_Valid_0_delay_1_61;
  reg                 io_A_Valid_0_delay_2_60;
  reg                 io_A_Valid_0_delay_3_59;
  reg                 io_A_Valid_0_delay_4_58;
  reg                 io_A_Valid_0_delay_5_57;
  reg                 io_A_Valid_0_delay_6_56;
  reg                 io_A_Valid_0_delay_7_55;
  reg                 io_A_Valid_0_delay_8_54;
  reg                 io_A_Valid_0_delay_9_53;
  reg                 io_A_Valid_0_delay_10_52;
  reg                 io_A_Valid_0_delay_11_51;
  reg                 io_A_Valid_0_delay_12_50;
  reg                 io_A_Valid_0_delay_13_49;
  reg                 io_A_Valid_0_delay_14_48;
  reg                 io_A_Valid_0_delay_15_47;
  reg                 io_A_Valid_0_delay_16_46;
  reg                 io_A_Valid_0_delay_17_45;
  reg                 io_A_Valid_0_delay_18_44;
  reg                 io_A_Valid_0_delay_19_43;
  reg                 io_A_Valid_0_delay_20_42;
  reg                 io_A_Valid_0_delay_21_41;
  reg                 io_A_Valid_0_delay_22_40;
  reg                 io_A_Valid_0_delay_23_39;
  reg                 io_A_Valid_0_delay_24_38;
  reg                 io_A_Valid_0_delay_25_37;
  reg                 io_A_Valid_0_delay_26_36;
  reg                 io_A_Valid_0_delay_27_35;
  reg                 io_A_Valid_0_delay_28_34;
  reg                 io_A_Valid_0_delay_29_33;
  reg                 io_A_Valid_0_delay_30_32;
  reg                 io_A_Valid_0_delay_31_31;
  reg                 io_A_Valid_0_delay_32_30;
  reg                 io_A_Valid_0_delay_33_29;
  reg                 io_A_Valid_0_delay_34_28;
  reg                 io_A_Valid_0_delay_35_27;
  reg                 io_A_Valid_0_delay_36_26;
  reg                 io_A_Valid_0_delay_37_25;
  reg                 io_A_Valid_0_delay_38_24;
  reg                 io_A_Valid_0_delay_39_23;
  reg                 io_A_Valid_0_delay_40_22;
  reg                 io_A_Valid_0_delay_41_21;
  reg                 io_A_Valid_0_delay_42_20;
  reg                 io_A_Valid_0_delay_43_19;
  reg                 io_A_Valid_0_delay_44_18;
  reg                 io_A_Valid_0_delay_45_17;
  reg                 io_A_Valid_0_delay_46_16;
  reg                 io_A_Valid_0_delay_47_15;
  reg                 io_A_Valid_0_delay_48_14;
  reg                 io_A_Valid_0_delay_49_13;
  reg                 io_A_Valid_0_delay_50_12;
  reg                 io_A_Valid_0_delay_51_11;
  reg                 io_A_Valid_0_delay_52_10;
  reg                 io_A_Valid_0_delay_53_9;
  reg                 io_A_Valid_0_delay_54_8;
  reg                 io_A_Valid_0_delay_55_7;
  reg                 io_A_Valid_0_delay_56_6;
  reg                 io_A_Valid_0_delay_57_5;
  reg                 io_A_Valid_0_delay_58_4;
  reg                 io_A_Valid_0_delay_59_3;
  reg                 io_A_Valid_0_delay_60_2;
  reg                 io_A_Valid_0_delay_61_1;
  reg                 io_A_Valid_0_delay_62;
  reg                 io_A_Valid_0_delay_1_62;
  reg                 io_A_Valid_0_delay_2_61;
  reg                 io_A_Valid_0_delay_3_60;
  reg                 io_A_Valid_0_delay_4_59;
  reg                 io_A_Valid_0_delay_5_58;
  reg                 io_A_Valid_0_delay_6_57;
  reg                 io_A_Valid_0_delay_7_56;
  reg                 io_A_Valid_0_delay_8_55;
  reg                 io_A_Valid_0_delay_9_54;
  reg                 io_A_Valid_0_delay_10_53;
  reg                 io_A_Valid_0_delay_11_52;
  reg                 io_A_Valid_0_delay_12_51;
  reg                 io_A_Valid_0_delay_13_50;
  reg                 io_A_Valid_0_delay_14_49;
  reg                 io_A_Valid_0_delay_15_48;
  reg                 io_A_Valid_0_delay_16_47;
  reg                 io_A_Valid_0_delay_17_46;
  reg                 io_A_Valid_0_delay_18_45;
  reg                 io_A_Valid_0_delay_19_44;
  reg                 io_A_Valid_0_delay_20_43;
  reg                 io_A_Valid_0_delay_21_42;
  reg                 io_A_Valid_0_delay_22_41;
  reg                 io_A_Valid_0_delay_23_40;
  reg                 io_A_Valid_0_delay_24_39;
  reg                 io_A_Valid_0_delay_25_38;
  reg                 io_A_Valid_0_delay_26_37;
  reg                 io_A_Valid_0_delay_27_36;
  reg                 io_A_Valid_0_delay_28_35;
  reg                 io_A_Valid_0_delay_29_34;
  reg                 io_A_Valid_0_delay_30_33;
  reg                 io_A_Valid_0_delay_31_32;
  reg                 io_A_Valid_0_delay_32_31;
  reg                 io_A_Valid_0_delay_33_30;
  reg                 io_A_Valid_0_delay_34_29;
  reg                 io_A_Valid_0_delay_35_28;
  reg                 io_A_Valid_0_delay_36_27;
  reg                 io_A_Valid_0_delay_37_26;
  reg                 io_A_Valid_0_delay_38_25;
  reg                 io_A_Valid_0_delay_39_24;
  reg                 io_A_Valid_0_delay_40_23;
  reg                 io_A_Valid_0_delay_41_22;
  reg                 io_A_Valid_0_delay_42_21;
  reg                 io_A_Valid_0_delay_43_20;
  reg                 io_A_Valid_0_delay_44_19;
  reg                 io_A_Valid_0_delay_45_18;
  reg                 io_A_Valid_0_delay_46_17;
  reg                 io_A_Valid_0_delay_47_16;
  reg                 io_A_Valid_0_delay_48_15;
  reg                 io_A_Valid_0_delay_49_14;
  reg                 io_A_Valid_0_delay_50_13;
  reg                 io_A_Valid_0_delay_51_12;
  reg                 io_A_Valid_0_delay_52_11;
  reg                 io_A_Valid_0_delay_53_10;
  reg                 io_A_Valid_0_delay_54_9;
  reg                 io_A_Valid_0_delay_55_8;
  reg                 io_A_Valid_0_delay_56_7;
  reg                 io_A_Valid_0_delay_57_6;
  reg                 io_A_Valid_0_delay_58_5;
  reg                 io_A_Valid_0_delay_59_4;
  reg                 io_A_Valid_0_delay_60_3;
  reg                 io_A_Valid_0_delay_61_2;
  reg                 io_A_Valid_0_delay_62_1;
  reg                 io_A_Valid_0_delay_63;
  reg        [15:0]   io_signCount_regNextWhen_1;
  reg                 io_B_Valid_0_delay_1;
  reg                 io_A_Valid_1_delay_1;
  reg                 io_B_Valid_1_delay_1;
  reg                 io_A_Valid_1_delay_1_1;
  reg                 io_A_Valid_1_delay_2;
  reg                 io_B_Valid_2_delay_1;
  reg                 io_A_Valid_1_delay_1_2;
  reg                 io_A_Valid_1_delay_2_1;
  reg                 io_A_Valid_1_delay_3;
  reg                 io_B_Valid_3_delay_1;
  reg                 io_A_Valid_1_delay_1_3;
  reg                 io_A_Valid_1_delay_2_2;
  reg                 io_A_Valid_1_delay_3_1;
  reg                 io_A_Valid_1_delay_4;
  reg                 io_B_Valid_4_delay_1;
  reg                 io_A_Valid_1_delay_1_4;
  reg                 io_A_Valid_1_delay_2_3;
  reg                 io_A_Valid_1_delay_3_2;
  reg                 io_A_Valid_1_delay_4_1;
  reg                 io_A_Valid_1_delay_5;
  reg                 io_B_Valid_5_delay_1;
  reg                 io_A_Valid_1_delay_1_5;
  reg                 io_A_Valid_1_delay_2_4;
  reg                 io_A_Valid_1_delay_3_3;
  reg                 io_A_Valid_1_delay_4_2;
  reg                 io_A_Valid_1_delay_5_1;
  reg                 io_A_Valid_1_delay_6;
  reg                 io_B_Valid_6_delay_1;
  reg                 io_A_Valid_1_delay_1_6;
  reg                 io_A_Valid_1_delay_2_5;
  reg                 io_A_Valid_1_delay_3_4;
  reg                 io_A_Valid_1_delay_4_3;
  reg                 io_A_Valid_1_delay_5_2;
  reg                 io_A_Valid_1_delay_6_1;
  reg                 io_A_Valid_1_delay_7;
  reg                 io_B_Valid_7_delay_1;
  reg                 io_A_Valid_1_delay_1_7;
  reg                 io_A_Valid_1_delay_2_6;
  reg                 io_A_Valid_1_delay_3_5;
  reg                 io_A_Valid_1_delay_4_4;
  reg                 io_A_Valid_1_delay_5_3;
  reg                 io_A_Valid_1_delay_6_2;
  reg                 io_A_Valid_1_delay_7_1;
  reg                 io_A_Valid_1_delay_8;
  reg                 io_B_Valid_8_delay_1;
  reg                 io_A_Valid_1_delay_1_8;
  reg                 io_A_Valid_1_delay_2_7;
  reg                 io_A_Valid_1_delay_3_6;
  reg                 io_A_Valid_1_delay_4_5;
  reg                 io_A_Valid_1_delay_5_4;
  reg                 io_A_Valid_1_delay_6_3;
  reg                 io_A_Valid_1_delay_7_2;
  reg                 io_A_Valid_1_delay_8_1;
  reg                 io_A_Valid_1_delay_9;
  reg                 io_B_Valid_9_delay_1;
  reg                 io_A_Valid_1_delay_1_9;
  reg                 io_A_Valid_1_delay_2_8;
  reg                 io_A_Valid_1_delay_3_7;
  reg                 io_A_Valid_1_delay_4_6;
  reg                 io_A_Valid_1_delay_5_5;
  reg                 io_A_Valid_1_delay_6_4;
  reg                 io_A_Valid_1_delay_7_3;
  reg                 io_A_Valid_1_delay_8_2;
  reg                 io_A_Valid_1_delay_9_1;
  reg                 io_A_Valid_1_delay_10;
  reg                 io_B_Valid_10_delay_1;
  reg                 io_A_Valid_1_delay_1_10;
  reg                 io_A_Valid_1_delay_2_9;
  reg                 io_A_Valid_1_delay_3_8;
  reg                 io_A_Valid_1_delay_4_7;
  reg                 io_A_Valid_1_delay_5_6;
  reg                 io_A_Valid_1_delay_6_5;
  reg                 io_A_Valid_1_delay_7_4;
  reg                 io_A_Valid_1_delay_8_3;
  reg                 io_A_Valid_1_delay_9_2;
  reg                 io_A_Valid_1_delay_10_1;
  reg                 io_A_Valid_1_delay_11;
  reg                 io_B_Valid_11_delay_1;
  reg                 io_A_Valid_1_delay_1_11;
  reg                 io_A_Valid_1_delay_2_10;
  reg                 io_A_Valid_1_delay_3_9;
  reg                 io_A_Valid_1_delay_4_8;
  reg                 io_A_Valid_1_delay_5_7;
  reg                 io_A_Valid_1_delay_6_6;
  reg                 io_A_Valid_1_delay_7_5;
  reg                 io_A_Valid_1_delay_8_4;
  reg                 io_A_Valid_1_delay_9_3;
  reg                 io_A_Valid_1_delay_10_2;
  reg                 io_A_Valid_1_delay_11_1;
  reg                 io_A_Valid_1_delay_12;
  reg                 io_B_Valid_12_delay_1;
  reg                 io_A_Valid_1_delay_1_12;
  reg                 io_A_Valid_1_delay_2_11;
  reg                 io_A_Valid_1_delay_3_10;
  reg                 io_A_Valid_1_delay_4_9;
  reg                 io_A_Valid_1_delay_5_8;
  reg                 io_A_Valid_1_delay_6_7;
  reg                 io_A_Valid_1_delay_7_6;
  reg                 io_A_Valid_1_delay_8_5;
  reg                 io_A_Valid_1_delay_9_4;
  reg                 io_A_Valid_1_delay_10_3;
  reg                 io_A_Valid_1_delay_11_2;
  reg                 io_A_Valid_1_delay_12_1;
  reg                 io_A_Valid_1_delay_13;
  reg                 io_B_Valid_13_delay_1;
  reg                 io_A_Valid_1_delay_1_13;
  reg                 io_A_Valid_1_delay_2_12;
  reg                 io_A_Valid_1_delay_3_11;
  reg                 io_A_Valid_1_delay_4_10;
  reg                 io_A_Valid_1_delay_5_9;
  reg                 io_A_Valid_1_delay_6_8;
  reg                 io_A_Valid_1_delay_7_7;
  reg                 io_A_Valid_1_delay_8_6;
  reg                 io_A_Valid_1_delay_9_5;
  reg                 io_A_Valid_1_delay_10_4;
  reg                 io_A_Valid_1_delay_11_3;
  reg                 io_A_Valid_1_delay_12_2;
  reg                 io_A_Valid_1_delay_13_1;
  reg                 io_A_Valid_1_delay_14;
  reg                 io_B_Valid_14_delay_1;
  reg                 io_A_Valid_1_delay_1_14;
  reg                 io_A_Valid_1_delay_2_13;
  reg                 io_A_Valid_1_delay_3_12;
  reg                 io_A_Valid_1_delay_4_11;
  reg                 io_A_Valid_1_delay_5_10;
  reg                 io_A_Valid_1_delay_6_9;
  reg                 io_A_Valid_1_delay_7_8;
  reg                 io_A_Valid_1_delay_8_7;
  reg                 io_A_Valid_1_delay_9_6;
  reg                 io_A_Valid_1_delay_10_5;
  reg                 io_A_Valid_1_delay_11_4;
  reg                 io_A_Valid_1_delay_12_3;
  reg                 io_A_Valid_1_delay_13_2;
  reg                 io_A_Valid_1_delay_14_1;
  reg                 io_A_Valid_1_delay_15;
  reg                 io_B_Valid_15_delay_1;
  reg                 io_A_Valid_1_delay_1_15;
  reg                 io_A_Valid_1_delay_2_14;
  reg                 io_A_Valid_1_delay_3_13;
  reg                 io_A_Valid_1_delay_4_12;
  reg                 io_A_Valid_1_delay_5_11;
  reg                 io_A_Valid_1_delay_6_10;
  reg                 io_A_Valid_1_delay_7_9;
  reg                 io_A_Valid_1_delay_8_8;
  reg                 io_A_Valid_1_delay_9_7;
  reg                 io_A_Valid_1_delay_10_6;
  reg                 io_A_Valid_1_delay_11_5;
  reg                 io_A_Valid_1_delay_12_4;
  reg                 io_A_Valid_1_delay_13_3;
  reg                 io_A_Valid_1_delay_14_2;
  reg                 io_A_Valid_1_delay_15_1;
  reg                 io_A_Valid_1_delay_16;
  reg                 io_B_Valid_16_delay_1;
  reg                 io_A_Valid_1_delay_1_16;
  reg                 io_A_Valid_1_delay_2_15;
  reg                 io_A_Valid_1_delay_3_14;
  reg                 io_A_Valid_1_delay_4_13;
  reg                 io_A_Valid_1_delay_5_12;
  reg                 io_A_Valid_1_delay_6_11;
  reg                 io_A_Valid_1_delay_7_10;
  reg                 io_A_Valid_1_delay_8_9;
  reg                 io_A_Valid_1_delay_9_8;
  reg                 io_A_Valid_1_delay_10_7;
  reg                 io_A_Valid_1_delay_11_6;
  reg                 io_A_Valid_1_delay_12_5;
  reg                 io_A_Valid_1_delay_13_4;
  reg                 io_A_Valid_1_delay_14_3;
  reg                 io_A_Valid_1_delay_15_2;
  reg                 io_A_Valid_1_delay_16_1;
  reg                 io_A_Valid_1_delay_17;
  reg                 io_B_Valid_17_delay_1;
  reg                 io_A_Valid_1_delay_1_17;
  reg                 io_A_Valid_1_delay_2_16;
  reg                 io_A_Valid_1_delay_3_15;
  reg                 io_A_Valid_1_delay_4_14;
  reg                 io_A_Valid_1_delay_5_13;
  reg                 io_A_Valid_1_delay_6_12;
  reg                 io_A_Valid_1_delay_7_11;
  reg                 io_A_Valid_1_delay_8_10;
  reg                 io_A_Valid_1_delay_9_9;
  reg                 io_A_Valid_1_delay_10_8;
  reg                 io_A_Valid_1_delay_11_7;
  reg                 io_A_Valid_1_delay_12_6;
  reg                 io_A_Valid_1_delay_13_5;
  reg                 io_A_Valid_1_delay_14_4;
  reg                 io_A_Valid_1_delay_15_3;
  reg                 io_A_Valid_1_delay_16_2;
  reg                 io_A_Valid_1_delay_17_1;
  reg                 io_A_Valid_1_delay_18;
  reg                 io_B_Valid_18_delay_1;
  reg                 io_A_Valid_1_delay_1_18;
  reg                 io_A_Valid_1_delay_2_17;
  reg                 io_A_Valid_1_delay_3_16;
  reg                 io_A_Valid_1_delay_4_15;
  reg                 io_A_Valid_1_delay_5_14;
  reg                 io_A_Valid_1_delay_6_13;
  reg                 io_A_Valid_1_delay_7_12;
  reg                 io_A_Valid_1_delay_8_11;
  reg                 io_A_Valid_1_delay_9_10;
  reg                 io_A_Valid_1_delay_10_9;
  reg                 io_A_Valid_1_delay_11_8;
  reg                 io_A_Valid_1_delay_12_7;
  reg                 io_A_Valid_1_delay_13_6;
  reg                 io_A_Valid_1_delay_14_5;
  reg                 io_A_Valid_1_delay_15_4;
  reg                 io_A_Valid_1_delay_16_3;
  reg                 io_A_Valid_1_delay_17_2;
  reg                 io_A_Valid_1_delay_18_1;
  reg                 io_A_Valid_1_delay_19;
  reg                 io_B_Valid_19_delay_1;
  reg                 io_A_Valid_1_delay_1_19;
  reg                 io_A_Valid_1_delay_2_18;
  reg                 io_A_Valid_1_delay_3_17;
  reg                 io_A_Valid_1_delay_4_16;
  reg                 io_A_Valid_1_delay_5_15;
  reg                 io_A_Valid_1_delay_6_14;
  reg                 io_A_Valid_1_delay_7_13;
  reg                 io_A_Valid_1_delay_8_12;
  reg                 io_A_Valid_1_delay_9_11;
  reg                 io_A_Valid_1_delay_10_10;
  reg                 io_A_Valid_1_delay_11_9;
  reg                 io_A_Valid_1_delay_12_8;
  reg                 io_A_Valid_1_delay_13_7;
  reg                 io_A_Valid_1_delay_14_6;
  reg                 io_A_Valid_1_delay_15_5;
  reg                 io_A_Valid_1_delay_16_4;
  reg                 io_A_Valid_1_delay_17_3;
  reg                 io_A_Valid_1_delay_18_2;
  reg                 io_A_Valid_1_delay_19_1;
  reg                 io_A_Valid_1_delay_20;
  reg                 io_B_Valid_20_delay_1;
  reg                 io_A_Valid_1_delay_1_20;
  reg                 io_A_Valid_1_delay_2_19;
  reg                 io_A_Valid_1_delay_3_18;
  reg                 io_A_Valid_1_delay_4_17;
  reg                 io_A_Valid_1_delay_5_16;
  reg                 io_A_Valid_1_delay_6_15;
  reg                 io_A_Valid_1_delay_7_14;
  reg                 io_A_Valid_1_delay_8_13;
  reg                 io_A_Valid_1_delay_9_12;
  reg                 io_A_Valid_1_delay_10_11;
  reg                 io_A_Valid_1_delay_11_10;
  reg                 io_A_Valid_1_delay_12_9;
  reg                 io_A_Valid_1_delay_13_8;
  reg                 io_A_Valid_1_delay_14_7;
  reg                 io_A_Valid_1_delay_15_6;
  reg                 io_A_Valid_1_delay_16_5;
  reg                 io_A_Valid_1_delay_17_4;
  reg                 io_A_Valid_1_delay_18_3;
  reg                 io_A_Valid_1_delay_19_2;
  reg                 io_A_Valid_1_delay_20_1;
  reg                 io_A_Valid_1_delay_21;
  reg                 io_B_Valid_21_delay_1;
  reg                 io_A_Valid_1_delay_1_21;
  reg                 io_A_Valid_1_delay_2_20;
  reg                 io_A_Valid_1_delay_3_19;
  reg                 io_A_Valid_1_delay_4_18;
  reg                 io_A_Valid_1_delay_5_17;
  reg                 io_A_Valid_1_delay_6_16;
  reg                 io_A_Valid_1_delay_7_15;
  reg                 io_A_Valid_1_delay_8_14;
  reg                 io_A_Valid_1_delay_9_13;
  reg                 io_A_Valid_1_delay_10_12;
  reg                 io_A_Valid_1_delay_11_11;
  reg                 io_A_Valid_1_delay_12_10;
  reg                 io_A_Valid_1_delay_13_9;
  reg                 io_A_Valid_1_delay_14_8;
  reg                 io_A_Valid_1_delay_15_7;
  reg                 io_A_Valid_1_delay_16_6;
  reg                 io_A_Valid_1_delay_17_5;
  reg                 io_A_Valid_1_delay_18_4;
  reg                 io_A_Valid_1_delay_19_3;
  reg                 io_A_Valid_1_delay_20_2;
  reg                 io_A_Valid_1_delay_21_1;
  reg                 io_A_Valid_1_delay_22;
  reg                 io_B_Valid_22_delay_1;
  reg                 io_A_Valid_1_delay_1_22;
  reg                 io_A_Valid_1_delay_2_21;
  reg                 io_A_Valid_1_delay_3_20;
  reg                 io_A_Valid_1_delay_4_19;
  reg                 io_A_Valid_1_delay_5_18;
  reg                 io_A_Valid_1_delay_6_17;
  reg                 io_A_Valid_1_delay_7_16;
  reg                 io_A_Valid_1_delay_8_15;
  reg                 io_A_Valid_1_delay_9_14;
  reg                 io_A_Valid_1_delay_10_13;
  reg                 io_A_Valid_1_delay_11_12;
  reg                 io_A_Valid_1_delay_12_11;
  reg                 io_A_Valid_1_delay_13_10;
  reg                 io_A_Valid_1_delay_14_9;
  reg                 io_A_Valid_1_delay_15_8;
  reg                 io_A_Valid_1_delay_16_7;
  reg                 io_A_Valid_1_delay_17_6;
  reg                 io_A_Valid_1_delay_18_5;
  reg                 io_A_Valid_1_delay_19_4;
  reg                 io_A_Valid_1_delay_20_3;
  reg                 io_A_Valid_1_delay_21_2;
  reg                 io_A_Valid_1_delay_22_1;
  reg                 io_A_Valid_1_delay_23;
  reg                 io_B_Valid_23_delay_1;
  reg                 io_A_Valid_1_delay_1_23;
  reg                 io_A_Valid_1_delay_2_22;
  reg                 io_A_Valid_1_delay_3_21;
  reg                 io_A_Valid_1_delay_4_20;
  reg                 io_A_Valid_1_delay_5_19;
  reg                 io_A_Valid_1_delay_6_18;
  reg                 io_A_Valid_1_delay_7_17;
  reg                 io_A_Valid_1_delay_8_16;
  reg                 io_A_Valid_1_delay_9_15;
  reg                 io_A_Valid_1_delay_10_14;
  reg                 io_A_Valid_1_delay_11_13;
  reg                 io_A_Valid_1_delay_12_12;
  reg                 io_A_Valid_1_delay_13_11;
  reg                 io_A_Valid_1_delay_14_10;
  reg                 io_A_Valid_1_delay_15_9;
  reg                 io_A_Valid_1_delay_16_8;
  reg                 io_A_Valid_1_delay_17_7;
  reg                 io_A_Valid_1_delay_18_6;
  reg                 io_A_Valid_1_delay_19_5;
  reg                 io_A_Valid_1_delay_20_4;
  reg                 io_A_Valid_1_delay_21_3;
  reg                 io_A_Valid_1_delay_22_2;
  reg                 io_A_Valid_1_delay_23_1;
  reg                 io_A_Valid_1_delay_24;
  reg                 io_B_Valid_24_delay_1;
  reg                 io_A_Valid_1_delay_1_24;
  reg                 io_A_Valid_1_delay_2_23;
  reg                 io_A_Valid_1_delay_3_22;
  reg                 io_A_Valid_1_delay_4_21;
  reg                 io_A_Valid_1_delay_5_20;
  reg                 io_A_Valid_1_delay_6_19;
  reg                 io_A_Valid_1_delay_7_18;
  reg                 io_A_Valid_1_delay_8_17;
  reg                 io_A_Valid_1_delay_9_16;
  reg                 io_A_Valid_1_delay_10_15;
  reg                 io_A_Valid_1_delay_11_14;
  reg                 io_A_Valid_1_delay_12_13;
  reg                 io_A_Valid_1_delay_13_12;
  reg                 io_A_Valid_1_delay_14_11;
  reg                 io_A_Valid_1_delay_15_10;
  reg                 io_A_Valid_1_delay_16_9;
  reg                 io_A_Valid_1_delay_17_8;
  reg                 io_A_Valid_1_delay_18_7;
  reg                 io_A_Valid_1_delay_19_6;
  reg                 io_A_Valid_1_delay_20_5;
  reg                 io_A_Valid_1_delay_21_4;
  reg                 io_A_Valid_1_delay_22_3;
  reg                 io_A_Valid_1_delay_23_2;
  reg                 io_A_Valid_1_delay_24_1;
  reg                 io_A_Valid_1_delay_25;
  reg                 io_B_Valid_25_delay_1;
  reg                 io_A_Valid_1_delay_1_25;
  reg                 io_A_Valid_1_delay_2_24;
  reg                 io_A_Valid_1_delay_3_23;
  reg                 io_A_Valid_1_delay_4_22;
  reg                 io_A_Valid_1_delay_5_21;
  reg                 io_A_Valid_1_delay_6_20;
  reg                 io_A_Valid_1_delay_7_19;
  reg                 io_A_Valid_1_delay_8_18;
  reg                 io_A_Valid_1_delay_9_17;
  reg                 io_A_Valid_1_delay_10_16;
  reg                 io_A_Valid_1_delay_11_15;
  reg                 io_A_Valid_1_delay_12_14;
  reg                 io_A_Valid_1_delay_13_13;
  reg                 io_A_Valid_1_delay_14_12;
  reg                 io_A_Valid_1_delay_15_11;
  reg                 io_A_Valid_1_delay_16_10;
  reg                 io_A_Valid_1_delay_17_9;
  reg                 io_A_Valid_1_delay_18_8;
  reg                 io_A_Valid_1_delay_19_7;
  reg                 io_A_Valid_1_delay_20_6;
  reg                 io_A_Valid_1_delay_21_5;
  reg                 io_A_Valid_1_delay_22_4;
  reg                 io_A_Valid_1_delay_23_3;
  reg                 io_A_Valid_1_delay_24_2;
  reg                 io_A_Valid_1_delay_25_1;
  reg                 io_A_Valid_1_delay_26;
  reg                 io_B_Valid_26_delay_1;
  reg                 io_A_Valid_1_delay_1_26;
  reg                 io_A_Valid_1_delay_2_25;
  reg                 io_A_Valid_1_delay_3_24;
  reg                 io_A_Valid_1_delay_4_23;
  reg                 io_A_Valid_1_delay_5_22;
  reg                 io_A_Valid_1_delay_6_21;
  reg                 io_A_Valid_1_delay_7_20;
  reg                 io_A_Valid_1_delay_8_19;
  reg                 io_A_Valid_1_delay_9_18;
  reg                 io_A_Valid_1_delay_10_17;
  reg                 io_A_Valid_1_delay_11_16;
  reg                 io_A_Valid_1_delay_12_15;
  reg                 io_A_Valid_1_delay_13_14;
  reg                 io_A_Valid_1_delay_14_13;
  reg                 io_A_Valid_1_delay_15_12;
  reg                 io_A_Valid_1_delay_16_11;
  reg                 io_A_Valid_1_delay_17_10;
  reg                 io_A_Valid_1_delay_18_9;
  reg                 io_A_Valid_1_delay_19_8;
  reg                 io_A_Valid_1_delay_20_7;
  reg                 io_A_Valid_1_delay_21_6;
  reg                 io_A_Valid_1_delay_22_5;
  reg                 io_A_Valid_1_delay_23_4;
  reg                 io_A_Valid_1_delay_24_3;
  reg                 io_A_Valid_1_delay_25_2;
  reg                 io_A_Valid_1_delay_26_1;
  reg                 io_A_Valid_1_delay_27;
  reg                 io_B_Valid_27_delay_1;
  reg                 io_A_Valid_1_delay_1_27;
  reg                 io_A_Valid_1_delay_2_26;
  reg                 io_A_Valid_1_delay_3_25;
  reg                 io_A_Valid_1_delay_4_24;
  reg                 io_A_Valid_1_delay_5_23;
  reg                 io_A_Valid_1_delay_6_22;
  reg                 io_A_Valid_1_delay_7_21;
  reg                 io_A_Valid_1_delay_8_20;
  reg                 io_A_Valid_1_delay_9_19;
  reg                 io_A_Valid_1_delay_10_18;
  reg                 io_A_Valid_1_delay_11_17;
  reg                 io_A_Valid_1_delay_12_16;
  reg                 io_A_Valid_1_delay_13_15;
  reg                 io_A_Valid_1_delay_14_14;
  reg                 io_A_Valid_1_delay_15_13;
  reg                 io_A_Valid_1_delay_16_12;
  reg                 io_A_Valid_1_delay_17_11;
  reg                 io_A_Valid_1_delay_18_10;
  reg                 io_A_Valid_1_delay_19_9;
  reg                 io_A_Valid_1_delay_20_8;
  reg                 io_A_Valid_1_delay_21_7;
  reg                 io_A_Valid_1_delay_22_6;
  reg                 io_A_Valid_1_delay_23_5;
  reg                 io_A_Valid_1_delay_24_4;
  reg                 io_A_Valid_1_delay_25_3;
  reg                 io_A_Valid_1_delay_26_2;
  reg                 io_A_Valid_1_delay_27_1;
  reg                 io_A_Valid_1_delay_28;
  reg                 io_B_Valid_28_delay_1;
  reg                 io_A_Valid_1_delay_1_28;
  reg                 io_A_Valid_1_delay_2_27;
  reg                 io_A_Valid_1_delay_3_26;
  reg                 io_A_Valid_1_delay_4_25;
  reg                 io_A_Valid_1_delay_5_24;
  reg                 io_A_Valid_1_delay_6_23;
  reg                 io_A_Valid_1_delay_7_22;
  reg                 io_A_Valid_1_delay_8_21;
  reg                 io_A_Valid_1_delay_9_20;
  reg                 io_A_Valid_1_delay_10_19;
  reg                 io_A_Valid_1_delay_11_18;
  reg                 io_A_Valid_1_delay_12_17;
  reg                 io_A_Valid_1_delay_13_16;
  reg                 io_A_Valid_1_delay_14_15;
  reg                 io_A_Valid_1_delay_15_14;
  reg                 io_A_Valid_1_delay_16_13;
  reg                 io_A_Valid_1_delay_17_12;
  reg                 io_A_Valid_1_delay_18_11;
  reg                 io_A_Valid_1_delay_19_10;
  reg                 io_A_Valid_1_delay_20_9;
  reg                 io_A_Valid_1_delay_21_8;
  reg                 io_A_Valid_1_delay_22_7;
  reg                 io_A_Valid_1_delay_23_6;
  reg                 io_A_Valid_1_delay_24_5;
  reg                 io_A_Valid_1_delay_25_4;
  reg                 io_A_Valid_1_delay_26_3;
  reg                 io_A_Valid_1_delay_27_2;
  reg                 io_A_Valid_1_delay_28_1;
  reg                 io_A_Valid_1_delay_29;
  reg                 io_B_Valid_29_delay_1;
  reg                 io_A_Valid_1_delay_1_29;
  reg                 io_A_Valid_1_delay_2_28;
  reg                 io_A_Valid_1_delay_3_27;
  reg                 io_A_Valid_1_delay_4_26;
  reg                 io_A_Valid_1_delay_5_25;
  reg                 io_A_Valid_1_delay_6_24;
  reg                 io_A_Valid_1_delay_7_23;
  reg                 io_A_Valid_1_delay_8_22;
  reg                 io_A_Valid_1_delay_9_21;
  reg                 io_A_Valid_1_delay_10_20;
  reg                 io_A_Valid_1_delay_11_19;
  reg                 io_A_Valid_1_delay_12_18;
  reg                 io_A_Valid_1_delay_13_17;
  reg                 io_A_Valid_1_delay_14_16;
  reg                 io_A_Valid_1_delay_15_15;
  reg                 io_A_Valid_1_delay_16_14;
  reg                 io_A_Valid_1_delay_17_13;
  reg                 io_A_Valid_1_delay_18_12;
  reg                 io_A_Valid_1_delay_19_11;
  reg                 io_A_Valid_1_delay_20_10;
  reg                 io_A_Valid_1_delay_21_9;
  reg                 io_A_Valid_1_delay_22_8;
  reg                 io_A_Valid_1_delay_23_7;
  reg                 io_A_Valid_1_delay_24_6;
  reg                 io_A_Valid_1_delay_25_5;
  reg                 io_A_Valid_1_delay_26_4;
  reg                 io_A_Valid_1_delay_27_3;
  reg                 io_A_Valid_1_delay_28_2;
  reg                 io_A_Valid_1_delay_29_1;
  reg                 io_A_Valid_1_delay_30;
  reg                 io_B_Valid_30_delay_1;
  reg                 io_A_Valid_1_delay_1_30;
  reg                 io_A_Valid_1_delay_2_29;
  reg                 io_A_Valid_1_delay_3_28;
  reg                 io_A_Valid_1_delay_4_27;
  reg                 io_A_Valid_1_delay_5_26;
  reg                 io_A_Valid_1_delay_6_25;
  reg                 io_A_Valid_1_delay_7_24;
  reg                 io_A_Valid_1_delay_8_23;
  reg                 io_A_Valid_1_delay_9_22;
  reg                 io_A_Valid_1_delay_10_21;
  reg                 io_A_Valid_1_delay_11_20;
  reg                 io_A_Valid_1_delay_12_19;
  reg                 io_A_Valid_1_delay_13_18;
  reg                 io_A_Valid_1_delay_14_17;
  reg                 io_A_Valid_1_delay_15_16;
  reg                 io_A_Valid_1_delay_16_15;
  reg                 io_A_Valid_1_delay_17_14;
  reg                 io_A_Valid_1_delay_18_13;
  reg                 io_A_Valid_1_delay_19_12;
  reg                 io_A_Valid_1_delay_20_11;
  reg                 io_A_Valid_1_delay_21_10;
  reg                 io_A_Valid_1_delay_22_9;
  reg                 io_A_Valid_1_delay_23_8;
  reg                 io_A_Valid_1_delay_24_7;
  reg                 io_A_Valid_1_delay_25_6;
  reg                 io_A_Valid_1_delay_26_5;
  reg                 io_A_Valid_1_delay_27_4;
  reg                 io_A_Valid_1_delay_28_3;
  reg                 io_A_Valid_1_delay_29_2;
  reg                 io_A_Valid_1_delay_30_1;
  reg                 io_A_Valid_1_delay_31;
  reg                 io_B_Valid_31_delay_1;
  reg                 io_A_Valid_1_delay_1_31;
  reg                 io_A_Valid_1_delay_2_30;
  reg                 io_A_Valid_1_delay_3_29;
  reg                 io_A_Valid_1_delay_4_28;
  reg                 io_A_Valid_1_delay_5_27;
  reg                 io_A_Valid_1_delay_6_26;
  reg                 io_A_Valid_1_delay_7_25;
  reg                 io_A_Valid_1_delay_8_24;
  reg                 io_A_Valid_1_delay_9_23;
  reg                 io_A_Valid_1_delay_10_22;
  reg                 io_A_Valid_1_delay_11_21;
  reg                 io_A_Valid_1_delay_12_20;
  reg                 io_A_Valid_1_delay_13_19;
  reg                 io_A_Valid_1_delay_14_18;
  reg                 io_A_Valid_1_delay_15_17;
  reg                 io_A_Valid_1_delay_16_16;
  reg                 io_A_Valid_1_delay_17_15;
  reg                 io_A_Valid_1_delay_18_14;
  reg                 io_A_Valid_1_delay_19_13;
  reg                 io_A_Valid_1_delay_20_12;
  reg                 io_A_Valid_1_delay_21_11;
  reg                 io_A_Valid_1_delay_22_10;
  reg                 io_A_Valid_1_delay_23_9;
  reg                 io_A_Valid_1_delay_24_8;
  reg                 io_A_Valid_1_delay_25_7;
  reg                 io_A_Valid_1_delay_26_6;
  reg                 io_A_Valid_1_delay_27_5;
  reg                 io_A_Valid_1_delay_28_4;
  reg                 io_A_Valid_1_delay_29_3;
  reg                 io_A_Valid_1_delay_30_2;
  reg                 io_A_Valid_1_delay_31_1;
  reg                 io_A_Valid_1_delay_32;
  reg                 io_B_Valid_32_delay_1;
  reg                 io_A_Valid_1_delay_1_32;
  reg                 io_A_Valid_1_delay_2_31;
  reg                 io_A_Valid_1_delay_3_30;
  reg                 io_A_Valid_1_delay_4_29;
  reg                 io_A_Valid_1_delay_5_28;
  reg                 io_A_Valid_1_delay_6_27;
  reg                 io_A_Valid_1_delay_7_26;
  reg                 io_A_Valid_1_delay_8_25;
  reg                 io_A_Valid_1_delay_9_24;
  reg                 io_A_Valid_1_delay_10_23;
  reg                 io_A_Valid_1_delay_11_22;
  reg                 io_A_Valid_1_delay_12_21;
  reg                 io_A_Valid_1_delay_13_20;
  reg                 io_A_Valid_1_delay_14_19;
  reg                 io_A_Valid_1_delay_15_18;
  reg                 io_A_Valid_1_delay_16_17;
  reg                 io_A_Valid_1_delay_17_16;
  reg                 io_A_Valid_1_delay_18_15;
  reg                 io_A_Valid_1_delay_19_14;
  reg                 io_A_Valid_1_delay_20_13;
  reg                 io_A_Valid_1_delay_21_12;
  reg                 io_A_Valid_1_delay_22_11;
  reg                 io_A_Valid_1_delay_23_10;
  reg                 io_A_Valid_1_delay_24_9;
  reg                 io_A_Valid_1_delay_25_8;
  reg                 io_A_Valid_1_delay_26_7;
  reg                 io_A_Valid_1_delay_27_6;
  reg                 io_A_Valid_1_delay_28_5;
  reg                 io_A_Valid_1_delay_29_4;
  reg                 io_A_Valid_1_delay_30_3;
  reg                 io_A_Valid_1_delay_31_2;
  reg                 io_A_Valid_1_delay_32_1;
  reg                 io_A_Valid_1_delay_33;
  reg                 io_B_Valid_33_delay_1;
  reg                 io_A_Valid_1_delay_1_33;
  reg                 io_A_Valid_1_delay_2_32;
  reg                 io_A_Valid_1_delay_3_31;
  reg                 io_A_Valid_1_delay_4_30;
  reg                 io_A_Valid_1_delay_5_29;
  reg                 io_A_Valid_1_delay_6_28;
  reg                 io_A_Valid_1_delay_7_27;
  reg                 io_A_Valid_1_delay_8_26;
  reg                 io_A_Valid_1_delay_9_25;
  reg                 io_A_Valid_1_delay_10_24;
  reg                 io_A_Valid_1_delay_11_23;
  reg                 io_A_Valid_1_delay_12_22;
  reg                 io_A_Valid_1_delay_13_21;
  reg                 io_A_Valid_1_delay_14_20;
  reg                 io_A_Valid_1_delay_15_19;
  reg                 io_A_Valid_1_delay_16_18;
  reg                 io_A_Valid_1_delay_17_17;
  reg                 io_A_Valid_1_delay_18_16;
  reg                 io_A_Valid_1_delay_19_15;
  reg                 io_A_Valid_1_delay_20_14;
  reg                 io_A_Valid_1_delay_21_13;
  reg                 io_A_Valid_1_delay_22_12;
  reg                 io_A_Valid_1_delay_23_11;
  reg                 io_A_Valid_1_delay_24_10;
  reg                 io_A_Valid_1_delay_25_9;
  reg                 io_A_Valid_1_delay_26_8;
  reg                 io_A_Valid_1_delay_27_7;
  reg                 io_A_Valid_1_delay_28_6;
  reg                 io_A_Valid_1_delay_29_5;
  reg                 io_A_Valid_1_delay_30_4;
  reg                 io_A_Valid_1_delay_31_3;
  reg                 io_A_Valid_1_delay_32_2;
  reg                 io_A_Valid_1_delay_33_1;
  reg                 io_A_Valid_1_delay_34;
  reg                 io_B_Valid_34_delay_1;
  reg                 io_A_Valid_1_delay_1_34;
  reg                 io_A_Valid_1_delay_2_33;
  reg                 io_A_Valid_1_delay_3_32;
  reg                 io_A_Valid_1_delay_4_31;
  reg                 io_A_Valid_1_delay_5_30;
  reg                 io_A_Valid_1_delay_6_29;
  reg                 io_A_Valid_1_delay_7_28;
  reg                 io_A_Valid_1_delay_8_27;
  reg                 io_A_Valid_1_delay_9_26;
  reg                 io_A_Valid_1_delay_10_25;
  reg                 io_A_Valid_1_delay_11_24;
  reg                 io_A_Valid_1_delay_12_23;
  reg                 io_A_Valid_1_delay_13_22;
  reg                 io_A_Valid_1_delay_14_21;
  reg                 io_A_Valid_1_delay_15_20;
  reg                 io_A_Valid_1_delay_16_19;
  reg                 io_A_Valid_1_delay_17_18;
  reg                 io_A_Valid_1_delay_18_17;
  reg                 io_A_Valid_1_delay_19_16;
  reg                 io_A_Valid_1_delay_20_15;
  reg                 io_A_Valid_1_delay_21_14;
  reg                 io_A_Valid_1_delay_22_13;
  reg                 io_A_Valid_1_delay_23_12;
  reg                 io_A_Valid_1_delay_24_11;
  reg                 io_A_Valid_1_delay_25_10;
  reg                 io_A_Valid_1_delay_26_9;
  reg                 io_A_Valid_1_delay_27_8;
  reg                 io_A_Valid_1_delay_28_7;
  reg                 io_A_Valid_1_delay_29_6;
  reg                 io_A_Valid_1_delay_30_5;
  reg                 io_A_Valid_1_delay_31_4;
  reg                 io_A_Valid_1_delay_32_3;
  reg                 io_A_Valid_1_delay_33_2;
  reg                 io_A_Valid_1_delay_34_1;
  reg                 io_A_Valid_1_delay_35;
  reg                 io_B_Valid_35_delay_1;
  reg                 io_A_Valid_1_delay_1_35;
  reg                 io_A_Valid_1_delay_2_34;
  reg                 io_A_Valid_1_delay_3_33;
  reg                 io_A_Valid_1_delay_4_32;
  reg                 io_A_Valid_1_delay_5_31;
  reg                 io_A_Valid_1_delay_6_30;
  reg                 io_A_Valid_1_delay_7_29;
  reg                 io_A_Valid_1_delay_8_28;
  reg                 io_A_Valid_1_delay_9_27;
  reg                 io_A_Valid_1_delay_10_26;
  reg                 io_A_Valid_1_delay_11_25;
  reg                 io_A_Valid_1_delay_12_24;
  reg                 io_A_Valid_1_delay_13_23;
  reg                 io_A_Valid_1_delay_14_22;
  reg                 io_A_Valid_1_delay_15_21;
  reg                 io_A_Valid_1_delay_16_20;
  reg                 io_A_Valid_1_delay_17_19;
  reg                 io_A_Valid_1_delay_18_18;
  reg                 io_A_Valid_1_delay_19_17;
  reg                 io_A_Valid_1_delay_20_16;
  reg                 io_A_Valid_1_delay_21_15;
  reg                 io_A_Valid_1_delay_22_14;
  reg                 io_A_Valid_1_delay_23_13;
  reg                 io_A_Valid_1_delay_24_12;
  reg                 io_A_Valid_1_delay_25_11;
  reg                 io_A_Valid_1_delay_26_10;
  reg                 io_A_Valid_1_delay_27_9;
  reg                 io_A_Valid_1_delay_28_8;
  reg                 io_A_Valid_1_delay_29_7;
  reg                 io_A_Valid_1_delay_30_6;
  reg                 io_A_Valid_1_delay_31_5;
  reg                 io_A_Valid_1_delay_32_4;
  reg                 io_A_Valid_1_delay_33_3;
  reg                 io_A_Valid_1_delay_34_2;
  reg                 io_A_Valid_1_delay_35_1;
  reg                 io_A_Valid_1_delay_36;
  reg                 io_B_Valid_36_delay_1;
  reg                 io_A_Valid_1_delay_1_36;
  reg                 io_A_Valid_1_delay_2_35;
  reg                 io_A_Valid_1_delay_3_34;
  reg                 io_A_Valid_1_delay_4_33;
  reg                 io_A_Valid_1_delay_5_32;
  reg                 io_A_Valid_1_delay_6_31;
  reg                 io_A_Valid_1_delay_7_30;
  reg                 io_A_Valid_1_delay_8_29;
  reg                 io_A_Valid_1_delay_9_28;
  reg                 io_A_Valid_1_delay_10_27;
  reg                 io_A_Valid_1_delay_11_26;
  reg                 io_A_Valid_1_delay_12_25;
  reg                 io_A_Valid_1_delay_13_24;
  reg                 io_A_Valid_1_delay_14_23;
  reg                 io_A_Valid_1_delay_15_22;
  reg                 io_A_Valid_1_delay_16_21;
  reg                 io_A_Valid_1_delay_17_20;
  reg                 io_A_Valid_1_delay_18_19;
  reg                 io_A_Valid_1_delay_19_18;
  reg                 io_A_Valid_1_delay_20_17;
  reg                 io_A_Valid_1_delay_21_16;
  reg                 io_A_Valid_1_delay_22_15;
  reg                 io_A_Valid_1_delay_23_14;
  reg                 io_A_Valid_1_delay_24_13;
  reg                 io_A_Valid_1_delay_25_12;
  reg                 io_A_Valid_1_delay_26_11;
  reg                 io_A_Valid_1_delay_27_10;
  reg                 io_A_Valid_1_delay_28_9;
  reg                 io_A_Valid_1_delay_29_8;
  reg                 io_A_Valid_1_delay_30_7;
  reg                 io_A_Valid_1_delay_31_6;
  reg                 io_A_Valid_1_delay_32_5;
  reg                 io_A_Valid_1_delay_33_4;
  reg                 io_A_Valid_1_delay_34_3;
  reg                 io_A_Valid_1_delay_35_2;
  reg                 io_A_Valid_1_delay_36_1;
  reg                 io_A_Valid_1_delay_37;
  reg                 io_B_Valid_37_delay_1;
  reg                 io_A_Valid_1_delay_1_37;
  reg                 io_A_Valid_1_delay_2_36;
  reg                 io_A_Valid_1_delay_3_35;
  reg                 io_A_Valid_1_delay_4_34;
  reg                 io_A_Valid_1_delay_5_33;
  reg                 io_A_Valid_1_delay_6_32;
  reg                 io_A_Valid_1_delay_7_31;
  reg                 io_A_Valid_1_delay_8_30;
  reg                 io_A_Valid_1_delay_9_29;
  reg                 io_A_Valid_1_delay_10_28;
  reg                 io_A_Valid_1_delay_11_27;
  reg                 io_A_Valid_1_delay_12_26;
  reg                 io_A_Valid_1_delay_13_25;
  reg                 io_A_Valid_1_delay_14_24;
  reg                 io_A_Valid_1_delay_15_23;
  reg                 io_A_Valid_1_delay_16_22;
  reg                 io_A_Valid_1_delay_17_21;
  reg                 io_A_Valid_1_delay_18_20;
  reg                 io_A_Valid_1_delay_19_19;
  reg                 io_A_Valid_1_delay_20_18;
  reg                 io_A_Valid_1_delay_21_17;
  reg                 io_A_Valid_1_delay_22_16;
  reg                 io_A_Valid_1_delay_23_15;
  reg                 io_A_Valid_1_delay_24_14;
  reg                 io_A_Valid_1_delay_25_13;
  reg                 io_A_Valid_1_delay_26_12;
  reg                 io_A_Valid_1_delay_27_11;
  reg                 io_A_Valid_1_delay_28_10;
  reg                 io_A_Valid_1_delay_29_9;
  reg                 io_A_Valid_1_delay_30_8;
  reg                 io_A_Valid_1_delay_31_7;
  reg                 io_A_Valid_1_delay_32_6;
  reg                 io_A_Valid_1_delay_33_5;
  reg                 io_A_Valid_1_delay_34_4;
  reg                 io_A_Valid_1_delay_35_3;
  reg                 io_A_Valid_1_delay_36_2;
  reg                 io_A_Valid_1_delay_37_1;
  reg                 io_A_Valid_1_delay_38;
  reg                 io_B_Valid_38_delay_1;
  reg                 io_A_Valid_1_delay_1_38;
  reg                 io_A_Valid_1_delay_2_37;
  reg                 io_A_Valid_1_delay_3_36;
  reg                 io_A_Valid_1_delay_4_35;
  reg                 io_A_Valid_1_delay_5_34;
  reg                 io_A_Valid_1_delay_6_33;
  reg                 io_A_Valid_1_delay_7_32;
  reg                 io_A_Valid_1_delay_8_31;
  reg                 io_A_Valid_1_delay_9_30;
  reg                 io_A_Valid_1_delay_10_29;
  reg                 io_A_Valid_1_delay_11_28;
  reg                 io_A_Valid_1_delay_12_27;
  reg                 io_A_Valid_1_delay_13_26;
  reg                 io_A_Valid_1_delay_14_25;
  reg                 io_A_Valid_1_delay_15_24;
  reg                 io_A_Valid_1_delay_16_23;
  reg                 io_A_Valid_1_delay_17_22;
  reg                 io_A_Valid_1_delay_18_21;
  reg                 io_A_Valid_1_delay_19_20;
  reg                 io_A_Valid_1_delay_20_19;
  reg                 io_A_Valid_1_delay_21_18;
  reg                 io_A_Valid_1_delay_22_17;
  reg                 io_A_Valid_1_delay_23_16;
  reg                 io_A_Valid_1_delay_24_15;
  reg                 io_A_Valid_1_delay_25_14;
  reg                 io_A_Valid_1_delay_26_13;
  reg                 io_A_Valid_1_delay_27_12;
  reg                 io_A_Valid_1_delay_28_11;
  reg                 io_A_Valid_1_delay_29_10;
  reg                 io_A_Valid_1_delay_30_9;
  reg                 io_A_Valid_1_delay_31_8;
  reg                 io_A_Valid_1_delay_32_7;
  reg                 io_A_Valid_1_delay_33_6;
  reg                 io_A_Valid_1_delay_34_5;
  reg                 io_A_Valid_1_delay_35_4;
  reg                 io_A_Valid_1_delay_36_3;
  reg                 io_A_Valid_1_delay_37_2;
  reg                 io_A_Valid_1_delay_38_1;
  reg                 io_A_Valid_1_delay_39;
  reg                 io_B_Valid_39_delay_1;
  reg                 io_A_Valid_1_delay_1_39;
  reg                 io_A_Valid_1_delay_2_38;
  reg                 io_A_Valid_1_delay_3_37;
  reg                 io_A_Valid_1_delay_4_36;
  reg                 io_A_Valid_1_delay_5_35;
  reg                 io_A_Valid_1_delay_6_34;
  reg                 io_A_Valid_1_delay_7_33;
  reg                 io_A_Valid_1_delay_8_32;
  reg                 io_A_Valid_1_delay_9_31;
  reg                 io_A_Valid_1_delay_10_30;
  reg                 io_A_Valid_1_delay_11_29;
  reg                 io_A_Valid_1_delay_12_28;
  reg                 io_A_Valid_1_delay_13_27;
  reg                 io_A_Valid_1_delay_14_26;
  reg                 io_A_Valid_1_delay_15_25;
  reg                 io_A_Valid_1_delay_16_24;
  reg                 io_A_Valid_1_delay_17_23;
  reg                 io_A_Valid_1_delay_18_22;
  reg                 io_A_Valid_1_delay_19_21;
  reg                 io_A_Valid_1_delay_20_20;
  reg                 io_A_Valid_1_delay_21_19;
  reg                 io_A_Valid_1_delay_22_18;
  reg                 io_A_Valid_1_delay_23_17;
  reg                 io_A_Valid_1_delay_24_16;
  reg                 io_A_Valid_1_delay_25_15;
  reg                 io_A_Valid_1_delay_26_14;
  reg                 io_A_Valid_1_delay_27_13;
  reg                 io_A_Valid_1_delay_28_12;
  reg                 io_A_Valid_1_delay_29_11;
  reg                 io_A_Valid_1_delay_30_10;
  reg                 io_A_Valid_1_delay_31_9;
  reg                 io_A_Valid_1_delay_32_8;
  reg                 io_A_Valid_1_delay_33_7;
  reg                 io_A_Valid_1_delay_34_6;
  reg                 io_A_Valid_1_delay_35_5;
  reg                 io_A_Valid_1_delay_36_4;
  reg                 io_A_Valid_1_delay_37_3;
  reg                 io_A_Valid_1_delay_38_2;
  reg                 io_A_Valid_1_delay_39_1;
  reg                 io_A_Valid_1_delay_40;
  reg                 io_B_Valid_40_delay_1;
  reg                 io_A_Valid_1_delay_1_40;
  reg                 io_A_Valid_1_delay_2_39;
  reg                 io_A_Valid_1_delay_3_38;
  reg                 io_A_Valid_1_delay_4_37;
  reg                 io_A_Valid_1_delay_5_36;
  reg                 io_A_Valid_1_delay_6_35;
  reg                 io_A_Valid_1_delay_7_34;
  reg                 io_A_Valid_1_delay_8_33;
  reg                 io_A_Valid_1_delay_9_32;
  reg                 io_A_Valid_1_delay_10_31;
  reg                 io_A_Valid_1_delay_11_30;
  reg                 io_A_Valid_1_delay_12_29;
  reg                 io_A_Valid_1_delay_13_28;
  reg                 io_A_Valid_1_delay_14_27;
  reg                 io_A_Valid_1_delay_15_26;
  reg                 io_A_Valid_1_delay_16_25;
  reg                 io_A_Valid_1_delay_17_24;
  reg                 io_A_Valid_1_delay_18_23;
  reg                 io_A_Valid_1_delay_19_22;
  reg                 io_A_Valid_1_delay_20_21;
  reg                 io_A_Valid_1_delay_21_20;
  reg                 io_A_Valid_1_delay_22_19;
  reg                 io_A_Valid_1_delay_23_18;
  reg                 io_A_Valid_1_delay_24_17;
  reg                 io_A_Valid_1_delay_25_16;
  reg                 io_A_Valid_1_delay_26_15;
  reg                 io_A_Valid_1_delay_27_14;
  reg                 io_A_Valid_1_delay_28_13;
  reg                 io_A_Valid_1_delay_29_12;
  reg                 io_A_Valid_1_delay_30_11;
  reg                 io_A_Valid_1_delay_31_10;
  reg                 io_A_Valid_1_delay_32_9;
  reg                 io_A_Valid_1_delay_33_8;
  reg                 io_A_Valid_1_delay_34_7;
  reg                 io_A_Valid_1_delay_35_6;
  reg                 io_A_Valid_1_delay_36_5;
  reg                 io_A_Valid_1_delay_37_4;
  reg                 io_A_Valid_1_delay_38_3;
  reg                 io_A_Valid_1_delay_39_2;
  reg                 io_A_Valid_1_delay_40_1;
  reg                 io_A_Valid_1_delay_41;
  reg                 io_B_Valid_41_delay_1;
  reg                 io_A_Valid_1_delay_1_41;
  reg                 io_A_Valid_1_delay_2_40;
  reg                 io_A_Valid_1_delay_3_39;
  reg                 io_A_Valid_1_delay_4_38;
  reg                 io_A_Valid_1_delay_5_37;
  reg                 io_A_Valid_1_delay_6_36;
  reg                 io_A_Valid_1_delay_7_35;
  reg                 io_A_Valid_1_delay_8_34;
  reg                 io_A_Valid_1_delay_9_33;
  reg                 io_A_Valid_1_delay_10_32;
  reg                 io_A_Valid_1_delay_11_31;
  reg                 io_A_Valid_1_delay_12_30;
  reg                 io_A_Valid_1_delay_13_29;
  reg                 io_A_Valid_1_delay_14_28;
  reg                 io_A_Valid_1_delay_15_27;
  reg                 io_A_Valid_1_delay_16_26;
  reg                 io_A_Valid_1_delay_17_25;
  reg                 io_A_Valid_1_delay_18_24;
  reg                 io_A_Valid_1_delay_19_23;
  reg                 io_A_Valid_1_delay_20_22;
  reg                 io_A_Valid_1_delay_21_21;
  reg                 io_A_Valid_1_delay_22_20;
  reg                 io_A_Valid_1_delay_23_19;
  reg                 io_A_Valid_1_delay_24_18;
  reg                 io_A_Valid_1_delay_25_17;
  reg                 io_A_Valid_1_delay_26_16;
  reg                 io_A_Valid_1_delay_27_15;
  reg                 io_A_Valid_1_delay_28_14;
  reg                 io_A_Valid_1_delay_29_13;
  reg                 io_A_Valid_1_delay_30_12;
  reg                 io_A_Valid_1_delay_31_11;
  reg                 io_A_Valid_1_delay_32_10;
  reg                 io_A_Valid_1_delay_33_9;
  reg                 io_A_Valid_1_delay_34_8;
  reg                 io_A_Valid_1_delay_35_7;
  reg                 io_A_Valid_1_delay_36_6;
  reg                 io_A_Valid_1_delay_37_5;
  reg                 io_A_Valid_1_delay_38_4;
  reg                 io_A_Valid_1_delay_39_3;
  reg                 io_A_Valid_1_delay_40_2;
  reg                 io_A_Valid_1_delay_41_1;
  reg                 io_A_Valid_1_delay_42;
  reg                 io_B_Valid_42_delay_1;
  reg                 io_A_Valid_1_delay_1_42;
  reg                 io_A_Valid_1_delay_2_41;
  reg                 io_A_Valid_1_delay_3_40;
  reg                 io_A_Valid_1_delay_4_39;
  reg                 io_A_Valid_1_delay_5_38;
  reg                 io_A_Valid_1_delay_6_37;
  reg                 io_A_Valid_1_delay_7_36;
  reg                 io_A_Valid_1_delay_8_35;
  reg                 io_A_Valid_1_delay_9_34;
  reg                 io_A_Valid_1_delay_10_33;
  reg                 io_A_Valid_1_delay_11_32;
  reg                 io_A_Valid_1_delay_12_31;
  reg                 io_A_Valid_1_delay_13_30;
  reg                 io_A_Valid_1_delay_14_29;
  reg                 io_A_Valid_1_delay_15_28;
  reg                 io_A_Valid_1_delay_16_27;
  reg                 io_A_Valid_1_delay_17_26;
  reg                 io_A_Valid_1_delay_18_25;
  reg                 io_A_Valid_1_delay_19_24;
  reg                 io_A_Valid_1_delay_20_23;
  reg                 io_A_Valid_1_delay_21_22;
  reg                 io_A_Valid_1_delay_22_21;
  reg                 io_A_Valid_1_delay_23_20;
  reg                 io_A_Valid_1_delay_24_19;
  reg                 io_A_Valid_1_delay_25_18;
  reg                 io_A_Valid_1_delay_26_17;
  reg                 io_A_Valid_1_delay_27_16;
  reg                 io_A_Valid_1_delay_28_15;
  reg                 io_A_Valid_1_delay_29_14;
  reg                 io_A_Valid_1_delay_30_13;
  reg                 io_A_Valid_1_delay_31_12;
  reg                 io_A_Valid_1_delay_32_11;
  reg                 io_A_Valid_1_delay_33_10;
  reg                 io_A_Valid_1_delay_34_9;
  reg                 io_A_Valid_1_delay_35_8;
  reg                 io_A_Valid_1_delay_36_7;
  reg                 io_A_Valid_1_delay_37_6;
  reg                 io_A_Valid_1_delay_38_5;
  reg                 io_A_Valid_1_delay_39_4;
  reg                 io_A_Valid_1_delay_40_3;
  reg                 io_A_Valid_1_delay_41_2;
  reg                 io_A_Valid_1_delay_42_1;
  reg                 io_A_Valid_1_delay_43;
  reg                 io_B_Valid_43_delay_1;
  reg                 io_A_Valid_1_delay_1_43;
  reg                 io_A_Valid_1_delay_2_42;
  reg                 io_A_Valid_1_delay_3_41;
  reg                 io_A_Valid_1_delay_4_40;
  reg                 io_A_Valid_1_delay_5_39;
  reg                 io_A_Valid_1_delay_6_38;
  reg                 io_A_Valid_1_delay_7_37;
  reg                 io_A_Valid_1_delay_8_36;
  reg                 io_A_Valid_1_delay_9_35;
  reg                 io_A_Valid_1_delay_10_34;
  reg                 io_A_Valid_1_delay_11_33;
  reg                 io_A_Valid_1_delay_12_32;
  reg                 io_A_Valid_1_delay_13_31;
  reg                 io_A_Valid_1_delay_14_30;
  reg                 io_A_Valid_1_delay_15_29;
  reg                 io_A_Valid_1_delay_16_28;
  reg                 io_A_Valid_1_delay_17_27;
  reg                 io_A_Valid_1_delay_18_26;
  reg                 io_A_Valid_1_delay_19_25;
  reg                 io_A_Valid_1_delay_20_24;
  reg                 io_A_Valid_1_delay_21_23;
  reg                 io_A_Valid_1_delay_22_22;
  reg                 io_A_Valid_1_delay_23_21;
  reg                 io_A_Valid_1_delay_24_20;
  reg                 io_A_Valid_1_delay_25_19;
  reg                 io_A_Valid_1_delay_26_18;
  reg                 io_A_Valid_1_delay_27_17;
  reg                 io_A_Valid_1_delay_28_16;
  reg                 io_A_Valid_1_delay_29_15;
  reg                 io_A_Valid_1_delay_30_14;
  reg                 io_A_Valid_1_delay_31_13;
  reg                 io_A_Valid_1_delay_32_12;
  reg                 io_A_Valid_1_delay_33_11;
  reg                 io_A_Valid_1_delay_34_10;
  reg                 io_A_Valid_1_delay_35_9;
  reg                 io_A_Valid_1_delay_36_8;
  reg                 io_A_Valid_1_delay_37_7;
  reg                 io_A_Valid_1_delay_38_6;
  reg                 io_A_Valid_1_delay_39_5;
  reg                 io_A_Valid_1_delay_40_4;
  reg                 io_A_Valid_1_delay_41_3;
  reg                 io_A_Valid_1_delay_42_2;
  reg                 io_A_Valid_1_delay_43_1;
  reg                 io_A_Valid_1_delay_44;
  reg                 io_B_Valid_44_delay_1;
  reg                 io_A_Valid_1_delay_1_44;
  reg                 io_A_Valid_1_delay_2_43;
  reg                 io_A_Valid_1_delay_3_42;
  reg                 io_A_Valid_1_delay_4_41;
  reg                 io_A_Valid_1_delay_5_40;
  reg                 io_A_Valid_1_delay_6_39;
  reg                 io_A_Valid_1_delay_7_38;
  reg                 io_A_Valid_1_delay_8_37;
  reg                 io_A_Valid_1_delay_9_36;
  reg                 io_A_Valid_1_delay_10_35;
  reg                 io_A_Valid_1_delay_11_34;
  reg                 io_A_Valid_1_delay_12_33;
  reg                 io_A_Valid_1_delay_13_32;
  reg                 io_A_Valid_1_delay_14_31;
  reg                 io_A_Valid_1_delay_15_30;
  reg                 io_A_Valid_1_delay_16_29;
  reg                 io_A_Valid_1_delay_17_28;
  reg                 io_A_Valid_1_delay_18_27;
  reg                 io_A_Valid_1_delay_19_26;
  reg                 io_A_Valid_1_delay_20_25;
  reg                 io_A_Valid_1_delay_21_24;
  reg                 io_A_Valid_1_delay_22_23;
  reg                 io_A_Valid_1_delay_23_22;
  reg                 io_A_Valid_1_delay_24_21;
  reg                 io_A_Valid_1_delay_25_20;
  reg                 io_A_Valid_1_delay_26_19;
  reg                 io_A_Valid_1_delay_27_18;
  reg                 io_A_Valid_1_delay_28_17;
  reg                 io_A_Valid_1_delay_29_16;
  reg                 io_A_Valid_1_delay_30_15;
  reg                 io_A_Valid_1_delay_31_14;
  reg                 io_A_Valid_1_delay_32_13;
  reg                 io_A_Valid_1_delay_33_12;
  reg                 io_A_Valid_1_delay_34_11;
  reg                 io_A_Valid_1_delay_35_10;
  reg                 io_A_Valid_1_delay_36_9;
  reg                 io_A_Valid_1_delay_37_8;
  reg                 io_A_Valid_1_delay_38_7;
  reg                 io_A_Valid_1_delay_39_6;
  reg                 io_A_Valid_1_delay_40_5;
  reg                 io_A_Valid_1_delay_41_4;
  reg                 io_A_Valid_1_delay_42_3;
  reg                 io_A_Valid_1_delay_43_2;
  reg                 io_A_Valid_1_delay_44_1;
  reg                 io_A_Valid_1_delay_45;
  reg                 io_B_Valid_45_delay_1;
  reg                 io_A_Valid_1_delay_1_45;
  reg                 io_A_Valid_1_delay_2_44;
  reg                 io_A_Valid_1_delay_3_43;
  reg                 io_A_Valid_1_delay_4_42;
  reg                 io_A_Valid_1_delay_5_41;
  reg                 io_A_Valid_1_delay_6_40;
  reg                 io_A_Valid_1_delay_7_39;
  reg                 io_A_Valid_1_delay_8_38;
  reg                 io_A_Valid_1_delay_9_37;
  reg                 io_A_Valid_1_delay_10_36;
  reg                 io_A_Valid_1_delay_11_35;
  reg                 io_A_Valid_1_delay_12_34;
  reg                 io_A_Valid_1_delay_13_33;
  reg                 io_A_Valid_1_delay_14_32;
  reg                 io_A_Valid_1_delay_15_31;
  reg                 io_A_Valid_1_delay_16_30;
  reg                 io_A_Valid_1_delay_17_29;
  reg                 io_A_Valid_1_delay_18_28;
  reg                 io_A_Valid_1_delay_19_27;
  reg                 io_A_Valid_1_delay_20_26;
  reg                 io_A_Valid_1_delay_21_25;
  reg                 io_A_Valid_1_delay_22_24;
  reg                 io_A_Valid_1_delay_23_23;
  reg                 io_A_Valid_1_delay_24_22;
  reg                 io_A_Valid_1_delay_25_21;
  reg                 io_A_Valid_1_delay_26_20;
  reg                 io_A_Valid_1_delay_27_19;
  reg                 io_A_Valid_1_delay_28_18;
  reg                 io_A_Valid_1_delay_29_17;
  reg                 io_A_Valid_1_delay_30_16;
  reg                 io_A_Valid_1_delay_31_15;
  reg                 io_A_Valid_1_delay_32_14;
  reg                 io_A_Valid_1_delay_33_13;
  reg                 io_A_Valid_1_delay_34_12;
  reg                 io_A_Valid_1_delay_35_11;
  reg                 io_A_Valid_1_delay_36_10;
  reg                 io_A_Valid_1_delay_37_9;
  reg                 io_A_Valid_1_delay_38_8;
  reg                 io_A_Valid_1_delay_39_7;
  reg                 io_A_Valid_1_delay_40_6;
  reg                 io_A_Valid_1_delay_41_5;
  reg                 io_A_Valid_1_delay_42_4;
  reg                 io_A_Valid_1_delay_43_3;
  reg                 io_A_Valid_1_delay_44_2;
  reg                 io_A_Valid_1_delay_45_1;
  reg                 io_A_Valid_1_delay_46;
  reg                 io_B_Valid_46_delay_1;
  reg                 io_A_Valid_1_delay_1_46;
  reg                 io_A_Valid_1_delay_2_45;
  reg                 io_A_Valid_1_delay_3_44;
  reg                 io_A_Valid_1_delay_4_43;
  reg                 io_A_Valid_1_delay_5_42;
  reg                 io_A_Valid_1_delay_6_41;
  reg                 io_A_Valid_1_delay_7_40;
  reg                 io_A_Valid_1_delay_8_39;
  reg                 io_A_Valid_1_delay_9_38;
  reg                 io_A_Valid_1_delay_10_37;
  reg                 io_A_Valid_1_delay_11_36;
  reg                 io_A_Valid_1_delay_12_35;
  reg                 io_A_Valid_1_delay_13_34;
  reg                 io_A_Valid_1_delay_14_33;
  reg                 io_A_Valid_1_delay_15_32;
  reg                 io_A_Valid_1_delay_16_31;
  reg                 io_A_Valid_1_delay_17_30;
  reg                 io_A_Valid_1_delay_18_29;
  reg                 io_A_Valid_1_delay_19_28;
  reg                 io_A_Valid_1_delay_20_27;
  reg                 io_A_Valid_1_delay_21_26;
  reg                 io_A_Valid_1_delay_22_25;
  reg                 io_A_Valid_1_delay_23_24;
  reg                 io_A_Valid_1_delay_24_23;
  reg                 io_A_Valid_1_delay_25_22;
  reg                 io_A_Valid_1_delay_26_21;
  reg                 io_A_Valid_1_delay_27_20;
  reg                 io_A_Valid_1_delay_28_19;
  reg                 io_A_Valid_1_delay_29_18;
  reg                 io_A_Valid_1_delay_30_17;
  reg                 io_A_Valid_1_delay_31_16;
  reg                 io_A_Valid_1_delay_32_15;
  reg                 io_A_Valid_1_delay_33_14;
  reg                 io_A_Valid_1_delay_34_13;
  reg                 io_A_Valid_1_delay_35_12;
  reg                 io_A_Valid_1_delay_36_11;
  reg                 io_A_Valid_1_delay_37_10;
  reg                 io_A_Valid_1_delay_38_9;
  reg                 io_A_Valid_1_delay_39_8;
  reg                 io_A_Valid_1_delay_40_7;
  reg                 io_A_Valid_1_delay_41_6;
  reg                 io_A_Valid_1_delay_42_5;
  reg                 io_A_Valid_1_delay_43_4;
  reg                 io_A_Valid_1_delay_44_3;
  reg                 io_A_Valid_1_delay_45_2;
  reg                 io_A_Valid_1_delay_46_1;
  reg                 io_A_Valid_1_delay_47;
  reg                 io_B_Valid_47_delay_1;
  reg                 io_A_Valid_1_delay_1_47;
  reg                 io_A_Valid_1_delay_2_46;
  reg                 io_A_Valid_1_delay_3_45;
  reg                 io_A_Valid_1_delay_4_44;
  reg                 io_A_Valid_1_delay_5_43;
  reg                 io_A_Valid_1_delay_6_42;
  reg                 io_A_Valid_1_delay_7_41;
  reg                 io_A_Valid_1_delay_8_40;
  reg                 io_A_Valid_1_delay_9_39;
  reg                 io_A_Valid_1_delay_10_38;
  reg                 io_A_Valid_1_delay_11_37;
  reg                 io_A_Valid_1_delay_12_36;
  reg                 io_A_Valid_1_delay_13_35;
  reg                 io_A_Valid_1_delay_14_34;
  reg                 io_A_Valid_1_delay_15_33;
  reg                 io_A_Valid_1_delay_16_32;
  reg                 io_A_Valid_1_delay_17_31;
  reg                 io_A_Valid_1_delay_18_30;
  reg                 io_A_Valid_1_delay_19_29;
  reg                 io_A_Valid_1_delay_20_28;
  reg                 io_A_Valid_1_delay_21_27;
  reg                 io_A_Valid_1_delay_22_26;
  reg                 io_A_Valid_1_delay_23_25;
  reg                 io_A_Valid_1_delay_24_24;
  reg                 io_A_Valid_1_delay_25_23;
  reg                 io_A_Valid_1_delay_26_22;
  reg                 io_A_Valid_1_delay_27_21;
  reg                 io_A_Valid_1_delay_28_20;
  reg                 io_A_Valid_1_delay_29_19;
  reg                 io_A_Valid_1_delay_30_18;
  reg                 io_A_Valid_1_delay_31_17;
  reg                 io_A_Valid_1_delay_32_16;
  reg                 io_A_Valid_1_delay_33_15;
  reg                 io_A_Valid_1_delay_34_14;
  reg                 io_A_Valid_1_delay_35_13;
  reg                 io_A_Valid_1_delay_36_12;
  reg                 io_A_Valid_1_delay_37_11;
  reg                 io_A_Valid_1_delay_38_10;
  reg                 io_A_Valid_1_delay_39_9;
  reg                 io_A_Valid_1_delay_40_8;
  reg                 io_A_Valid_1_delay_41_7;
  reg                 io_A_Valid_1_delay_42_6;
  reg                 io_A_Valid_1_delay_43_5;
  reg                 io_A_Valid_1_delay_44_4;
  reg                 io_A_Valid_1_delay_45_3;
  reg                 io_A_Valid_1_delay_46_2;
  reg                 io_A_Valid_1_delay_47_1;
  reg                 io_A_Valid_1_delay_48;
  reg                 io_B_Valid_48_delay_1;
  reg                 io_A_Valid_1_delay_1_48;
  reg                 io_A_Valid_1_delay_2_47;
  reg                 io_A_Valid_1_delay_3_46;
  reg                 io_A_Valid_1_delay_4_45;
  reg                 io_A_Valid_1_delay_5_44;
  reg                 io_A_Valid_1_delay_6_43;
  reg                 io_A_Valid_1_delay_7_42;
  reg                 io_A_Valid_1_delay_8_41;
  reg                 io_A_Valid_1_delay_9_40;
  reg                 io_A_Valid_1_delay_10_39;
  reg                 io_A_Valid_1_delay_11_38;
  reg                 io_A_Valid_1_delay_12_37;
  reg                 io_A_Valid_1_delay_13_36;
  reg                 io_A_Valid_1_delay_14_35;
  reg                 io_A_Valid_1_delay_15_34;
  reg                 io_A_Valid_1_delay_16_33;
  reg                 io_A_Valid_1_delay_17_32;
  reg                 io_A_Valid_1_delay_18_31;
  reg                 io_A_Valid_1_delay_19_30;
  reg                 io_A_Valid_1_delay_20_29;
  reg                 io_A_Valid_1_delay_21_28;
  reg                 io_A_Valid_1_delay_22_27;
  reg                 io_A_Valid_1_delay_23_26;
  reg                 io_A_Valid_1_delay_24_25;
  reg                 io_A_Valid_1_delay_25_24;
  reg                 io_A_Valid_1_delay_26_23;
  reg                 io_A_Valid_1_delay_27_22;
  reg                 io_A_Valid_1_delay_28_21;
  reg                 io_A_Valid_1_delay_29_20;
  reg                 io_A_Valid_1_delay_30_19;
  reg                 io_A_Valid_1_delay_31_18;
  reg                 io_A_Valid_1_delay_32_17;
  reg                 io_A_Valid_1_delay_33_16;
  reg                 io_A_Valid_1_delay_34_15;
  reg                 io_A_Valid_1_delay_35_14;
  reg                 io_A_Valid_1_delay_36_13;
  reg                 io_A_Valid_1_delay_37_12;
  reg                 io_A_Valid_1_delay_38_11;
  reg                 io_A_Valid_1_delay_39_10;
  reg                 io_A_Valid_1_delay_40_9;
  reg                 io_A_Valid_1_delay_41_8;
  reg                 io_A_Valid_1_delay_42_7;
  reg                 io_A_Valid_1_delay_43_6;
  reg                 io_A_Valid_1_delay_44_5;
  reg                 io_A_Valid_1_delay_45_4;
  reg                 io_A_Valid_1_delay_46_3;
  reg                 io_A_Valid_1_delay_47_2;
  reg                 io_A_Valid_1_delay_48_1;
  reg                 io_A_Valid_1_delay_49;
  reg                 io_B_Valid_49_delay_1;
  reg                 io_A_Valid_1_delay_1_49;
  reg                 io_A_Valid_1_delay_2_48;
  reg                 io_A_Valid_1_delay_3_47;
  reg                 io_A_Valid_1_delay_4_46;
  reg                 io_A_Valid_1_delay_5_45;
  reg                 io_A_Valid_1_delay_6_44;
  reg                 io_A_Valid_1_delay_7_43;
  reg                 io_A_Valid_1_delay_8_42;
  reg                 io_A_Valid_1_delay_9_41;
  reg                 io_A_Valid_1_delay_10_40;
  reg                 io_A_Valid_1_delay_11_39;
  reg                 io_A_Valid_1_delay_12_38;
  reg                 io_A_Valid_1_delay_13_37;
  reg                 io_A_Valid_1_delay_14_36;
  reg                 io_A_Valid_1_delay_15_35;
  reg                 io_A_Valid_1_delay_16_34;
  reg                 io_A_Valid_1_delay_17_33;
  reg                 io_A_Valid_1_delay_18_32;
  reg                 io_A_Valid_1_delay_19_31;
  reg                 io_A_Valid_1_delay_20_30;
  reg                 io_A_Valid_1_delay_21_29;
  reg                 io_A_Valid_1_delay_22_28;
  reg                 io_A_Valid_1_delay_23_27;
  reg                 io_A_Valid_1_delay_24_26;
  reg                 io_A_Valid_1_delay_25_25;
  reg                 io_A_Valid_1_delay_26_24;
  reg                 io_A_Valid_1_delay_27_23;
  reg                 io_A_Valid_1_delay_28_22;
  reg                 io_A_Valid_1_delay_29_21;
  reg                 io_A_Valid_1_delay_30_20;
  reg                 io_A_Valid_1_delay_31_19;
  reg                 io_A_Valid_1_delay_32_18;
  reg                 io_A_Valid_1_delay_33_17;
  reg                 io_A_Valid_1_delay_34_16;
  reg                 io_A_Valid_1_delay_35_15;
  reg                 io_A_Valid_1_delay_36_14;
  reg                 io_A_Valid_1_delay_37_13;
  reg                 io_A_Valid_1_delay_38_12;
  reg                 io_A_Valid_1_delay_39_11;
  reg                 io_A_Valid_1_delay_40_10;
  reg                 io_A_Valid_1_delay_41_9;
  reg                 io_A_Valid_1_delay_42_8;
  reg                 io_A_Valid_1_delay_43_7;
  reg                 io_A_Valid_1_delay_44_6;
  reg                 io_A_Valid_1_delay_45_5;
  reg                 io_A_Valid_1_delay_46_4;
  reg                 io_A_Valid_1_delay_47_3;
  reg                 io_A_Valid_1_delay_48_2;
  reg                 io_A_Valid_1_delay_49_1;
  reg                 io_A_Valid_1_delay_50;
  reg                 io_B_Valid_50_delay_1;
  reg                 io_A_Valid_1_delay_1_50;
  reg                 io_A_Valid_1_delay_2_49;
  reg                 io_A_Valid_1_delay_3_48;
  reg                 io_A_Valid_1_delay_4_47;
  reg                 io_A_Valid_1_delay_5_46;
  reg                 io_A_Valid_1_delay_6_45;
  reg                 io_A_Valid_1_delay_7_44;
  reg                 io_A_Valid_1_delay_8_43;
  reg                 io_A_Valid_1_delay_9_42;
  reg                 io_A_Valid_1_delay_10_41;
  reg                 io_A_Valid_1_delay_11_40;
  reg                 io_A_Valid_1_delay_12_39;
  reg                 io_A_Valid_1_delay_13_38;
  reg                 io_A_Valid_1_delay_14_37;
  reg                 io_A_Valid_1_delay_15_36;
  reg                 io_A_Valid_1_delay_16_35;
  reg                 io_A_Valid_1_delay_17_34;
  reg                 io_A_Valid_1_delay_18_33;
  reg                 io_A_Valid_1_delay_19_32;
  reg                 io_A_Valid_1_delay_20_31;
  reg                 io_A_Valid_1_delay_21_30;
  reg                 io_A_Valid_1_delay_22_29;
  reg                 io_A_Valid_1_delay_23_28;
  reg                 io_A_Valid_1_delay_24_27;
  reg                 io_A_Valid_1_delay_25_26;
  reg                 io_A_Valid_1_delay_26_25;
  reg                 io_A_Valid_1_delay_27_24;
  reg                 io_A_Valid_1_delay_28_23;
  reg                 io_A_Valid_1_delay_29_22;
  reg                 io_A_Valid_1_delay_30_21;
  reg                 io_A_Valid_1_delay_31_20;
  reg                 io_A_Valid_1_delay_32_19;
  reg                 io_A_Valid_1_delay_33_18;
  reg                 io_A_Valid_1_delay_34_17;
  reg                 io_A_Valid_1_delay_35_16;
  reg                 io_A_Valid_1_delay_36_15;
  reg                 io_A_Valid_1_delay_37_14;
  reg                 io_A_Valid_1_delay_38_13;
  reg                 io_A_Valid_1_delay_39_12;
  reg                 io_A_Valid_1_delay_40_11;
  reg                 io_A_Valid_1_delay_41_10;
  reg                 io_A_Valid_1_delay_42_9;
  reg                 io_A_Valid_1_delay_43_8;
  reg                 io_A_Valid_1_delay_44_7;
  reg                 io_A_Valid_1_delay_45_6;
  reg                 io_A_Valid_1_delay_46_5;
  reg                 io_A_Valid_1_delay_47_4;
  reg                 io_A_Valid_1_delay_48_3;
  reg                 io_A_Valid_1_delay_49_2;
  reg                 io_A_Valid_1_delay_50_1;
  reg                 io_A_Valid_1_delay_51;
  reg                 io_B_Valid_51_delay_1;
  reg                 io_A_Valid_1_delay_1_51;
  reg                 io_A_Valid_1_delay_2_50;
  reg                 io_A_Valid_1_delay_3_49;
  reg                 io_A_Valid_1_delay_4_48;
  reg                 io_A_Valid_1_delay_5_47;
  reg                 io_A_Valid_1_delay_6_46;
  reg                 io_A_Valid_1_delay_7_45;
  reg                 io_A_Valid_1_delay_8_44;
  reg                 io_A_Valid_1_delay_9_43;
  reg                 io_A_Valid_1_delay_10_42;
  reg                 io_A_Valid_1_delay_11_41;
  reg                 io_A_Valid_1_delay_12_40;
  reg                 io_A_Valid_1_delay_13_39;
  reg                 io_A_Valid_1_delay_14_38;
  reg                 io_A_Valid_1_delay_15_37;
  reg                 io_A_Valid_1_delay_16_36;
  reg                 io_A_Valid_1_delay_17_35;
  reg                 io_A_Valid_1_delay_18_34;
  reg                 io_A_Valid_1_delay_19_33;
  reg                 io_A_Valid_1_delay_20_32;
  reg                 io_A_Valid_1_delay_21_31;
  reg                 io_A_Valid_1_delay_22_30;
  reg                 io_A_Valid_1_delay_23_29;
  reg                 io_A_Valid_1_delay_24_28;
  reg                 io_A_Valid_1_delay_25_27;
  reg                 io_A_Valid_1_delay_26_26;
  reg                 io_A_Valid_1_delay_27_25;
  reg                 io_A_Valid_1_delay_28_24;
  reg                 io_A_Valid_1_delay_29_23;
  reg                 io_A_Valid_1_delay_30_22;
  reg                 io_A_Valid_1_delay_31_21;
  reg                 io_A_Valid_1_delay_32_20;
  reg                 io_A_Valid_1_delay_33_19;
  reg                 io_A_Valid_1_delay_34_18;
  reg                 io_A_Valid_1_delay_35_17;
  reg                 io_A_Valid_1_delay_36_16;
  reg                 io_A_Valid_1_delay_37_15;
  reg                 io_A_Valid_1_delay_38_14;
  reg                 io_A_Valid_1_delay_39_13;
  reg                 io_A_Valid_1_delay_40_12;
  reg                 io_A_Valid_1_delay_41_11;
  reg                 io_A_Valid_1_delay_42_10;
  reg                 io_A_Valid_1_delay_43_9;
  reg                 io_A_Valid_1_delay_44_8;
  reg                 io_A_Valid_1_delay_45_7;
  reg                 io_A_Valid_1_delay_46_6;
  reg                 io_A_Valid_1_delay_47_5;
  reg                 io_A_Valid_1_delay_48_4;
  reg                 io_A_Valid_1_delay_49_3;
  reg                 io_A_Valid_1_delay_50_2;
  reg                 io_A_Valid_1_delay_51_1;
  reg                 io_A_Valid_1_delay_52;
  reg                 io_B_Valid_52_delay_1;
  reg                 io_A_Valid_1_delay_1_52;
  reg                 io_A_Valid_1_delay_2_51;
  reg                 io_A_Valid_1_delay_3_50;
  reg                 io_A_Valid_1_delay_4_49;
  reg                 io_A_Valid_1_delay_5_48;
  reg                 io_A_Valid_1_delay_6_47;
  reg                 io_A_Valid_1_delay_7_46;
  reg                 io_A_Valid_1_delay_8_45;
  reg                 io_A_Valid_1_delay_9_44;
  reg                 io_A_Valid_1_delay_10_43;
  reg                 io_A_Valid_1_delay_11_42;
  reg                 io_A_Valid_1_delay_12_41;
  reg                 io_A_Valid_1_delay_13_40;
  reg                 io_A_Valid_1_delay_14_39;
  reg                 io_A_Valid_1_delay_15_38;
  reg                 io_A_Valid_1_delay_16_37;
  reg                 io_A_Valid_1_delay_17_36;
  reg                 io_A_Valid_1_delay_18_35;
  reg                 io_A_Valid_1_delay_19_34;
  reg                 io_A_Valid_1_delay_20_33;
  reg                 io_A_Valid_1_delay_21_32;
  reg                 io_A_Valid_1_delay_22_31;
  reg                 io_A_Valid_1_delay_23_30;
  reg                 io_A_Valid_1_delay_24_29;
  reg                 io_A_Valid_1_delay_25_28;
  reg                 io_A_Valid_1_delay_26_27;
  reg                 io_A_Valid_1_delay_27_26;
  reg                 io_A_Valid_1_delay_28_25;
  reg                 io_A_Valid_1_delay_29_24;
  reg                 io_A_Valid_1_delay_30_23;
  reg                 io_A_Valid_1_delay_31_22;
  reg                 io_A_Valid_1_delay_32_21;
  reg                 io_A_Valid_1_delay_33_20;
  reg                 io_A_Valid_1_delay_34_19;
  reg                 io_A_Valid_1_delay_35_18;
  reg                 io_A_Valid_1_delay_36_17;
  reg                 io_A_Valid_1_delay_37_16;
  reg                 io_A_Valid_1_delay_38_15;
  reg                 io_A_Valid_1_delay_39_14;
  reg                 io_A_Valid_1_delay_40_13;
  reg                 io_A_Valid_1_delay_41_12;
  reg                 io_A_Valid_1_delay_42_11;
  reg                 io_A_Valid_1_delay_43_10;
  reg                 io_A_Valid_1_delay_44_9;
  reg                 io_A_Valid_1_delay_45_8;
  reg                 io_A_Valid_1_delay_46_7;
  reg                 io_A_Valid_1_delay_47_6;
  reg                 io_A_Valid_1_delay_48_5;
  reg                 io_A_Valid_1_delay_49_4;
  reg                 io_A_Valid_1_delay_50_3;
  reg                 io_A_Valid_1_delay_51_2;
  reg                 io_A_Valid_1_delay_52_1;
  reg                 io_A_Valid_1_delay_53;
  reg                 io_B_Valid_53_delay_1;
  reg                 io_A_Valid_1_delay_1_53;
  reg                 io_A_Valid_1_delay_2_52;
  reg                 io_A_Valid_1_delay_3_51;
  reg                 io_A_Valid_1_delay_4_50;
  reg                 io_A_Valid_1_delay_5_49;
  reg                 io_A_Valid_1_delay_6_48;
  reg                 io_A_Valid_1_delay_7_47;
  reg                 io_A_Valid_1_delay_8_46;
  reg                 io_A_Valid_1_delay_9_45;
  reg                 io_A_Valid_1_delay_10_44;
  reg                 io_A_Valid_1_delay_11_43;
  reg                 io_A_Valid_1_delay_12_42;
  reg                 io_A_Valid_1_delay_13_41;
  reg                 io_A_Valid_1_delay_14_40;
  reg                 io_A_Valid_1_delay_15_39;
  reg                 io_A_Valid_1_delay_16_38;
  reg                 io_A_Valid_1_delay_17_37;
  reg                 io_A_Valid_1_delay_18_36;
  reg                 io_A_Valid_1_delay_19_35;
  reg                 io_A_Valid_1_delay_20_34;
  reg                 io_A_Valid_1_delay_21_33;
  reg                 io_A_Valid_1_delay_22_32;
  reg                 io_A_Valid_1_delay_23_31;
  reg                 io_A_Valid_1_delay_24_30;
  reg                 io_A_Valid_1_delay_25_29;
  reg                 io_A_Valid_1_delay_26_28;
  reg                 io_A_Valid_1_delay_27_27;
  reg                 io_A_Valid_1_delay_28_26;
  reg                 io_A_Valid_1_delay_29_25;
  reg                 io_A_Valid_1_delay_30_24;
  reg                 io_A_Valid_1_delay_31_23;
  reg                 io_A_Valid_1_delay_32_22;
  reg                 io_A_Valid_1_delay_33_21;
  reg                 io_A_Valid_1_delay_34_20;
  reg                 io_A_Valid_1_delay_35_19;
  reg                 io_A_Valid_1_delay_36_18;
  reg                 io_A_Valid_1_delay_37_17;
  reg                 io_A_Valid_1_delay_38_16;
  reg                 io_A_Valid_1_delay_39_15;
  reg                 io_A_Valid_1_delay_40_14;
  reg                 io_A_Valid_1_delay_41_13;
  reg                 io_A_Valid_1_delay_42_12;
  reg                 io_A_Valid_1_delay_43_11;
  reg                 io_A_Valid_1_delay_44_10;
  reg                 io_A_Valid_1_delay_45_9;
  reg                 io_A_Valid_1_delay_46_8;
  reg                 io_A_Valid_1_delay_47_7;
  reg                 io_A_Valid_1_delay_48_6;
  reg                 io_A_Valid_1_delay_49_5;
  reg                 io_A_Valid_1_delay_50_4;
  reg                 io_A_Valid_1_delay_51_3;
  reg                 io_A_Valid_1_delay_52_2;
  reg                 io_A_Valid_1_delay_53_1;
  reg                 io_A_Valid_1_delay_54;
  reg                 io_B_Valid_54_delay_1;
  reg                 io_A_Valid_1_delay_1_54;
  reg                 io_A_Valid_1_delay_2_53;
  reg                 io_A_Valid_1_delay_3_52;
  reg                 io_A_Valid_1_delay_4_51;
  reg                 io_A_Valid_1_delay_5_50;
  reg                 io_A_Valid_1_delay_6_49;
  reg                 io_A_Valid_1_delay_7_48;
  reg                 io_A_Valid_1_delay_8_47;
  reg                 io_A_Valid_1_delay_9_46;
  reg                 io_A_Valid_1_delay_10_45;
  reg                 io_A_Valid_1_delay_11_44;
  reg                 io_A_Valid_1_delay_12_43;
  reg                 io_A_Valid_1_delay_13_42;
  reg                 io_A_Valid_1_delay_14_41;
  reg                 io_A_Valid_1_delay_15_40;
  reg                 io_A_Valid_1_delay_16_39;
  reg                 io_A_Valid_1_delay_17_38;
  reg                 io_A_Valid_1_delay_18_37;
  reg                 io_A_Valid_1_delay_19_36;
  reg                 io_A_Valid_1_delay_20_35;
  reg                 io_A_Valid_1_delay_21_34;
  reg                 io_A_Valid_1_delay_22_33;
  reg                 io_A_Valid_1_delay_23_32;
  reg                 io_A_Valid_1_delay_24_31;
  reg                 io_A_Valid_1_delay_25_30;
  reg                 io_A_Valid_1_delay_26_29;
  reg                 io_A_Valid_1_delay_27_28;
  reg                 io_A_Valid_1_delay_28_27;
  reg                 io_A_Valid_1_delay_29_26;
  reg                 io_A_Valid_1_delay_30_25;
  reg                 io_A_Valid_1_delay_31_24;
  reg                 io_A_Valid_1_delay_32_23;
  reg                 io_A_Valid_1_delay_33_22;
  reg                 io_A_Valid_1_delay_34_21;
  reg                 io_A_Valid_1_delay_35_20;
  reg                 io_A_Valid_1_delay_36_19;
  reg                 io_A_Valid_1_delay_37_18;
  reg                 io_A_Valid_1_delay_38_17;
  reg                 io_A_Valid_1_delay_39_16;
  reg                 io_A_Valid_1_delay_40_15;
  reg                 io_A_Valid_1_delay_41_14;
  reg                 io_A_Valid_1_delay_42_13;
  reg                 io_A_Valid_1_delay_43_12;
  reg                 io_A_Valid_1_delay_44_11;
  reg                 io_A_Valid_1_delay_45_10;
  reg                 io_A_Valid_1_delay_46_9;
  reg                 io_A_Valid_1_delay_47_8;
  reg                 io_A_Valid_1_delay_48_7;
  reg                 io_A_Valid_1_delay_49_6;
  reg                 io_A_Valid_1_delay_50_5;
  reg                 io_A_Valid_1_delay_51_4;
  reg                 io_A_Valid_1_delay_52_3;
  reg                 io_A_Valid_1_delay_53_2;
  reg                 io_A_Valid_1_delay_54_1;
  reg                 io_A_Valid_1_delay_55;
  reg                 io_B_Valid_55_delay_1;
  reg                 io_A_Valid_1_delay_1_55;
  reg                 io_A_Valid_1_delay_2_54;
  reg                 io_A_Valid_1_delay_3_53;
  reg                 io_A_Valid_1_delay_4_52;
  reg                 io_A_Valid_1_delay_5_51;
  reg                 io_A_Valid_1_delay_6_50;
  reg                 io_A_Valid_1_delay_7_49;
  reg                 io_A_Valid_1_delay_8_48;
  reg                 io_A_Valid_1_delay_9_47;
  reg                 io_A_Valid_1_delay_10_46;
  reg                 io_A_Valid_1_delay_11_45;
  reg                 io_A_Valid_1_delay_12_44;
  reg                 io_A_Valid_1_delay_13_43;
  reg                 io_A_Valid_1_delay_14_42;
  reg                 io_A_Valid_1_delay_15_41;
  reg                 io_A_Valid_1_delay_16_40;
  reg                 io_A_Valid_1_delay_17_39;
  reg                 io_A_Valid_1_delay_18_38;
  reg                 io_A_Valid_1_delay_19_37;
  reg                 io_A_Valid_1_delay_20_36;
  reg                 io_A_Valid_1_delay_21_35;
  reg                 io_A_Valid_1_delay_22_34;
  reg                 io_A_Valid_1_delay_23_33;
  reg                 io_A_Valid_1_delay_24_32;
  reg                 io_A_Valid_1_delay_25_31;
  reg                 io_A_Valid_1_delay_26_30;
  reg                 io_A_Valid_1_delay_27_29;
  reg                 io_A_Valid_1_delay_28_28;
  reg                 io_A_Valid_1_delay_29_27;
  reg                 io_A_Valid_1_delay_30_26;
  reg                 io_A_Valid_1_delay_31_25;
  reg                 io_A_Valid_1_delay_32_24;
  reg                 io_A_Valid_1_delay_33_23;
  reg                 io_A_Valid_1_delay_34_22;
  reg                 io_A_Valid_1_delay_35_21;
  reg                 io_A_Valid_1_delay_36_20;
  reg                 io_A_Valid_1_delay_37_19;
  reg                 io_A_Valid_1_delay_38_18;
  reg                 io_A_Valid_1_delay_39_17;
  reg                 io_A_Valid_1_delay_40_16;
  reg                 io_A_Valid_1_delay_41_15;
  reg                 io_A_Valid_1_delay_42_14;
  reg                 io_A_Valid_1_delay_43_13;
  reg                 io_A_Valid_1_delay_44_12;
  reg                 io_A_Valid_1_delay_45_11;
  reg                 io_A_Valid_1_delay_46_10;
  reg                 io_A_Valid_1_delay_47_9;
  reg                 io_A_Valid_1_delay_48_8;
  reg                 io_A_Valid_1_delay_49_7;
  reg                 io_A_Valid_1_delay_50_6;
  reg                 io_A_Valid_1_delay_51_5;
  reg                 io_A_Valid_1_delay_52_4;
  reg                 io_A_Valid_1_delay_53_3;
  reg                 io_A_Valid_1_delay_54_2;
  reg                 io_A_Valid_1_delay_55_1;
  reg                 io_A_Valid_1_delay_56;
  reg                 io_B_Valid_56_delay_1;
  reg                 io_A_Valid_1_delay_1_56;
  reg                 io_A_Valid_1_delay_2_55;
  reg                 io_A_Valid_1_delay_3_54;
  reg                 io_A_Valid_1_delay_4_53;
  reg                 io_A_Valid_1_delay_5_52;
  reg                 io_A_Valid_1_delay_6_51;
  reg                 io_A_Valid_1_delay_7_50;
  reg                 io_A_Valid_1_delay_8_49;
  reg                 io_A_Valid_1_delay_9_48;
  reg                 io_A_Valid_1_delay_10_47;
  reg                 io_A_Valid_1_delay_11_46;
  reg                 io_A_Valid_1_delay_12_45;
  reg                 io_A_Valid_1_delay_13_44;
  reg                 io_A_Valid_1_delay_14_43;
  reg                 io_A_Valid_1_delay_15_42;
  reg                 io_A_Valid_1_delay_16_41;
  reg                 io_A_Valid_1_delay_17_40;
  reg                 io_A_Valid_1_delay_18_39;
  reg                 io_A_Valid_1_delay_19_38;
  reg                 io_A_Valid_1_delay_20_37;
  reg                 io_A_Valid_1_delay_21_36;
  reg                 io_A_Valid_1_delay_22_35;
  reg                 io_A_Valid_1_delay_23_34;
  reg                 io_A_Valid_1_delay_24_33;
  reg                 io_A_Valid_1_delay_25_32;
  reg                 io_A_Valid_1_delay_26_31;
  reg                 io_A_Valid_1_delay_27_30;
  reg                 io_A_Valid_1_delay_28_29;
  reg                 io_A_Valid_1_delay_29_28;
  reg                 io_A_Valid_1_delay_30_27;
  reg                 io_A_Valid_1_delay_31_26;
  reg                 io_A_Valid_1_delay_32_25;
  reg                 io_A_Valid_1_delay_33_24;
  reg                 io_A_Valid_1_delay_34_23;
  reg                 io_A_Valid_1_delay_35_22;
  reg                 io_A_Valid_1_delay_36_21;
  reg                 io_A_Valid_1_delay_37_20;
  reg                 io_A_Valid_1_delay_38_19;
  reg                 io_A_Valid_1_delay_39_18;
  reg                 io_A_Valid_1_delay_40_17;
  reg                 io_A_Valid_1_delay_41_16;
  reg                 io_A_Valid_1_delay_42_15;
  reg                 io_A_Valid_1_delay_43_14;
  reg                 io_A_Valid_1_delay_44_13;
  reg                 io_A_Valid_1_delay_45_12;
  reg                 io_A_Valid_1_delay_46_11;
  reg                 io_A_Valid_1_delay_47_10;
  reg                 io_A_Valid_1_delay_48_9;
  reg                 io_A_Valid_1_delay_49_8;
  reg                 io_A_Valid_1_delay_50_7;
  reg                 io_A_Valid_1_delay_51_6;
  reg                 io_A_Valid_1_delay_52_5;
  reg                 io_A_Valid_1_delay_53_4;
  reg                 io_A_Valid_1_delay_54_3;
  reg                 io_A_Valid_1_delay_55_2;
  reg                 io_A_Valid_1_delay_56_1;
  reg                 io_A_Valid_1_delay_57;
  reg                 io_B_Valid_57_delay_1;
  reg                 io_A_Valid_1_delay_1_57;
  reg                 io_A_Valid_1_delay_2_56;
  reg                 io_A_Valid_1_delay_3_55;
  reg                 io_A_Valid_1_delay_4_54;
  reg                 io_A_Valid_1_delay_5_53;
  reg                 io_A_Valid_1_delay_6_52;
  reg                 io_A_Valid_1_delay_7_51;
  reg                 io_A_Valid_1_delay_8_50;
  reg                 io_A_Valid_1_delay_9_49;
  reg                 io_A_Valid_1_delay_10_48;
  reg                 io_A_Valid_1_delay_11_47;
  reg                 io_A_Valid_1_delay_12_46;
  reg                 io_A_Valid_1_delay_13_45;
  reg                 io_A_Valid_1_delay_14_44;
  reg                 io_A_Valid_1_delay_15_43;
  reg                 io_A_Valid_1_delay_16_42;
  reg                 io_A_Valid_1_delay_17_41;
  reg                 io_A_Valid_1_delay_18_40;
  reg                 io_A_Valid_1_delay_19_39;
  reg                 io_A_Valid_1_delay_20_38;
  reg                 io_A_Valid_1_delay_21_37;
  reg                 io_A_Valid_1_delay_22_36;
  reg                 io_A_Valid_1_delay_23_35;
  reg                 io_A_Valid_1_delay_24_34;
  reg                 io_A_Valid_1_delay_25_33;
  reg                 io_A_Valid_1_delay_26_32;
  reg                 io_A_Valid_1_delay_27_31;
  reg                 io_A_Valid_1_delay_28_30;
  reg                 io_A_Valid_1_delay_29_29;
  reg                 io_A_Valid_1_delay_30_28;
  reg                 io_A_Valid_1_delay_31_27;
  reg                 io_A_Valid_1_delay_32_26;
  reg                 io_A_Valid_1_delay_33_25;
  reg                 io_A_Valid_1_delay_34_24;
  reg                 io_A_Valid_1_delay_35_23;
  reg                 io_A_Valid_1_delay_36_22;
  reg                 io_A_Valid_1_delay_37_21;
  reg                 io_A_Valid_1_delay_38_20;
  reg                 io_A_Valid_1_delay_39_19;
  reg                 io_A_Valid_1_delay_40_18;
  reg                 io_A_Valid_1_delay_41_17;
  reg                 io_A_Valid_1_delay_42_16;
  reg                 io_A_Valid_1_delay_43_15;
  reg                 io_A_Valid_1_delay_44_14;
  reg                 io_A_Valid_1_delay_45_13;
  reg                 io_A_Valid_1_delay_46_12;
  reg                 io_A_Valid_1_delay_47_11;
  reg                 io_A_Valid_1_delay_48_10;
  reg                 io_A_Valid_1_delay_49_9;
  reg                 io_A_Valid_1_delay_50_8;
  reg                 io_A_Valid_1_delay_51_7;
  reg                 io_A_Valid_1_delay_52_6;
  reg                 io_A_Valid_1_delay_53_5;
  reg                 io_A_Valid_1_delay_54_4;
  reg                 io_A_Valid_1_delay_55_3;
  reg                 io_A_Valid_1_delay_56_2;
  reg                 io_A_Valid_1_delay_57_1;
  reg                 io_A_Valid_1_delay_58;
  reg                 io_B_Valid_58_delay_1;
  reg                 io_A_Valid_1_delay_1_58;
  reg                 io_A_Valid_1_delay_2_57;
  reg                 io_A_Valid_1_delay_3_56;
  reg                 io_A_Valid_1_delay_4_55;
  reg                 io_A_Valid_1_delay_5_54;
  reg                 io_A_Valid_1_delay_6_53;
  reg                 io_A_Valid_1_delay_7_52;
  reg                 io_A_Valid_1_delay_8_51;
  reg                 io_A_Valid_1_delay_9_50;
  reg                 io_A_Valid_1_delay_10_49;
  reg                 io_A_Valid_1_delay_11_48;
  reg                 io_A_Valid_1_delay_12_47;
  reg                 io_A_Valid_1_delay_13_46;
  reg                 io_A_Valid_1_delay_14_45;
  reg                 io_A_Valid_1_delay_15_44;
  reg                 io_A_Valid_1_delay_16_43;
  reg                 io_A_Valid_1_delay_17_42;
  reg                 io_A_Valid_1_delay_18_41;
  reg                 io_A_Valid_1_delay_19_40;
  reg                 io_A_Valid_1_delay_20_39;
  reg                 io_A_Valid_1_delay_21_38;
  reg                 io_A_Valid_1_delay_22_37;
  reg                 io_A_Valid_1_delay_23_36;
  reg                 io_A_Valid_1_delay_24_35;
  reg                 io_A_Valid_1_delay_25_34;
  reg                 io_A_Valid_1_delay_26_33;
  reg                 io_A_Valid_1_delay_27_32;
  reg                 io_A_Valid_1_delay_28_31;
  reg                 io_A_Valid_1_delay_29_30;
  reg                 io_A_Valid_1_delay_30_29;
  reg                 io_A_Valid_1_delay_31_28;
  reg                 io_A_Valid_1_delay_32_27;
  reg                 io_A_Valid_1_delay_33_26;
  reg                 io_A_Valid_1_delay_34_25;
  reg                 io_A_Valid_1_delay_35_24;
  reg                 io_A_Valid_1_delay_36_23;
  reg                 io_A_Valid_1_delay_37_22;
  reg                 io_A_Valid_1_delay_38_21;
  reg                 io_A_Valid_1_delay_39_20;
  reg                 io_A_Valid_1_delay_40_19;
  reg                 io_A_Valid_1_delay_41_18;
  reg                 io_A_Valid_1_delay_42_17;
  reg                 io_A_Valid_1_delay_43_16;
  reg                 io_A_Valid_1_delay_44_15;
  reg                 io_A_Valid_1_delay_45_14;
  reg                 io_A_Valid_1_delay_46_13;
  reg                 io_A_Valid_1_delay_47_12;
  reg                 io_A_Valid_1_delay_48_11;
  reg                 io_A_Valid_1_delay_49_10;
  reg                 io_A_Valid_1_delay_50_9;
  reg                 io_A_Valid_1_delay_51_8;
  reg                 io_A_Valid_1_delay_52_7;
  reg                 io_A_Valid_1_delay_53_6;
  reg                 io_A_Valid_1_delay_54_5;
  reg                 io_A_Valid_1_delay_55_4;
  reg                 io_A_Valid_1_delay_56_3;
  reg                 io_A_Valid_1_delay_57_2;
  reg                 io_A_Valid_1_delay_58_1;
  reg                 io_A_Valid_1_delay_59;
  reg                 io_B_Valid_59_delay_1;
  reg                 io_A_Valid_1_delay_1_59;
  reg                 io_A_Valid_1_delay_2_58;
  reg                 io_A_Valid_1_delay_3_57;
  reg                 io_A_Valid_1_delay_4_56;
  reg                 io_A_Valid_1_delay_5_55;
  reg                 io_A_Valid_1_delay_6_54;
  reg                 io_A_Valid_1_delay_7_53;
  reg                 io_A_Valid_1_delay_8_52;
  reg                 io_A_Valid_1_delay_9_51;
  reg                 io_A_Valid_1_delay_10_50;
  reg                 io_A_Valid_1_delay_11_49;
  reg                 io_A_Valid_1_delay_12_48;
  reg                 io_A_Valid_1_delay_13_47;
  reg                 io_A_Valid_1_delay_14_46;
  reg                 io_A_Valid_1_delay_15_45;
  reg                 io_A_Valid_1_delay_16_44;
  reg                 io_A_Valid_1_delay_17_43;
  reg                 io_A_Valid_1_delay_18_42;
  reg                 io_A_Valid_1_delay_19_41;
  reg                 io_A_Valid_1_delay_20_40;
  reg                 io_A_Valid_1_delay_21_39;
  reg                 io_A_Valid_1_delay_22_38;
  reg                 io_A_Valid_1_delay_23_37;
  reg                 io_A_Valid_1_delay_24_36;
  reg                 io_A_Valid_1_delay_25_35;
  reg                 io_A_Valid_1_delay_26_34;
  reg                 io_A_Valid_1_delay_27_33;
  reg                 io_A_Valid_1_delay_28_32;
  reg                 io_A_Valid_1_delay_29_31;
  reg                 io_A_Valid_1_delay_30_30;
  reg                 io_A_Valid_1_delay_31_29;
  reg                 io_A_Valid_1_delay_32_28;
  reg                 io_A_Valid_1_delay_33_27;
  reg                 io_A_Valid_1_delay_34_26;
  reg                 io_A_Valid_1_delay_35_25;
  reg                 io_A_Valid_1_delay_36_24;
  reg                 io_A_Valid_1_delay_37_23;
  reg                 io_A_Valid_1_delay_38_22;
  reg                 io_A_Valid_1_delay_39_21;
  reg                 io_A_Valid_1_delay_40_20;
  reg                 io_A_Valid_1_delay_41_19;
  reg                 io_A_Valid_1_delay_42_18;
  reg                 io_A_Valid_1_delay_43_17;
  reg                 io_A_Valid_1_delay_44_16;
  reg                 io_A_Valid_1_delay_45_15;
  reg                 io_A_Valid_1_delay_46_14;
  reg                 io_A_Valid_1_delay_47_13;
  reg                 io_A_Valid_1_delay_48_12;
  reg                 io_A_Valid_1_delay_49_11;
  reg                 io_A_Valid_1_delay_50_10;
  reg                 io_A_Valid_1_delay_51_9;
  reg                 io_A_Valid_1_delay_52_8;
  reg                 io_A_Valid_1_delay_53_7;
  reg                 io_A_Valid_1_delay_54_6;
  reg                 io_A_Valid_1_delay_55_5;
  reg                 io_A_Valid_1_delay_56_4;
  reg                 io_A_Valid_1_delay_57_3;
  reg                 io_A_Valid_1_delay_58_2;
  reg                 io_A_Valid_1_delay_59_1;
  reg                 io_A_Valid_1_delay_60;
  reg                 io_B_Valid_60_delay_1;
  reg                 io_A_Valid_1_delay_1_60;
  reg                 io_A_Valid_1_delay_2_59;
  reg                 io_A_Valid_1_delay_3_58;
  reg                 io_A_Valid_1_delay_4_57;
  reg                 io_A_Valid_1_delay_5_56;
  reg                 io_A_Valid_1_delay_6_55;
  reg                 io_A_Valid_1_delay_7_54;
  reg                 io_A_Valid_1_delay_8_53;
  reg                 io_A_Valid_1_delay_9_52;
  reg                 io_A_Valid_1_delay_10_51;
  reg                 io_A_Valid_1_delay_11_50;
  reg                 io_A_Valid_1_delay_12_49;
  reg                 io_A_Valid_1_delay_13_48;
  reg                 io_A_Valid_1_delay_14_47;
  reg                 io_A_Valid_1_delay_15_46;
  reg                 io_A_Valid_1_delay_16_45;
  reg                 io_A_Valid_1_delay_17_44;
  reg                 io_A_Valid_1_delay_18_43;
  reg                 io_A_Valid_1_delay_19_42;
  reg                 io_A_Valid_1_delay_20_41;
  reg                 io_A_Valid_1_delay_21_40;
  reg                 io_A_Valid_1_delay_22_39;
  reg                 io_A_Valid_1_delay_23_38;
  reg                 io_A_Valid_1_delay_24_37;
  reg                 io_A_Valid_1_delay_25_36;
  reg                 io_A_Valid_1_delay_26_35;
  reg                 io_A_Valid_1_delay_27_34;
  reg                 io_A_Valid_1_delay_28_33;
  reg                 io_A_Valid_1_delay_29_32;
  reg                 io_A_Valid_1_delay_30_31;
  reg                 io_A_Valid_1_delay_31_30;
  reg                 io_A_Valid_1_delay_32_29;
  reg                 io_A_Valid_1_delay_33_28;
  reg                 io_A_Valid_1_delay_34_27;
  reg                 io_A_Valid_1_delay_35_26;
  reg                 io_A_Valid_1_delay_36_25;
  reg                 io_A_Valid_1_delay_37_24;
  reg                 io_A_Valid_1_delay_38_23;
  reg                 io_A_Valid_1_delay_39_22;
  reg                 io_A_Valid_1_delay_40_21;
  reg                 io_A_Valid_1_delay_41_20;
  reg                 io_A_Valid_1_delay_42_19;
  reg                 io_A_Valid_1_delay_43_18;
  reg                 io_A_Valid_1_delay_44_17;
  reg                 io_A_Valid_1_delay_45_16;
  reg                 io_A_Valid_1_delay_46_15;
  reg                 io_A_Valid_1_delay_47_14;
  reg                 io_A_Valid_1_delay_48_13;
  reg                 io_A_Valid_1_delay_49_12;
  reg                 io_A_Valid_1_delay_50_11;
  reg                 io_A_Valid_1_delay_51_10;
  reg                 io_A_Valid_1_delay_52_9;
  reg                 io_A_Valid_1_delay_53_8;
  reg                 io_A_Valid_1_delay_54_7;
  reg                 io_A_Valid_1_delay_55_6;
  reg                 io_A_Valid_1_delay_56_5;
  reg                 io_A_Valid_1_delay_57_4;
  reg                 io_A_Valid_1_delay_58_3;
  reg                 io_A_Valid_1_delay_59_2;
  reg                 io_A_Valid_1_delay_60_1;
  reg                 io_A_Valid_1_delay_61;
  reg                 io_B_Valid_61_delay_1;
  reg                 io_A_Valid_1_delay_1_61;
  reg                 io_A_Valid_1_delay_2_60;
  reg                 io_A_Valid_1_delay_3_59;
  reg                 io_A_Valid_1_delay_4_58;
  reg                 io_A_Valid_1_delay_5_57;
  reg                 io_A_Valid_1_delay_6_56;
  reg                 io_A_Valid_1_delay_7_55;
  reg                 io_A_Valid_1_delay_8_54;
  reg                 io_A_Valid_1_delay_9_53;
  reg                 io_A_Valid_1_delay_10_52;
  reg                 io_A_Valid_1_delay_11_51;
  reg                 io_A_Valid_1_delay_12_50;
  reg                 io_A_Valid_1_delay_13_49;
  reg                 io_A_Valid_1_delay_14_48;
  reg                 io_A_Valid_1_delay_15_47;
  reg                 io_A_Valid_1_delay_16_46;
  reg                 io_A_Valid_1_delay_17_45;
  reg                 io_A_Valid_1_delay_18_44;
  reg                 io_A_Valid_1_delay_19_43;
  reg                 io_A_Valid_1_delay_20_42;
  reg                 io_A_Valid_1_delay_21_41;
  reg                 io_A_Valid_1_delay_22_40;
  reg                 io_A_Valid_1_delay_23_39;
  reg                 io_A_Valid_1_delay_24_38;
  reg                 io_A_Valid_1_delay_25_37;
  reg                 io_A_Valid_1_delay_26_36;
  reg                 io_A_Valid_1_delay_27_35;
  reg                 io_A_Valid_1_delay_28_34;
  reg                 io_A_Valid_1_delay_29_33;
  reg                 io_A_Valid_1_delay_30_32;
  reg                 io_A_Valid_1_delay_31_31;
  reg                 io_A_Valid_1_delay_32_30;
  reg                 io_A_Valid_1_delay_33_29;
  reg                 io_A_Valid_1_delay_34_28;
  reg                 io_A_Valid_1_delay_35_27;
  reg                 io_A_Valid_1_delay_36_26;
  reg                 io_A_Valid_1_delay_37_25;
  reg                 io_A_Valid_1_delay_38_24;
  reg                 io_A_Valid_1_delay_39_23;
  reg                 io_A_Valid_1_delay_40_22;
  reg                 io_A_Valid_1_delay_41_21;
  reg                 io_A_Valid_1_delay_42_20;
  reg                 io_A_Valid_1_delay_43_19;
  reg                 io_A_Valid_1_delay_44_18;
  reg                 io_A_Valid_1_delay_45_17;
  reg                 io_A_Valid_1_delay_46_16;
  reg                 io_A_Valid_1_delay_47_15;
  reg                 io_A_Valid_1_delay_48_14;
  reg                 io_A_Valid_1_delay_49_13;
  reg                 io_A_Valid_1_delay_50_12;
  reg                 io_A_Valid_1_delay_51_11;
  reg                 io_A_Valid_1_delay_52_10;
  reg                 io_A_Valid_1_delay_53_9;
  reg                 io_A_Valid_1_delay_54_8;
  reg                 io_A_Valid_1_delay_55_7;
  reg                 io_A_Valid_1_delay_56_6;
  reg                 io_A_Valid_1_delay_57_5;
  reg                 io_A_Valid_1_delay_58_4;
  reg                 io_A_Valid_1_delay_59_3;
  reg                 io_A_Valid_1_delay_60_2;
  reg                 io_A_Valid_1_delay_61_1;
  reg                 io_A_Valid_1_delay_62;
  reg                 io_B_Valid_62_delay_1;
  reg                 io_A_Valid_1_delay_1_62;
  reg                 io_A_Valid_1_delay_2_61;
  reg                 io_A_Valid_1_delay_3_60;
  reg                 io_A_Valid_1_delay_4_59;
  reg                 io_A_Valid_1_delay_5_58;
  reg                 io_A_Valid_1_delay_6_57;
  reg                 io_A_Valid_1_delay_7_56;
  reg                 io_A_Valid_1_delay_8_55;
  reg                 io_A_Valid_1_delay_9_54;
  reg                 io_A_Valid_1_delay_10_53;
  reg                 io_A_Valid_1_delay_11_52;
  reg                 io_A_Valid_1_delay_12_51;
  reg                 io_A_Valid_1_delay_13_50;
  reg                 io_A_Valid_1_delay_14_49;
  reg                 io_A_Valid_1_delay_15_48;
  reg                 io_A_Valid_1_delay_16_47;
  reg                 io_A_Valid_1_delay_17_46;
  reg                 io_A_Valid_1_delay_18_45;
  reg                 io_A_Valid_1_delay_19_44;
  reg                 io_A_Valid_1_delay_20_43;
  reg                 io_A_Valid_1_delay_21_42;
  reg                 io_A_Valid_1_delay_22_41;
  reg                 io_A_Valid_1_delay_23_40;
  reg                 io_A_Valid_1_delay_24_39;
  reg                 io_A_Valid_1_delay_25_38;
  reg                 io_A_Valid_1_delay_26_37;
  reg                 io_A_Valid_1_delay_27_36;
  reg                 io_A_Valid_1_delay_28_35;
  reg                 io_A_Valid_1_delay_29_34;
  reg                 io_A_Valid_1_delay_30_33;
  reg                 io_A_Valid_1_delay_31_32;
  reg                 io_A_Valid_1_delay_32_31;
  reg                 io_A_Valid_1_delay_33_30;
  reg                 io_A_Valid_1_delay_34_29;
  reg                 io_A_Valid_1_delay_35_28;
  reg                 io_A_Valid_1_delay_36_27;
  reg                 io_A_Valid_1_delay_37_26;
  reg                 io_A_Valid_1_delay_38_25;
  reg                 io_A_Valid_1_delay_39_24;
  reg                 io_A_Valid_1_delay_40_23;
  reg                 io_A_Valid_1_delay_41_22;
  reg                 io_A_Valid_1_delay_42_21;
  reg                 io_A_Valid_1_delay_43_20;
  reg                 io_A_Valid_1_delay_44_19;
  reg                 io_A_Valid_1_delay_45_18;
  reg                 io_A_Valid_1_delay_46_17;
  reg                 io_A_Valid_1_delay_47_16;
  reg                 io_A_Valid_1_delay_48_15;
  reg                 io_A_Valid_1_delay_49_14;
  reg                 io_A_Valid_1_delay_50_13;
  reg                 io_A_Valid_1_delay_51_12;
  reg                 io_A_Valid_1_delay_52_11;
  reg                 io_A_Valid_1_delay_53_10;
  reg                 io_A_Valid_1_delay_54_9;
  reg                 io_A_Valid_1_delay_55_8;
  reg                 io_A_Valid_1_delay_56_7;
  reg                 io_A_Valid_1_delay_57_6;
  reg                 io_A_Valid_1_delay_58_5;
  reg                 io_A_Valid_1_delay_59_4;
  reg                 io_A_Valid_1_delay_60_3;
  reg                 io_A_Valid_1_delay_61_2;
  reg                 io_A_Valid_1_delay_62_1;
  reg                 io_A_Valid_1_delay_63;
  reg                 io_B_Valid_63_delay_1;
  reg        [15:0]   io_signCount_regNextWhen_2;
  reg                 io_B_Valid_0_delay_1_1;
  reg                 io_B_Valid_0_delay_2;
  reg                 io_A_Valid_2_delay_1;
  reg                 io_B_Valid_1_delay_1_1;
  reg                 io_B_Valid_1_delay_2;
  reg                 io_A_Valid_2_delay_1_1;
  reg                 io_A_Valid_2_delay_2;
  reg                 io_B_Valid_2_delay_1_1;
  reg                 io_B_Valid_2_delay_2;
  reg                 io_A_Valid_2_delay_1_2;
  reg                 io_A_Valid_2_delay_2_1;
  reg                 io_A_Valid_2_delay_3;
  reg                 io_B_Valid_3_delay_1_1;
  reg                 io_B_Valid_3_delay_2;
  reg                 io_A_Valid_2_delay_1_3;
  reg                 io_A_Valid_2_delay_2_2;
  reg                 io_A_Valid_2_delay_3_1;
  reg                 io_A_Valid_2_delay_4;
  reg                 io_B_Valid_4_delay_1_1;
  reg                 io_B_Valid_4_delay_2;
  reg                 io_A_Valid_2_delay_1_4;
  reg                 io_A_Valid_2_delay_2_3;
  reg                 io_A_Valid_2_delay_3_2;
  reg                 io_A_Valid_2_delay_4_1;
  reg                 io_A_Valid_2_delay_5;
  reg                 io_B_Valid_5_delay_1_1;
  reg                 io_B_Valid_5_delay_2;
  reg                 io_A_Valid_2_delay_1_5;
  reg                 io_A_Valid_2_delay_2_4;
  reg                 io_A_Valid_2_delay_3_3;
  reg                 io_A_Valid_2_delay_4_2;
  reg                 io_A_Valid_2_delay_5_1;
  reg                 io_A_Valid_2_delay_6;
  reg                 io_B_Valid_6_delay_1_1;
  reg                 io_B_Valid_6_delay_2;
  reg                 io_A_Valid_2_delay_1_6;
  reg                 io_A_Valid_2_delay_2_5;
  reg                 io_A_Valid_2_delay_3_4;
  reg                 io_A_Valid_2_delay_4_3;
  reg                 io_A_Valid_2_delay_5_2;
  reg                 io_A_Valid_2_delay_6_1;
  reg                 io_A_Valid_2_delay_7;
  reg                 io_B_Valid_7_delay_1_1;
  reg                 io_B_Valid_7_delay_2;
  reg                 io_A_Valid_2_delay_1_7;
  reg                 io_A_Valid_2_delay_2_6;
  reg                 io_A_Valid_2_delay_3_5;
  reg                 io_A_Valid_2_delay_4_4;
  reg                 io_A_Valid_2_delay_5_3;
  reg                 io_A_Valid_2_delay_6_2;
  reg                 io_A_Valid_2_delay_7_1;
  reg                 io_A_Valid_2_delay_8;
  reg                 io_B_Valid_8_delay_1_1;
  reg                 io_B_Valid_8_delay_2;
  reg                 io_A_Valid_2_delay_1_8;
  reg                 io_A_Valid_2_delay_2_7;
  reg                 io_A_Valid_2_delay_3_6;
  reg                 io_A_Valid_2_delay_4_5;
  reg                 io_A_Valid_2_delay_5_4;
  reg                 io_A_Valid_2_delay_6_3;
  reg                 io_A_Valid_2_delay_7_2;
  reg                 io_A_Valid_2_delay_8_1;
  reg                 io_A_Valid_2_delay_9;
  reg                 io_B_Valid_9_delay_1_1;
  reg                 io_B_Valid_9_delay_2;
  reg                 io_A_Valid_2_delay_1_9;
  reg                 io_A_Valid_2_delay_2_8;
  reg                 io_A_Valid_2_delay_3_7;
  reg                 io_A_Valid_2_delay_4_6;
  reg                 io_A_Valid_2_delay_5_5;
  reg                 io_A_Valid_2_delay_6_4;
  reg                 io_A_Valid_2_delay_7_3;
  reg                 io_A_Valid_2_delay_8_2;
  reg                 io_A_Valid_2_delay_9_1;
  reg                 io_A_Valid_2_delay_10;
  reg                 io_B_Valid_10_delay_1_1;
  reg                 io_B_Valid_10_delay_2;
  reg                 io_A_Valid_2_delay_1_10;
  reg                 io_A_Valid_2_delay_2_9;
  reg                 io_A_Valid_2_delay_3_8;
  reg                 io_A_Valid_2_delay_4_7;
  reg                 io_A_Valid_2_delay_5_6;
  reg                 io_A_Valid_2_delay_6_5;
  reg                 io_A_Valid_2_delay_7_4;
  reg                 io_A_Valid_2_delay_8_3;
  reg                 io_A_Valid_2_delay_9_2;
  reg                 io_A_Valid_2_delay_10_1;
  reg                 io_A_Valid_2_delay_11;
  reg                 io_B_Valid_11_delay_1_1;
  reg                 io_B_Valid_11_delay_2;
  reg                 io_A_Valid_2_delay_1_11;
  reg                 io_A_Valid_2_delay_2_10;
  reg                 io_A_Valid_2_delay_3_9;
  reg                 io_A_Valid_2_delay_4_8;
  reg                 io_A_Valid_2_delay_5_7;
  reg                 io_A_Valid_2_delay_6_6;
  reg                 io_A_Valid_2_delay_7_5;
  reg                 io_A_Valid_2_delay_8_4;
  reg                 io_A_Valid_2_delay_9_3;
  reg                 io_A_Valid_2_delay_10_2;
  reg                 io_A_Valid_2_delay_11_1;
  reg                 io_A_Valid_2_delay_12;
  reg                 io_B_Valid_12_delay_1_1;
  reg                 io_B_Valid_12_delay_2;
  reg                 io_A_Valid_2_delay_1_12;
  reg                 io_A_Valid_2_delay_2_11;
  reg                 io_A_Valid_2_delay_3_10;
  reg                 io_A_Valid_2_delay_4_9;
  reg                 io_A_Valid_2_delay_5_8;
  reg                 io_A_Valid_2_delay_6_7;
  reg                 io_A_Valid_2_delay_7_6;
  reg                 io_A_Valid_2_delay_8_5;
  reg                 io_A_Valid_2_delay_9_4;
  reg                 io_A_Valid_2_delay_10_3;
  reg                 io_A_Valid_2_delay_11_2;
  reg                 io_A_Valid_2_delay_12_1;
  reg                 io_A_Valid_2_delay_13;
  reg                 io_B_Valid_13_delay_1_1;
  reg                 io_B_Valid_13_delay_2;
  reg                 io_A_Valid_2_delay_1_13;
  reg                 io_A_Valid_2_delay_2_12;
  reg                 io_A_Valid_2_delay_3_11;
  reg                 io_A_Valid_2_delay_4_10;
  reg                 io_A_Valid_2_delay_5_9;
  reg                 io_A_Valid_2_delay_6_8;
  reg                 io_A_Valid_2_delay_7_7;
  reg                 io_A_Valid_2_delay_8_6;
  reg                 io_A_Valid_2_delay_9_5;
  reg                 io_A_Valid_2_delay_10_4;
  reg                 io_A_Valid_2_delay_11_3;
  reg                 io_A_Valid_2_delay_12_2;
  reg                 io_A_Valid_2_delay_13_1;
  reg                 io_A_Valid_2_delay_14;
  reg                 io_B_Valid_14_delay_1_1;
  reg                 io_B_Valid_14_delay_2;
  reg                 io_A_Valid_2_delay_1_14;
  reg                 io_A_Valid_2_delay_2_13;
  reg                 io_A_Valid_2_delay_3_12;
  reg                 io_A_Valid_2_delay_4_11;
  reg                 io_A_Valid_2_delay_5_10;
  reg                 io_A_Valid_2_delay_6_9;
  reg                 io_A_Valid_2_delay_7_8;
  reg                 io_A_Valid_2_delay_8_7;
  reg                 io_A_Valid_2_delay_9_6;
  reg                 io_A_Valid_2_delay_10_5;
  reg                 io_A_Valid_2_delay_11_4;
  reg                 io_A_Valid_2_delay_12_3;
  reg                 io_A_Valid_2_delay_13_2;
  reg                 io_A_Valid_2_delay_14_1;
  reg                 io_A_Valid_2_delay_15;
  reg                 io_B_Valid_15_delay_1_1;
  reg                 io_B_Valid_15_delay_2;
  reg                 io_A_Valid_2_delay_1_15;
  reg                 io_A_Valid_2_delay_2_14;
  reg                 io_A_Valid_2_delay_3_13;
  reg                 io_A_Valid_2_delay_4_12;
  reg                 io_A_Valid_2_delay_5_11;
  reg                 io_A_Valid_2_delay_6_10;
  reg                 io_A_Valid_2_delay_7_9;
  reg                 io_A_Valid_2_delay_8_8;
  reg                 io_A_Valid_2_delay_9_7;
  reg                 io_A_Valid_2_delay_10_6;
  reg                 io_A_Valid_2_delay_11_5;
  reg                 io_A_Valid_2_delay_12_4;
  reg                 io_A_Valid_2_delay_13_3;
  reg                 io_A_Valid_2_delay_14_2;
  reg                 io_A_Valid_2_delay_15_1;
  reg                 io_A_Valid_2_delay_16;
  reg                 io_B_Valid_16_delay_1_1;
  reg                 io_B_Valid_16_delay_2;
  reg                 io_A_Valid_2_delay_1_16;
  reg                 io_A_Valid_2_delay_2_15;
  reg                 io_A_Valid_2_delay_3_14;
  reg                 io_A_Valid_2_delay_4_13;
  reg                 io_A_Valid_2_delay_5_12;
  reg                 io_A_Valid_2_delay_6_11;
  reg                 io_A_Valid_2_delay_7_10;
  reg                 io_A_Valid_2_delay_8_9;
  reg                 io_A_Valid_2_delay_9_8;
  reg                 io_A_Valid_2_delay_10_7;
  reg                 io_A_Valid_2_delay_11_6;
  reg                 io_A_Valid_2_delay_12_5;
  reg                 io_A_Valid_2_delay_13_4;
  reg                 io_A_Valid_2_delay_14_3;
  reg                 io_A_Valid_2_delay_15_2;
  reg                 io_A_Valid_2_delay_16_1;
  reg                 io_A_Valid_2_delay_17;
  reg                 io_B_Valid_17_delay_1_1;
  reg                 io_B_Valid_17_delay_2;
  reg                 io_A_Valid_2_delay_1_17;
  reg                 io_A_Valid_2_delay_2_16;
  reg                 io_A_Valid_2_delay_3_15;
  reg                 io_A_Valid_2_delay_4_14;
  reg                 io_A_Valid_2_delay_5_13;
  reg                 io_A_Valid_2_delay_6_12;
  reg                 io_A_Valid_2_delay_7_11;
  reg                 io_A_Valid_2_delay_8_10;
  reg                 io_A_Valid_2_delay_9_9;
  reg                 io_A_Valid_2_delay_10_8;
  reg                 io_A_Valid_2_delay_11_7;
  reg                 io_A_Valid_2_delay_12_6;
  reg                 io_A_Valid_2_delay_13_5;
  reg                 io_A_Valid_2_delay_14_4;
  reg                 io_A_Valid_2_delay_15_3;
  reg                 io_A_Valid_2_delay_16_2;
  reg                 io_A_Valid_2_delay_17_1;
  reg                 io_A_Valid_2_delay_18;
  reg                 io_B_Valid_18_delay_1_1;
  reg                 io_B_Valid_18_delay_2;
  reg                 io_A_Valid_2_delay_1_18;
  reg                 io_A_Valid_2_delay_2_17;
  reg                 io_A_Valid_2_delay_3_16;
  reg                 io_A_Valid_2_delay_4_15;
  reg                 io_A_Valid_2_delay_5_14;
  reg                 io_A_Valid_2_delay_6_13;
  reg                 io_A_Valid_2_delay_7_12;
  reg                 io_A_Valid_2_delay_8_11;
  reg                 io_A_Valid_2_delay_9_10;
  reg                 io_A_Valid_2_delay_10_9;
  reg                 io_A_Valid_2_delay_11_8;
  reg                 io_A_Valid_2_delay_12_7;
  reg                 io_A_Valid_2_delay_13_6;
  reg                 io_A_Valid_2_delay_14_5;
  reg                 io_A_Valid_2_delay_15_4;
  reg                 io_A_Valid_2_delay_16_3;
  reg                 io_A_Valid_2_delay_17_2;
  reg                 io_A_Valid_2_delay_18_1;
  reg                 io_A_Valid_2_delay_19;
  reg                 io_B_Valid_19_delay_1_1;
  reg                 io_B_Valid_19_delay_2;
  reg                 io_A_Valid_2_delay_1_19;
  reg                 io_A_Valid_2_delay_2_18;
  reg                 io_A_Valid_2_delay_3_17;
  reg                 io_A_Valid_2_delay_4_16;
  reg                 io_A_Valid_2_delay_5_15;
  reg                 io_A_Valid_2_delay_6_14;
  reg                 io_A_Valid_2_delay_7_13;
  reg                 io_A_Valid_2_delay_8_12;
  reg                 io_A_Valid_2_delay_9_11;
  reg                 io_A_Valid_2_delay_10_10;
  reg                 io_A_Valid_2_delay_11_9;
  reg                 io_A_Valid_2_delay_12_8;
  reg                 io_A_Valid_2_delay_13_7;
  reg                 io_A_Valid_2_delay_14_6;
  reg                 io_A_Valid_2_delay_15_5;
  reg                 io_A_Valid_2_delay_16_4;
  reg                 io_A_Valid_2_delay_17_3;
  reg                 io_A_Valid_2_delay_18_2;
  reg                 io_A_Valid_2_delay_19_1;
  reg                 io_A_Valid_2_delay_20;
  reg                 io_B_Valid_20_delay_1_1;
  reg                 io_B_Valid_20_delay_2;
  reg                 io_A_Valid_2_delay_1_20;
  reg                 io_A_Valid_2_delay_2_19;
  reg                 io_A_Valid_2_delay_3_18;
  reg                 io_A_Valid_2_delay_4_17;
  reg                 io_A_Valid_2_delay_5_16;
  reg                 io_A_Valid_2_delay_6_15;
  reg                 io_A_Valid_2_delay_7_14;
  reg                 io_A_Valid_2_delay_8_13;
  reg                 io_A_Valid_2_delay_9_12;
  reg                 io_A_Valid_2_delay_10_11;
  reg                 io_A_Valid_2_delay_11_10;
  reg                 io_A_Valid_2_delay_12_9;
  reg                 io_A_Valid_2_delay_13_8;
  reg                 io_A_Valid_2_delay_14_7;
  reg                 io_A_Valid_2_delay_15_6;
  reg                 io_A_Valid_2_delay_16_5;
  reg                 io_A_Valid_2_delay_17_4;
  reg                 io_A_Valid_2_delay_18_3;
  reg                 io_A_Valid_2_delay_19_2;
  reg                 io_A_Valid_2_delay_20_1;
  reg                 io_A_Valid_2_delay_21;
  reg                 io_B_Valid_21_delay_1_1;
  reg                 io_B_Valid_21_delay_2;
  reg                 io_A_Valid_2_delay_1_21;
  reg                 io_A_Valid_2_delay_2_20;
  reg                 io_A_Valid_2_delay_3_19;
  reg                 io_A_Valid_2_delay_4_18;
  reg                 io_A_Valid_2_delay_5_17;
  reg                 io_A_Valid_2_delay_6_16;
  reg                 io_A_Valid_2_delay_7_15;
  reg                 io_A_Valid_2_delay_8_14;
  reg                 io_A_Valid_2_delay_9_13;
  reg                 io_A_Valid_2_delay_10_12;
  reg                 io_A_Valid_2_delay_11_11;
  reg                 io_A_Valid_2_delay_12_10;
  reg                 io_A_Valid_2_delay_13_9;
  reg                 io_A_Valid_2_delay_14_8;
  reg                 io_A_Valid_2_delay_15_7;
  reg                 io_A_Valid_2_delay_16_6;
  reg                 io_A_Valid_2_delay_17_5;
  reg                 io_A_Valid_2_delay_18_4;
  reg                 io_A_Valid_2_delay_19_3;
  reg                 io_A_Valid_2_delay_20_2;
  reg                 io_A_Valid_2_delay_21_1;
  reg                 io_A_Valid_2_delay_22;
  reg                 io_B_Valid_22_delay_1_1;
  reg                 io_B_Valid_22_delay_2;
  reg                 io_A_Valid_2_delay_1_22;
  reg                 io_A_Valid_2_delay_2_21;
  reg                 io_A_Valid_2_delay_3_20;
  reg                 io_A_Valid_2_delay_4_19;
  reg                 io_A_Valid_2_delay_5_18;
  reg                 io_A_Valid_2_delay_6_17;
  reg                 io_A_Valid_2_delay_7_16;
  reg                 io_A_Valid_2_delay_8_15;
  reg                 io_A_Valid_2_delay_9_14;
  reg                 io_A_Valid_2_delay_10_13;
  reg                 io_A_Valid_2_delay_11_12;
  reg                 io_A_Valid_2_delay_12_11;
  reg                 io_A_Valid_2_delay_13_10;
  reg                 io_A_Valid_2_delay_14_9;
  reg                 io_A_Valid_2_delay_15_8;
  reg                 io_A_Valid_2_delay_16_7;
  reg                 io_A_Valid_2_delay_17_6;
  reg                 io_A_Valid_2_delay_18_5;
  reg                 io_A_Valid_2_delay_19_4;
  reg                 io_A_Valid_2_delay_20_3;
  reg                 io_A_Valid_2_delay_21_2;
  reg                 io_A_Valid_2_delay_22_1;
  reg                 io_A_Valid_2_delay_23;
  reg                 io_B_Valid_23_delay_1_1;
  reg                 io_B_Valid_23_delay_2;
  reg                 io_A_Valid_2_delay_1_23;
  reg                 io_A_Valid_2_delay_2_22;
  reg                 io_A_Valid_2_delay_3_21;
  reg                 io_A_Valid_2_delay_4_20;
  reg                 io_A_Valid_2_delay_5_19;
  reg                 io_A_Valid_2_delay_6_18;
  reg                 io_A_Valid_2_delay_7_17;
  reg                 io_A_Valid_2_delay_8_16;
  reg                 io_A_Valid_2_delay_9_15;
  reg                 io_A_Valid_2_delay_10_14;
  reg                 io_A_Valid_2_delay_11_13;
  reg                 io_A_Valid_2_delay_12_12;
  reg                 io_A_Valid_2_delay_13_11;
  reg                 io_A_Valid_2_delay_14_10;
  reg                 io_A_Valid_2_delay_15_9;
  reg                 io_A_Valid_2_delay_16_8;
  reg                 io_A_Valid_2_delay_17_7;
  reg                 io_A_Valid_2_delay_18_6;
  reg                 io_A_Valid_2_delay_19_5;
  reg                 io_A_Valid_2_delay_20_4;
  reg                 io_A_Valid_2_delay_21_3;
  reg                 io_A_Valid_2_delay_22_2;
  reg                 io_A_Valid_2_delay_23_1;
  reg                 io_A_Valid_2_delay_24;
  reg                 io_B_Valid_24_delay_1_1;
  reg                 io_B_Valid_24_delay_2;
  reg                 io_A_Valid_2_delay_1_24;
  reg                 io_A_Valid_2_delay_2_23;
  reg                 io_A_Valid_2_delay_3_22;
  reg                 io_A_Valid_2_delay_4_21;
  reg                 io_A_Valid_2_delay_5_20;
  reg                 io_A_Valid_2_delay_6_19;
  reg                 io_A_Valid_2_delay_7_18;
  reg                 io_A_Valid_2_delay_8_17;
  reg                 io_A_Valid_2_delay_9_16;
  reg                 io_A_Valid_2_delay_10_15;
  reg                 io_A_Valid_2_delay_11_14;
  reg                 io_A_Valid_2_delay_12_13;
  reg                 io_A_Valid_2_delay_13_12;
  reg                 io_A_Valid_2_delay_14_11;
  reg                 io_A_Valid_2_delay_15_10;
  reg                 io_A_Valid_2_delay_16_9;
  reg                 io_A_Valid_2_delay_17_8;
  reg                 io_A_Valid_2_delay_18_7;
  reg                 io_A_Valid_2_delay_19_6;
  reg                 io_A_Valid_2_delay_20_5;
  reg                 io_A_Valid_2_delay_21_4;
  reg                 io_A_Valid_2_delay_22_3;
  reg                 io_A_Valid_2_delay_23_2;
  reg                 io_A_Valid_2_delay_24_1;
  reg                 io_A_Valid_2_delay_25;
  reg                 io_B_Valid_25_delay_1_1;
  reg                 io_B_Valid_25_delay_2;
  reg                 io_A_Valid_2_delay_1_25;
  reg                 io_A_Valid_2_delay_2_24;
  reg                 io_A_Valid_2_delay_3_23;
  reg                 io_A_Valid_2_delay_4_22;
  reg                 io_A_Valid_2_delay_5_21;
  reg                 io_A_Valid_2_delay_6_20;
  reg                 io_A_Valid_2_delay_7_19;
  reg                 io_A_Valid_2_delay_8_18;
  reg                 io_A_Valid_2_delay_9_17;
  reg                 io_A_Valid_2_delay_10_16;
  reg                 io_A_Valid_2_delay_11_15;
  reg                 io_A_Valid_2_delay_12_14;
  reg                 io_A_Valid_2_delay_13_13;
  reg                 io_A_Valid_2_delay_14_12;
  reg                 io_A_Valid_2_delay_15_11;
  reg                 io_A_Valid_2_delay_16_10;
  reg                 io_A_Valid_2_delay_17_9;
  reg                 io_A_Valid_2_delay_18_8;
  reg                 io_A_Valid_2_delay_19_7;
  reg                 io_A_Valid_2_delay_20_6;
  reg                 io_A_Valid_2_delay_21_5;
  reg                 io_A_Valid_2_delay_22_4;
  reg                 io_A_Valid_2_delay_23_3;
  reg                 io_A_Valid_2_delay_24_2;
  reg                 io_A_Valid_2_delay_25_1;
  reg                 io_A_Valid_2_delay_26;
  reg                 io_B_Valid_26_delay_1_1;
  reg                 io_B_Valid_26_delay_2;
  reg                 io_A_Valid_2_delay_1_26;
  reg                 io_A_Valid_2_delay_2_25;
  reg                 io_A_Valid_2_delay_3_24;
  reg                 io_A_Valid_2_delay_4_23;
  reg                 io_A_Valid_2_delay_5_22;
  reg                 io_A_Valid_2_delay_6_21;
  reg                 io_A_Valid_2_delay_7_20;
  reg                 io_A_Valid_2_delay_8_19;
  reg                 io_A_Valid_2_delay_9_18;
  reg                 io_A_Valid_2_delay_10_17;
  reg                 io_A_Valid_2_delay_11_16;
  reg                 io_A_Valid_2_delay_12_15;
  reg                 io_A_Valid_2_delay_13_14;
  reg                 io_A_Valid_2_delay_14_13;
  reg                 io_A_Valid_2_delay_15_12;
  reg                 io_A_Valid_2_delay_16_11;
  reg                 io_A_Valid_2_delay_17_10;
  reg                 io_A_Valid_2_delay_18_9;
  reg                 io_A_Valid_2_delay_19_8;
  reg                 io_A_Valid_2_delay_20_7;
  reg                 io_A_Valid_2_delay_21_6;
  reg                 io_A_Valid_2_delay_22_5;
  reg                 io_A_Valid_2_delay_23_4;
  reg                 io_A_Valid_2_delay_24_3;
  reg                 io_A_Valid_2_delay_25_2;
  reg                 io_A_Valid_2_delay_26_1;
  reg                 io_A_Valid_2_delay_27;
  reg                 io_B_Valid_27_delay_1_1;
  reg                 io_B_Valid_27_delay_2;
  reg                 io_A_Valid_2_delay_1_27;
  reg                 io_A_Valid_2_delay_2_26;
  reg                 io_A_Valid_2_delay_3_25;
  reg                 io_A_Valid_2_delay_4_24;
  reg                 io_A_Valid_2_delay_5_23;
  reg                 io_A_Valid_2_delay_6_22;
  reg                 io_A_Valid_2_delay_7_21;
  reg                 io_A_Valid_2_delay_8_20;
  reg                 io_A_Valid_2_delay_9_19;
  reg                 io_A_Valid_2_delay_10_18;
  reg                 io_A_Valid_2_delay_11_17;
  reg                 io_A_Valid_2_delay_12_16;
  reg                 io_A_Valid_2_delay_13_15;
  reg                 io_A_Valid_2_delay_14_14;
  reg                 io_A_Valid_2_delay_15_13;
  reg                 io_A_Valid_2_delay_16_12;
  reg                 io_A_Valid_2_delay_17_11;
  reg                 io_A_Valid_2_delay_18_10;
  reg                 io_A_Valid_2_delay_19_9;
  reg                 io_A_Valid_2_delay_20_8;
  reg                 io_A_Valid_2_delay_21_7;
  reg                 io_A_Valid_2_delay_22_6;
  reg                 io_A_Valid_2_delay_23_5;
  reg                 io_A_Valid_2_delay_24_4;
  reg                 io_A_Valid_2_delay_25_3;
  reg                 io_A_Valid_2_delay_26_2;
  reg                 io_A_Valid_2_delay_27_1;
  reg                 io_A_Valid_2_delay_28;
  reg                 io_B_Valid_28_delay_1_1;
  reg                 io_B_Valid_28_delay_2;
  reg                 io_A_Valid_2_delay_1_28;
  reg                 io_A_Valid_2_delay_2_27;
  reg                 io_A_Valid_2_delay_3_26;
  reg                 io_A_Valid_2_delay_4_25;
  reg                 io_A_Valid_2_delay_5_24;
  reg                 io_A_Valid_2_delay_6_23;
  reg                 io_A_Valid_2_delay_7_22;
  reg                 io_A_Valid_2_delay_8_21;
  reg                 io_A_Valid_2_delay_9_20;
  reg                 io_A_Valid_2_delay_10_19;
  reg                 io_A_Valid_2_delay_11_18;
  reg                 io_A_Valid_2_delay_12_17;
  reg                 io_A_Valid_2_delay_13_16;
  reg                 io_A_Valid_2_delay_14_15;
  reg                 io_A_Valid_2_delay_15_14;
  reg                 io_A_Valid_2_delay_16_13;
  reg                 io_A_Valid_2_delay_17_12;
  reg                 io_A_Valid_2_delay_18_11;
  reg                 io_A_Valid_2_delay_19_10;
  reg                 io_A_Valid_2_delay_20_9;
  reg                 io_A_Valid_2_delay_21_8;
  reg                 io_A_Valid_2_delay_22_7;
  reg                 io_A_Valid_2_delay_23_6;
  reg                 io_A_Valid_2_delay_24_5;
  reg                 io_A_Valid_2_delay_25_4;
  reg                 io_A_Valid_2_delay_26_3;
  reg                 io_A_Valid_2_delay_27_2;
  reg                 io_A_Valid_2_delay_28_1;
  reg                 io_A_Valid_2_delay_29;
  reg                 io_B_Valid_29_delay_1_1;
  reg                 io_B_Valid_29_delay_2;
  reg                 io_A_Valid_2_delay_1_29;
  reg                 io_A_Valid_2_delay_2_28;
  reg                 io_A_Valid_2_delay_3_27;
  reg                 io_A_Valid_2_delay_4_26;
  reg                 io_A_Valid_2_delay_5_25;
  reg                 io_A_Valid_2_delay_6_24;
  reg                 io_A_Valid_2_delay_7_23;
  reg                 io_A_Valid_2_delay_8_22;
  reg                 io_A_Valid_2_delay_9_21;
  reg                 io_A_Valid_2_delay_10_20;
  reg                 io_A_Valid_2_delay_11_19;
  reg                 io_A_Valid_2_delay_12_18;
  reg                 io_A_Valid_2_delay_13_17;
  reg                 io_A_Valid_2_delay_14_16;
  reg                 io_A_Valid_2_delay_15_15;
  reg                 io_A_Valid_2_delay_16_14;
  reg                 io_A_Valid_2_delay_17_13;
  reg                 io_A_Valid_2_delay_18_12;
  reg                 io_A_Valid_2_delay_19_11;
  reg                 io_A_Valid_2_delay_20_10;
  reg                 io_A_Valid_2_delay_21_9;
  reg                 io_A_Valid_2_delay_22_8;
  reg                 io_A_Valid_2_delay_23_7;
  reg                 io_A_Valid_2_delay_24_6;
  reg                 io_A_Valid_2_delay_25_5;
  reg                 io_A_Valid_2_delay_26_4;
  reg                 io_A_Valid_2_delay_27_3;
  reg                 io_A_Valid_2_delay_28_2;
  reg                 io_A_Valid_2_delay_29_1;
  reg                 io_A_Valid_2_delay_30;
  reg                 io_B_Valid_30_delay_1_1;
  reg                 io_B_Valid_30_delay_2;
  reg                 io_A_Valid_2_delay_1_30;
  reg                 io_A_Valid_2_delay_2_29;
  reg                 io_A_Valid_2_delay_3_28;
  reg                 io_A_Valid_2_delay_4_27;
  reg                 io_A_Valid_2_delay_5_26;
  reg                 io_A_Valid_2_delay_6_25;
  reg                 io_A_Valid_2_delay_7_24;
  reg                 io_A_Valid_2_delay_8_23;
  reg                 io_A_Valid_2_delay_9_22;
  reg                 io_A_Valid_2_delay_10_21;
  reg                 io_A_Valid_2_delay_11_20;
  reg                 io_A_Valid_2_delay_12_19;
  reg                 io_A_Valid_2_delay_13_18;
  reg                 io_A_Valid_2_delay_14_17;
  reg                 io_A_Valid_2_delay_15_16;
  reg                 io_A_Valid_2_delay_16_15;
  reg                 io_A_Valid_2_delay_17_14;
  reg                 io_A_Valid_2_delay_18_13;
  reg                 io_A_Valid_2_delay_19_12;
  reg                 io_A_Valid_2_delay_20_11;
  reg                 io_A_Valid_2_delay_21_10;
  reg                 io_A_Valid_2_delay_22_9;
  reg                 io_A_Valid_2_delay_23_8;
  reg                 io_A_Valid_2_delay_24_7;
  reg                 io_A_Valid_2_delay_25_6;
  reg                 io_A_Valid_2_delay_26_5;
  reg                 io_A_Valid_2_delay_27_4;
  reg                 io_A_Valid_2_delay_28_3;
  reg                 io_A_Valid_2_delay_29_2;
  reg                 io_A_Valid_2_delay_30_1;
  reg                 io_A_Valid_2_delay_31;
  reg                 io_B_Valid_31_delay_1_1;
  reg                 io_B_Valid_31_delay_2;
  reg                 io_A_Valid_2_delay_1_31;
  reg                 io_A_Valid_2_delay_2_30;
  reg                 io_A_Valid_2_delay_3_29;
  reg                 io_A_Valid_2_delay_4_28;
  reg                 io_A_Valid_2_delay_5_27;
  reg                 io_A_Valid_2_delay_6_26;
  reg                 io_A_Valid_2_delay_7_25;
  reg                 io_A_Valid_2_delay_8_24;
  reg                 io_A_Valid_2_delay_9_23;
  reg                 io_A_Valid_2_delay_10_22;
  reg                 io_A_Valid_2_delay_11_21;
  reg                 io_A_Valid_2_delay_12_20;
  reg                 io_A_Valid_2_delay_13_19;
  reg                 io_A_Valid_2_delay_14_18;
  reg                 io_A_Valid_2_delay_15_17;
  reg                 io_A_Valid_2_delay_16_16;
  reg                 io_A_Valid_2_delay_17_15;
  reg                 io_A_Valid_2_delay_18_14;
  reg                 io_A_Valid_2_delay_19_13;
  reg                 io_A_Valid_2_delay_20_12;
  reg                 io_A_Valid_2_delay_21_11;
  reg                 io_A_Valid_2_delay_22_10;
  reg                 io_A_Valid_2_delay_23_9;
  reg                 io_A_Valid_2_delay_24_8;
  reg                 io_A_Valid_2_delay_25_7;
  reg                 io_A_Valid_2_delay_26_6;
  reg                 io_A_Valid_2_delay_27_5;
  reg                 io_A_Valid_2_delay_28_4;
  reg                 io_A_Valid_2_delay_29_3;
  reg                 io_A_Valid_2_delay_30_2;
  reg                 io_A_Valid_2_delay_31_1;
  reg                 io_A_Valid_2_delay_32;
  reg                 io_B_Valid_32_delay_1_1;
  reg                 io_B_Valid_32_delay_2;
  reg                 io_A_Valid_2_delay_1_32;
  reg                 io_A_Valid_2_delay_2_31;
  reg                 io_A_Valid_2_delay_3_30;
  reg                 io_A_Valid_2_delay_4_29;
  reg                 io_A_Valid_2_delay_5_28;
  reg                 io_A_Valid_2_delay_6_27;
  reg                 io_A_Valid_2_delay_7_26;
  reg                 io_A_Valid_2_delay_8_25;
  reg                 io_A_Valid_2_delay_9_24;
  reg                 io_A_Valid_2_delay_10_23;
  reg                 io_A_Valid_2_delay_11_22;
  reg                 io_A_Valid_2_delay_12_21;
  reg                 io_A_Valid_2_delay_13_20;
  reg                 io_A_Valid_2_delay_14_19;
  reg                 io_A_Valid_2_delay_15_18;
  reg                 io_A_Valid_2_delay_16_17;
  reg                 io_A_Valid_2_delay_17_16;
  reg                 io_A_Valid_2_delay_18_15;
  reg                 io_A_Valid_2_delay_19_14;
  reg                 io_A_Valid_2_delay_20_13;
  reg                 io_A_Valid_2_delay_21_12;
  reg                 io_A_Valid_2_delay_22_11;
  reg                 io_A_Valid_2_delay_23_10;
  reg                 io_A_Valid_2_delay_24_9;
  reg                 io_A_Valid_2_delay_25_8;
  reg                 io_A_Valid_2_delay_26_7;
  reg                 io_A_Valid_2_delay_27_6;
  reg                 io_A_Valid_2_delay_28_5;
  reg                 io_A_Valid_2_delay_29_4;
  reg                 io_A_Valid_2_delay_30_3;
  reg                 io_A_Valid_2_delay_31_2;
  reg                 io_A_Valid_2_delay_32_1;
  reg                 io_A_Valid_2_delay_33;
  reg                 io_B_Valid_33_delay_1_1;
  reg                 io_B_Valid_33_delay_2;
  reg                 io_A_Valid_2_delay_1_33;
  reg                 io_A_Valid_2_delay_2_32;
  reg                 io_A_Valid_2_delay_3_31;
  reg                 io_A_Valid_2_delay_4_30;
  reg                 io_A_Valid_2_delay_5_29;
  reg                 io_A_Valid_2_delay_6_28;
  reg                 io_A_Valid_2_delay_7_27;
  reg                 io_A_Valid_2_delay_8_26;
  reg                 io_A_Valid_2_delay_9_25;
  reg                 io_A_Valid_2_delay_10_24;
  reg                 io_A_Valid_2_delay_11_23;
  reg                 io_A_Valid_2_delay_12_22;
  reg                 io_A_Valid_2_delay_13_21;
  reg                 io_A_Valid_2_delay_14_20;
  reg                 io_A_Valid_2_delay_15_19;
  reg                 io_A_Valid_2_delay_16_18;
  reg                 io_A_Valid_2_delay_17_17;
  reg                 io_A_Valid_2_delay_18_16;
  reg                 io_A_Valid_2_delay_19_15;
  reg                 io_A_Valid_2_delay_20_14;
  reg                 io_A_Valid_2_delay_21_13;
  reg                 io_A_Valid_2_delay_22_12;
  reg                 io_A_Valid_2_delay_23_11;
  reg                 io_A_Valid_2_delay_24_10;
  reg                 io_A_Valid_2_delay_25_9;
  reg                 io_A_Valid_2_delay_26_8;
  reg                 io_A_Valid_2_delay_27_7;
  reg                 io_A_Valid_2_delay_28_6;
  reg                 io_A_Valid_2_delay_29_5;
  reg                 io_A_Valid_2_delay_30_4;
  reg                 io_A_Valid_2_delay_31_3;
  reg                 io_A_Valid_2_delay_32_2;
  reg                 io_A_Valid_2_delay_33_1;
  reg                 io_A_Valid_2_delay_34;
  reg                 io_B_Valid_34_delay_1_1;
  reg                 io_B_Valid_34_delay_2;
  reg                 io_A_Valid_2_delay_1_34;
  reg                 io_A_Valid_2_delay_2_33;
  reg                 io_A_Valid_2_delay_3_32;
  reg                 io_A_Valid_2_delay_4_31;
  reg                 io_A_Valid_2_delay_5_30;
  reg                 io_A_Valid_2_delay_6_29;
  reg                 io_A_Valid_2_delay_7_28;
  reg                 io_A_Valid_2_delay_8_27;
  reg                 io_A_Valid_2_delay_9_26;
  reg                 io_A_Valid_2_delay_10_25;
  reg                 io_A_Valid_2_delay_11_24;
  reg                 io_A_Valid_2_delay_12_23;
  reg                 io_A_Valid_2_delay_13_22;
  reg                 io_A_Valid_2_delay_14_21;
  reg                 io_A_Valid_2_delay_15_20;
  reg                 io_A_Valid_2_delay_16_19;
  reg                 io_A_Valid_2_delay_17_18;
  reg                 io_A_Valid_2_delay_18_17;
  reg                 io_A_Valid_2_delay_19_16;
  reg                 io_A_Valid_2_delay_20_15;
  reg                 io_A_Valid_2_delay_21_14;
  reg                 io_A_Valid_2_delay_22_13;
  reg                 io_A_Valid_2_delay_23_12;
  reg                 io_A_Valid_2_delay_24_11;
  reg                 io_A_Valid_2_delay_25_10;
  reg                 io_A_Valid_2_delay_26_9;
  reg                 io_A_Valid_2_delay_27_8;
  reg                 io_A_Valid_2_delay_28_7;
  reg                 io_A_Valid_2_delay_29_6;
  reg                 io_A_Valid_2_delay_30_5;
  reg                 io_A_Valid_2_delay_31_4;
  reg                 io_A_Valid_2_delay_32_3;
  reg                 io_A_Valid_2_delay_33_2;
  reg                 io_A_Valid_2_delay_34_1;
  reg                 io_A_Valid_2_delay_35;
  reg                 io_B_Valid_35_delay_1_1;
  reg                 io_B_Valid_35_delay_2;
  reg                 io_A_Valid_2_delay_1_35;
  reg                 io_A_Valid_2_delay_2_34;
  reg                 io_A_Valid_2_delay_3_33;
  reg                 io_A_Valid_2_delay_4_32;
  reg                 io_A_Valid_2_delay_5_31;
  reg                 io_A_Valid_2_delay_6_30;
  reg                 io_A_Valid_2_delay_7_29;
  reg                 io_A_Valid_2_delay_8_28;
  reg                 io_A_Valid_2_delay_9_27;
  reg                 io_A_Valid_2_delay_10_26;
  reg                 io_A_Valid_2_delay_11_25;
  reg                 io_A_Valid_2_delay_12_24;
  reg                 io_A_Valid_2_delay_13_23;
  reg                 io_A_Valid_2_delay_14_22;
  reg                 io_A_Valid_2_delay_15_21;
  reg                 io_A_Valid_2_delay_16_20;
  reg                 io_A_Valid_2_delay_17_19;
  reg                 io_A_Valid_2_delay_18_18;
  reg                 io_A_Valid_2_delay_19_17;
  reg                 io_A_Valid_2_delay_20_16;
  reg                 io_A_Valid_2_delay_21_15;
  reg                 io_A_Valid_2_delay_22_14;
  reg                 io_A_Valid_2_delay_23_13;
  reg                 io_A_Valid_2_delay_24_12;
  reg                 io_A_Valid_2_delay_25_11;
  reg                 io_A_Valid_2_delay_26_10;
  reg                 io_A_Valid_2_delay_27_9;
  reg                 io_A_Valid_2_delay_28_8;
  reg                 io_A_Valid_2_delay_29_7;
  reg                 io_A_Valid_2_delay_30_6;
  reg                 io_A_Valid_2_delay_31_5;
  reg                 io_A_Valid_2_delay_32_4;
  reg                 io_A_Valid_2_delay_33_3;
  reg                 io_A_Valid_2_delay_34_2;
  reg                 io_A_Valid_2_delay_35_1;
  reg                 io_A_Valid_2_delay_36;
  reg                 io_B_Valid_36_delay_1_1;
  reg                 io_B_Valid_36_delay_2;
  reg                 io_A_Valid_2_delay_1_36;
  reg                 io_A_Valid_2_delay_2_35;
  reg                 io_A_Valid_2_delay_3_34;
  reg                 io_A_Valid_2_delay_4_33;
  reg                 io_A_Valid_2_delay_5_32;
  reg                 io_A_Valid_2_delay_6_31;
  reg                 io_A_Valid_2_delay_7_30;
  reg                 io_A_Valid_2_delay_8_29;
  reg                 io_A_Valid_2_delay_9_28;
  reg                 io_A_Valid_2_delay_10_27;
  reg                 io_A_Valid_2_delay_11_26;
  reg                 io_A_Valid_2_delay_12_25;
  reg                 io_A_Valid_2_delay_13_24;
  reg                 io_A_Valid_2_delay_14_23;
  reg                 io_A_Valid_2_delay_15_22;
  reg                 io_A_Valid_2_delay_16_21;
  reg                 io_A_Valid_2_delay_17_20;
  reg                 io_A_Valid_2_delay_18_19;
  reg                 io_A_Valid_2_delay_19_18;
  reg                 io_A_Valid_2_delay_20_17;
  reg                 io_A_Valid_2_delay_21_16;
  reg                 io_A_Valid_2_delay_22_15;
  reg                 io_A_Valid_2_delay_23_14;
  reg                 io_A_Valid_2_delay_24_13;
  reg                 io_A_Valid_2_delay_25_12;
  reg                 io_A_Valid_2_delay_26_11;
  reg                 io_A_Valid_2_delay_27_10;
  reg                 io_A_Valid_2_delay_28_9;
  reg                 io_A_Valid_2_delay_29_8;
  reg                 io_A_Valid_2_delay_30_7;
  reg                 io_A_Valid_2_delay_31_6;
  reg                 io_A_Valid_2_delay_32_5;
  reg                 io_A_Valid_2_delay_33_4;
  reg                 io_A_Valid_2_delay_34_3;
  reg                 io_A_Valid_2_delay_35_2;
  reg                 io_A_Valid_2_delay_36_1;
  reg                 io_A_Valid_2_delay_37;
  reg                 io_B_Valid_37_delay_1_1;
  reg                 io_B_Valid_37_delay_2;
  reg                 io_A_Valid_2_delay_1_37;
  reg                 io_A_Valid_2_delay_2_36;
  reg                 io_A_Valid_2_delay_3_35;
  reg                 io_A_Valid_2_delay_4_34;
  reg                 io_A_Valid_2_delay_5_33;
  reg                 io_A_Valid_2_delay_6_32;
  reg                 io_A_Valid_2_delay_7_31;
  reg                 io_A_Valid_2_delay_8_30;
  reg                 io_A_Valid_2_delay_9_29;
  reg                 io_A_Valid_2_delay_10_28;
  reg                 io_A_Valid_2_delay_11_27;
  reg                 io_A_Valid_2_delay_12_26;
  reg                 io_A_Valid_2_delay_13_25;
  reg                 io_A_Valid_2_delay_14_24;
  reg                 io_A_Valid_2_delay_15_23;
  reg                 io_A_Valid_2_delay_16_22;
  reg                 io_A_Valid_2_delay_17_21;
  reg                 io_A_Valid_2_delay_18_20;
  reg                 io_A_Valid_2_delay_19_19;
  reg                 io_A_Valid_2_delay_20_18;
  reg                 io_A_Valid_2_delay_21_17;
  reg                 io_A_Valid_2_delay_22_16;
  reg                 io_A_Valid_2_delay_23_15;
  reg                 io_A_Valid_2_delay_24_14;
  reg                 io_A_Valid_2_delay_25_13;
  reg                 io_A_Valid_2_delay_26_12;
  reg                 io_A_Valid_2_delay_27_11;
  reg                 io_A_Valid_2_delay_28_10;
  reg                 io_A_Valid_2_delay_29_9;
  reg                 io_A_Valid_2_delay_30_8;
  reg                 io_A_Valid_2_delay_31_7;
  reg                 io_A_Valid_2_delay_32_6;
  reg                 io_A_Valid_2_delay_33_5;
  reg                 io_A_Valid_2_delay_34_4;
  reg                 io_A_Valid_2_delay_35_3;
  reg                 io_A_Valid_2_delay_36_2;
  reg                 io_A_Valid_2_delay_37_1;
  reg                 io_A_Valid_2_delay_38;
  reg                 io_B_Valid_38_delay_1_1;
  reg                 io_B_Valid_38_delay_2;
  reg                 io_A_Valid_2_delay_1_38;
  reg                 io_A_Valid_2_delay_2_37;
  reg                 io_A_Valid_2_delay_3_36;
  reg                 io_A_Valid_2_delay_4_35;
  reg                 io_A_Valid_2_delay_5_34;
  reg                 io_A_Valid_2_delay_6_33;
  reg                 io_A_Valid_2_delay_7_32;
  reg                 io_A_Valid_2_delay_8_31;
  reg                 io_A_Valid_2_delay_9_30;
  reg                 io_A_Valid_2_delay_10_29;
  reg                 io_A_Valid_2_delay_11_28;
  reg                 io_A_Valid_2_delay_12_27;
  reg                 io_A_Valid_2_delay_13_26;
  reg                 io_A_Valid_2_delay_14_25;
  reg                 io_A_Valid_2_delay_15_24;
  reg                 io_A_Valid_2_delay_16_23;
  reg                 io_A_Valid_2_delay_17_22;
  reg                 io_A_Valid_2_delay_18_21;
  reg                 io_A_Valid_2_delay_19_20;
  reg                 io_A_Valid_2_delay_20_19;
  reg                 io_A_Valid_2_delay_21_18;
  reg                 io_A_Valid_2_delay_22_17;
  reg                 io_A_Valid_2_delay_23_16;
  reg                 io_A_Valid_2_delay_24_15;
  reg                 io_A_Valid_2_delay_25_14;
  reg                 io_A_Valid_2_delay_26_13;
  reg                 io_A_Valid_2_delay_27_12;
  reg                 io_A_Valid_2_delay_28_11;
  reg                 io_A_Valid_2_delay_29_10;
  reg                 io_A_Valid_2_delay_30_9;
  reg                 io_A_Valid_2_delay_31_8;
  reg                 io_A_Valid_2_delay_32_7;
  reg                 io_A_Valid_2_delay_33_6;
  reg                 io_A_Valid_2_delay_34_5;
  reg                 io_A_Valid_2_delay_35_4;
  reg                 io_A_Valid_2_delay_36_3;
  reg                 io_A_Valid_2_delay_37_2;
  reg                 io_A_Valid_2_delay_38_1;
  reg                 io_A_Valid_2_delay_39;
  reg                 io_B_Valid_39_delay_1_1;
  reg                 io_B_Valid_39_delay_2;
  reg                 io_A_Valid_2_delay_1_39;
  reg                 io_A_Valid_2_delay_2_38;
  reg                 io_A_Valid_2_delay_3_37;
  reg                 io_A_Valid_2_delay_4_36;
  reg                 io_A_Valid_2_delay_5_35;
  reg                 io_A_Valid_2_delay_6_34;
  reg                 io_A_Valid_2_delay_7_33;
  reg                 io_A_Valid_2_delay_8_32;
  reg                 io_A_Valid_2_delay_9_31;
  reg                 io_A_Valid_2_delay_10_30;
  reg                 io_A_Valid_2_delay_11_29;
  reg                 io_A_Valid_2_delay_12_28;
  reg                 io_A_Valid_2_delay_13_27;
  reg                 io_A_Valid_2_delay_14_26;
  reg                 io_A_Valid_2_delay_15_25;
  reg                 io_A_Valid_2_delay_16_24;
  reg                 io_A_Valid_2_delay_17_23;
  reg                 io_A_Valid_2_delay_18_22;
  reg                 io_A_Valid_2_delay_19_21;
  reg                 io_A_Valid_2_delay_20_20;
  reg                 io_A_Valid_2_delay_21_19;
  reg                 io_A_Valid_2_delay_22_18;
  reg                 io_A_Valid_2_delay_23_17;
  reg                 io_A_Valid_2_delay_24_16;
  reg                 io_A_Valid_2_delay_25_15;
  reg                 io_A_Valid_2_delay_26_14;
  reg                 io_A_Valid_2_delay_27_13;
  reg                 io_A_Valid_2_delay_28_12;
  reg                 io_A_Valid_2_delay_29_11;
  reg                 io_A_Valid_2_delay_30_10;
  reg                 io_A_Valid_2_delay_31_9;
  reg                 io_A_Valid_2_delay_32_8;
  reg                 io_A_Valid_2_delay_33_7;
  reg                 io_A_Valid_2_delay_34_6;
  reg                 io_A_Valid_2_delay_35_5;
  reg                 io_A_Valid_2_delay_36_4;
  reg                 io_A_Valid_2_delay_37_3;
  reg                 io_A_Valid_2_delay_38_2;
  reg                 io_A_Valid_2_delay_39_1;
  reg                 io_A_Valid_2_delay_40;
  reg                 io_B_Valid_40_delay_1_1;
  reg                 io_B_Valid_40_delay_2;
  reg                 io_A_Valid_2_delay_1_40;
  reg                 io_A_Valid_2_delay_2_39;
  reg                 io_A_Valid_2_delay_3_38;
  reg                 io_A_Valid_2_delay_4_37;
  reg                 io_A_Valid_2_delay_5_36;
  reg                 io_A_Valid_2_delay_6_35;
  reg                 io_A_Valid_2_delay_7_34;
  reg                 io_A_Valid_2_delay_8_33;
  reg                 io_A_Valid_2_delay_9_32;
  reg                 io_A_Valid_2_delay_10_31;
  reg                 io_A_Valid_2_delay_11_30;
  reg                 io_A_Valid_2_delay_12_29;
  reg                 io_A_Valid_2_delay_13_28;
  reg                 io_A_Valid_2_delay_14_27;
  reg                 io_A_Valid_2_delay_15_26;
  reg                 io_A_Valid_2_delay_16_25;
  reg                 io_A_Valid_2_delay_17_24;
  reg                 io_A_Valid_2_delay_18_23;
  reg                 io_A_Valid_2_delay_19_22;
  reg                 io_A_Valid_2_delay_20_21;
  reg                 io_A_Valid_2_delay_21_20;
  reg                 io_A_Valid_2_delay_22_19;
  reg                 io_A_Valid_2_delay_23_18;
  reg                 io_A_Valid_2_delay_24_17;
  reg                 io_A_Valid_2_delay_25_16;
  reg                 io_A_Valid_2_delay_26_15;
  reg                 io_A_Valid_2_delay_27_14;
  reg                 io_A_Valid_2_delay_28_13;
  reg                 io_A_Valid_2_delay_29_12;
  reg                 io_A_Valid_2_delay_30_11;
  reg                 io_A_Valid_2_delay_31_10;
  reg                 io_A_Valid_2_delay_32_9;
  reg                 io_A_Valid_2_delay_33_8;
  reg                 io_A_Valid_2_delay_34_7;
  reg                 io_A_Valid_2_delay_35_6;
  reg                 io_A_Valid_2_delay_36_5;
  reg                 io_A_Valid_2_delay_37_4;
  reg                 io_A_Valid_2_delay_38_3;
  reg                 io_A_Valid_2_delay_39_2;
  reg                 io_A_Valid_2_delay_40_1;
  reg                 io_A_Valid_2_delay_41;
  reg                 io_B_Valid_41_delay_1_1;
  reg                 io_B_Valid_41_delay_2;
  reg                 io_A_Valid_2_delay_1_41;
  reg                 io_A_Valid_2_delay_2_40;
  reg                 io_A_Valid_2_delay_3_39;
  reg                 io_A_Valid_2_delay_4_38;
  reg                 io_A_Valid_2_delay_5_37;
  reg                 io_A_Valid_2_delay_6_36;
  reg                 io_A_Valid_2_delay_7_35;
  reg                 io_A_Valid_2_delay_8_34;
  reg                 io_A_Valid_2_delay_9_33;
  reg                 io_A_Valid_2_delay_10_32;
  reg                 io_A_Valid_2_delay_11_31;
  reg                 io_A_Valid_2_delay_12_30;
  reg                 io_A_Valid_2_delay_13_29;
  reg                 io_A_Valid_2_delay_14_28;
  reg                 io_A_Valid_2_delay_15_27;
  reg                 io_A_Valid_2_delay_16_26;
  reg                 io_A_Valid_2_delay_17_25;
  reg                 io_A_Valid_2_delay_18_24;
  reg                 io_A_Valid_2_delay_19_23;
  reg                 io_A_Valid_2_delay_20_22;
  reg                 io_A_Valid_2_delay_21_21;
  reg                 io_A_Valid_2_delay_22_20;
  reg                 io_A_Valid_2_delay_23_19;
  reg                 io_A_Valid_2_delay_24_18;
  reg                 io_A_Valid_2_delay_25_17;
  reg                 io_A_Valid_2_delay_26_16;
  reg                 io_A_Valid_2_delay_27_15;
  reg                 io_A_Valid_2_delay_28_14;
  reg                 io_A_Valid_2_delay_29_13;
  reg                 io_A_Valid_2_delay_30_12;
  reg                 io_A_Valid_2_delay_31_11;
  reg                 io_A_Valid_2_delay_32_10;
  reg                 io_A_Valid_2_delay_33_9;
  reg                 io_A_Valid_2_delay_34_8;
  reg                 io_A_Valid_2_delay_35_7;
  reg                 io_A_Valid_2_delay_36_6;
  reg                 io_A_Valid_2_delay_37_5;
  reg                 io_A_Valid_2_delay_38_4;
  reg                 io_A_Valid_2_delay_39_3;
  reg                 io_A_Valid_2_delay_40_2;
  reg                 io_A_Valid_2_delay_41_1;
  reg                 io_A_Valid_2_delay_42;
  reg                 io_B_Valid_42_delay_1_1;
  reg                 io_B_Valid_42_delay_2;
  reg                 io_A_Valid_2_delay_1_42;
  reg                 io_A_Valid_2_delay_2_41;
  reg                 io_A_Valid_2_delay_3_40;
  reg                 io_A_Valid_2_delay_4_39;
  reg                 io_A_Valid_2_delay_5_38;
  reg                 io_A_Valid_2_delay_6_37;
  reg                 io_A_Valid_2_delay_7_36;
  reg                 io_A_Valid_2_delay_8_35;
  reg                 io_A_Valid_2_delay_9_34;
  reg                 io_A_Valid_2_delay_10_33;
  reg                 io_A_Valid_2_delay_11_32;
  reg                 io_A_Valid_2_delay_12_31;
  reg                 io_A_Valid_2_delay_13_30;
  reg                 io_A_Valid_2_delay_14_29;
  reg                 io_A_Valid_2_delay_15_28;
  reg                 io_A_Valid_2_delay_16_27;
  reg                 io_A_Valid_2_delay_17_26;
  reg                 io_A_Valid_2_delay_18_25;
  reg                 io_A_Valid_2_delay_19_24;
  reg                 io_A_Valid_2_delay_20_23;
  reg                 io_A_Valid_2_delay_21_22;
  reg                 io_A_Valid_2_delay_22_21;
  reg                 io_A_Valid_2_delay_23_20;
  reg                 io_A_Valid_2_delay_24_19;
  reg                 io_A_Valid_2_delay_25_18;
  reg                 io_A_Valid_2_delay_26_17;
  reg                 io_A_Valid_2_delay_27_16;
  reg                 io_A_Valid_2_delay_28_15;
  reg                 io_A_Valid_2_delay_29_14;
  reg                 io_A_Valid_2_delay_30_13;
  reg                 io_A_Valid_2_delay_31_12;
  reg                 io_A_Valid_2_delay_32_11;
  reg                 io_A_Valid_2_delay_33_10;
  reg                 io_A_Valid_2_delay_34_9;
  reg                 io_A_Valid_2_delay_35_8;
  reg                 io_A_Valid_2_delay_36_7;
  reg                 io_A_Valid_2_delay_37_6;
  reg                 io_A_Valid_2_delay_38_5;
  reg                 io_A_Valid_2_delay_39_4;
  reg                 io_A_Valid_2_delay_40_3;
  reg                 io_A_Valid_2_delay_41_2;
  reg                 io_A_Valid_2_delay_42_1;
  reg                 io_A_Valid_2_delay_43;
  reg                 io_B_Valid_43_delay_1_1;
  reg                 io_B_Valid_43_delay_2;
  reg                 io_A_Valid_2_delay_1_43;
  reg                 io_A_Valid_2_delay_2_42;
  reg                 io_A_Valid_2_delay_3_41;
  reg                 io_A_Valid_2_delay_4_40;
  reg                 io_A_Valid_2_delay_5_39;
  reg                 io_A_Valid_2_delay_6_38;
  reg                 io_A_Valid_2_delay_7_37;
  reg                 io_A_Valid_2_delay_8_36;
  reg                 io_A_Valid_2_delay_9_35;
  reg                 io_A_Valid_2_delay_10_34;
  reg                 io_A_Valid_2_delay_11_33;
  reg                 io_A_Valid_2_delay_12_32;
  reg                 io_A_Valid_2_delay_13_31;
  reg                 io_A_Valid_2_delay_14_30;
  reg                 io_A_Valid_2_delay_15_29;
  reg                 io_A_Valid_2_delay_16_28;
  reg                 io_A_Valid_2_delay_17_27;
  reg                 io_A_Valid_2_delay_18_26;
  reg                 io_A_Valid_2_delay_19_25;
  reg                 io_A_Valid_2_delay_20_24;
  reg                 io_A_Valid_2_delay_21_23;
  reg                 io_A_Valid_2_delay_22_22;
  reg                 io_A_Valid_2_delay_23_21;
  reg                 io_A_Valid_2_delay_24_20;
  reg                 io_A_Valid_2_delay_25_19;
  reg                 io_A_Valid_2_delay_26_18;
  reg                 io_A_Valid_2_delay_27_17;
  reg                 io_A_Valid_2_delay_28_16;
  reg                 io_A_Valid_2_delay_29_15;
  reg                 io_A_Valid_2_delay_30_14;
  reg                 io_A_Valid_2_delay_31_13;
  reg                 io_A_Valid_2_delay_32_12;
  reg                 io_A_Valid_2_delay_33_11;
  reg                 io_A_Valid_2_delay_34_10;
  reg                 io_A_Valid_2_delay_35_9;
  reg                 io_A_Valid_2_delay_36_8;
  reg                 io_A_Valid_2_delay_37_7;
  reg                 io_A_Valid_2_delay_38_6;
  reg                 io_A_Valid_2_delay_39_5;
  reg                 io_A_Valid_2_delay_40_4;
  reg                 io_A_Valid_2_delay_41_3;
  reg                 io_A_Valid_2_delay_42_2;
  reg                 io_A_Valid_2_delay_43_1;
  reg                 io_A_Valid_2_delay_44;
  reg                 io_B_Valid_44_delay_1_1;
  reg                 io_B_Valid_44_delay_2;
  reg                 io_A_Valid_2_delay_1_44;
  reg                 io_A_Valid_2_delay_2_43;
  reg                 io_A_Valid_2_delay_3_42;
  reg                 io_A_Valid_2_delay_4_41;
  reg                 io_A_Valid_2_delay_5_40;
  reg                 io_A_Valid_2_delay_6_39;
  reg                 io_A_Valid_2_delay_7_38;
  reg                 io_A_Valid_2_delay_8_37;
  reg                 io_A_Valid_2_delay_9_36;
  reg                 io_A_Valid_2_delay_10_35;
  reg                 io_A_Valid_2_delay_11_34;
  reg                 io_A_Valid_2_delay_12_33;
  reg                 io_A_Valid_2_delay_13_32;
  reg                 io_A_Valid_2_delay_14_31;
  reg                 io_A_Valid_2_delay_15_30;
  reg                 io_A_Valid_2_delay_16_29;
  reg                 io_A_Valid_2_delay_17_28;
  reg                 io_A_Valid_2_delay_18_27;
  reg                 io_A_Valid_2_delay_19_26;
  reg                 io_A_Valid_2_delay_20_25;
  reg                 io_A_Valid_2_delay_21_24;
  reg                 io_A_Valid_2_delay_22_23;
  reg                 io_A_Valid_2_delay_23_22;
  reg                 io_A_Valid_2_delay_24_21;
  reg                 io_A_Valid_2_delay_25_20;
  reg                 io_A_Valid_2_delay_26_19;
  reg                 io_A_Valid_2_delay_27_18;
  reg                 io_A_Valid_2_delay_28_17;
  reg                 io_A_Valid_2_delay_29_16;
  reg                 io_A_Valid_2_delay_30_15;
  reg                 io_A_Valid_2_delay_31_14;
  reg                 io_A_Valid_2_delay_32_13;
  reg                 io_A_Valid_2_delay_33_12;
  reg                 io_A_Valid_2_delay_34_11;
  reg                 io_A_Valid_2_delay_35_10;
  reg                 io_A_Valid_2_delay_36_9;
  reg                 io_A_Valid_2_delay_37_8;
  reg                 io_A_Valid_2_delay_38_7;
  reg                 io_A_Valid_2_delay_39_6;
  reg                 io_A_Valid_2_delay_40_5;
  reg                 io_A_Valid_2_delay_41_4;
  reg                 io_A_Valid_2_delay_42_3;
  reg                 io_A_Valid_2_delay_43_2;
  reg                 io_A_Valid_2_delay_44_1;
  reg                 io_A_Valid_2_delay_45;
  reg                 io_B_Valid_45_delay_1_1;
  reg                 io_B_Valid_45_delay_2;
  reg                 io_A_Valid_2_delay_1_45;
  reg                 io_A_Valid_2_delay_2_44;
  reg                 io_A_Valid_2_delay_3_43;
  reg                 io_A_Valid_2_delay_4_42;
  reg                 io_A_Valid_2_delay_5_41;
  reg                 io_A_Valid_2_delay_6_40;
  reg                 io_A_Valid_2_delay_7_39;
  reg                 io_A_Valid_2_delay_8_38;
  reg                 io_A_Valid_2_delay_9_37;
  reg                 io_A_Valid_2_delay_10_36;
  reg                 io_A_Valid_2_delay_11_35;
  reg                 io_A_Valid_2_delay_12_34;
  reg                 io_A_Valid_2_delay_13_33;
  reg                 io_A_Valid_2_delay_14_32;
  reg                 io_A_Valid_2_delay_15_31;
  reg                 io_A_Valid_2_delay_16_30;
  reg                 io_A_Valid_2_delay_17_29;
  reg                 io_A_Valid_2_delay_18_28;
  reg                 io_A_Valid_2_delay_19_27;
  reg                 io_A_Valid_2_delay_20_26;
  reg                 io_A_Valid_2_delay_21_25;
  reg                 io_A_Valid_2_delay_22_24;
  reg                 io_A_Valid_2_delay_23_23;
  reg                 io_A_Valid_2_delay_24_22;
  reg                 io_A_Valid_2_delay_25_21;
  reg                 io_A_Valid_2_delay_26_20;
  reg                 io_A_Valid_2_delay_27_19;
  reg                 io_A_Valid_2_delay_28_18;
  reg                 io_A_Valid_2_delay_29_17;
  reg                 io_A_Valid_2_delay_30_16;
  reg                 io_A_Valid_2_delay_31_15;
  reg                 io_A_Valid_2_delay_32_14;
  reg                 io_A_Valid_2_delay_33_13;
  reg                 io_A_Valid_2_delay_34_12;
  reg                 io_A_Valid_2_delay_35_11;
  reg                 io_A_Valid_2_delay_36_10;
  reg                 io_A_Valid_2_delay_37_9;
  reg                 io_A_Valid_2_delay_38_8;
  reg                 io_A_Valid_2_delay_39_7;
  reg                 io_A_Valid_2_delay_40_6;
  reg                 io_A_Valid_2_delay_41_5;
  reg                 io_A_Valid_2_delay_42_4;
  reg                 io_A_Valid_2_delay_43_3;
  reg                 io_A_Valid_2_delay_44_2;
  reg                 io_A_Valid_2_delay_45_1;
  reg                 io_A_Valid_2_delay_46;
  reg                 io_B_Valid_46_delay_1_1;
  reg                 io_B_Valid_46_delay_2;
  reg                 io_A_Valid_2_delay_1_46;
  reg                 io_A_Valid_2_delay_2_45;
  reg                 io_A_Valid_2_delay_3_44;
  reg                 io_A_Valid_2_delay_4_43;
  reg                 io_A_Valid_2_delay_5_42;
  reg                 io_A_Valid_2_delay_6_41;
  reg                 io_A_Valid_2_delay_7_40;
  reg                 io_A_Valid_2_delay_8_39;
  reg                 io_A_Valid_2_delay_9_38;
  reg                 io_A_Valid_2_delay_10_37;
  reg                 io_A_Valid_2_delay_11_36;
  reg                 io_A_Valid_2_delay_12_35;
  reg                 io_A_Valid_2_delay_13_34;
  reg                 io_A_Valid_2_delay_14_33;
  reg                 io_A_Valid_2_delay_15_32;
  reg                 io_A_Valid_2_delay_16_31;
  reg                 io_A_Valid_2_delay_17_30;
  reg                 io_A_Valid_2_delay_18_29;
  reg                 io_A_Valid_2_delay_19_28;
  reg                 io_A_Valid_2_delay_20_27;
  reg                 io_A_Valid_2_delay_21_26;
  reg                 io_A_Valid_2_delay_22_25;
  reg                 io_A_Valid_2_delay_23_24;
  reg                 io_A_Valid_2_delay_24_23;
  reg                 io_A_Valid_2_delay_25_22;
  reg                 io_A_Valid_2_delay_26_21;
  reg                 io_A_Valid_2_delay_27_20;
  reg                 io_A_Valid_2_delay_28_19;
  reg                 io_A_Valid_2_delay_29_18;
  reg                 io_A_Valid_2_delay_30_17;
  reg                 io_A_Valid_2_delay_31_16;
  reg                 io_A_Valid_2_delay_32_15;
  reg                 io_A_Valid_2_delay_33_14;
  reg                 io_A_Valid_2_delay_34_13;
  reg                 io_A_Valid_2_delay_35_12;
  reg                 io_A_Valid_2_delay_36_11;
  reg                 io_A_Valid_2_delay_37_10;
  reg                 io_A_Valid_2_delay_38_9;
  reg                 io_A_Valid_2_delay_39_8;
  reg                 io_A_Valid_2_delay_40_7;
  reg                 io_A_Valid_2_delay_41_6;
  reg                 io_A_Valid_2_delay_42_5;
  reg                 io_A_Valid_2_delay_43_4;
  reg                 io_A_Valid_2_delay_44_3;
  reg                 io_A_Valid_2_delay_45_2;
  reg                 io_A_Valid_2_delay_46_1;
  reg                 io_A_Valid_2_delay_47;
  reg                 io_B_Valid_47_delay_1_1;
  reg                 io_B_Valid_47_delay_2;
  reg                 io_A_Valid_2_delay_1_47;
  reg                 io_A_Valid_2_delay_2_46;
  reg                 io_A_Valid_2_delay_3_45;
  reg                 io_A_Valid_2_delay_4_44;
  reg                 io_A_Valid_2_delay_5_43;
  reg                 io_A_Valid_2_delay_6_42;
  reg                 io_A_Valid_2_delay_7_41;
  reg                 io_A_Valid_2_delay_8_40;
  reg                 io_A_Valid_2_delay_9_39;
  reg                 io_A_Valid_2_delay_10_38;
  reg                 io_A_Valid_2_delay_11_37;
  reg                 io_A_Valid_2_delay_12_36;
  reg                 io_A_Valid_2_delay_13_35;
  reg                 io_A_Valid_2_delay_14_34;
  reg                 io_A_Valid_2_delay_15_33;
  reg                 io_A_Valid_2_delay_16_32;
  reg                 io_A_Valid_2_delay_17_31;
  reg                 io_A_Valid_2_delay_18_30;
  reg                 io_A_Valid_2_delay_19_29;
  reg                 io_A_Valid_2_delay_20_28;
  reg                 io_A_Valid_2_delay_21_27;
  reg                 io_A_Valid_2_delay_22_26;
  reg                 io_A_Valid_2_delay_23_25;
  reg                 io_A_Valid_2_delay_24_24;
  reg                 io_A_Valid_2_delay_25_23;
  reg                 io_A_Valid_2_delay_26_22;
  reg                 io_A_Valid_2_delay_27_21;
  reg                 io_A_Valid_2_delay_28_20;
  reg                 io_A_Valid_2_delay_29_19;
  reg                 io_A_Valid_2_delay_30_18;
  reg                 io_A_Valid_2_delay_31_17;
  reg                 io_A_Valid_2_delay_32_16;
  reg                 io_A_Valid_2_delay_33_15;
  reg                 io_A_Valid_2_delay_34_14;
  reg                 io_A_Valid_2_delay_35_13;
  reg                 io_A_Valid_2_delay_36_12;
  reg                 io_A_Valid_2_delay_37_11;
  reg                 io_A_Valid_2_delay_38_10;
  reg                 io_A_Valid_2_delay_39_9;
  reg                 io_A_Valid_2_delay_40_8;
  reg                 io_A_Valid_2_delay_41_7;
  reg                 io_A_Valid_2_delay_42_6;
  reg                 io_A_Valid_2_delay_43_5;
  reg                 io_A_Valid_2_delay_44_4;
  reg                 io_A_Valid_2_delay_45_3;
  reg                 io_A_Valid_2_delay_46_2;
  reg                 io_A_Valid_2_delay_47_1;
  reg                 io_A_Valid_2_delay_48;
  reg                 io_B_Valid_48_delay_1_1;
  reg                 io_B_Valid_48_delay_2;
  reg                 io_A_Valid_2_delay_1_48;
  reg                 io_A_Valid_2_delay_2_47;
  reg                 io_A_Valid_2_delay_3_46;
  reg                 io_A_Valid_2_delay_4_45;
  reg                 io_A_Valid_2_delay_5_44;
  reg                 io_A_Valid_2_delay_6_43;
  reg                 io_A_Valid_2_delay_7_42;
  reg                 io_A_Valid_2_delay_8_41;
  reg                 io_A_Valid_2_delay_9_40;
  reg                 io_A_Valid_2_delay_10_39;
  reg                 io_A_Valid_2_delay_11_38;
  reg                 io_A_Valid_2_delay_12_37;
  reg                 io_A_Valid_2_delay_13_36;
  reg                 io_A_Valid_2_delay_14_35;
  reg                 io_A_Valid_2_delay_15_34;
  reg                 io_A_Valid_2_delay_16_33;
  reg                 io_A_Valid_2_delay_17_32;
  reg                 io_A_Valid_2_delay_18_31;
  reg                 io_A_Valid_2_delay_19_30;
  reg                 io_A_Valid_2_delay_20_29;
  reg                 io_A_Valid_2_delay_21_28;
  reg                 io_A_Valid_2_delay_22_27;
  reg                 io_A_Valid_2_delay_23_26;
  reg                 io_A_Valid_2_delay_24_25;
  reg                 io_A_Valid_2_delay_25_24;
  reg                 io_A_Valid_2_delay_26_23;
  reg                 io_A_Valid_2_delay_27_22;
  reg                 io_A_Valid_2_delay_28_21;
  reg                 io_A_Valid_2_delay_29_20;
  reg                 io_A_Valid_2_delay_30_19;
  reg                 io_A_Valid_2_delay_31_18;
  reg                 io_A_Valid_2_delay_32_17;
  reg                 io_A_Valid_2_delay_33_16;
  reg                 io_A_Valid_2_delay_34_15;
  reg                 io_A_Valid_2_delay_35_14;
  reg                 io_A_Valid_2_delay_36_13;
  reg                 io_A_Valid_2_delay_37_12;
  reg                 io_A_Valid_2_delay_38_11;
  reg                 io_A_Valid_2_delay_39_10;
  reg                 io_A_Valid_2_delay_40_9;
  reg                 io_A_Valid_2_delay_41_8;
  reg                 io_A_Valid_2_delay_42_7;
  reg                 io_A_Valid_2_delay_43_6;
  reg                 io_A_Valid_2_delay_44_5;
  reg                 io_A_Valid_2_delay_45_4;
  reg                 io_A_Valid_2_delay_46_3;
  reg                 io_A_Valid_2_delay_47_2;
  reg                 io_A_Valid_2_delay_48_1;
  reg                 io_A_Valid_2_delay_49;
  reg                 io_B_Valid_49_delay_1_1;
  reg                 io_B_Valid_49_delay_2;
  reg                 io_A_Valid_2_delay_1_49;
  reg                 io_A_Valid_2_delay_2_48;
  reg                 io_A_Valid_2_delay_3_47;
  reg                 io_A_Valid_2_delay_4_46;
  reg                 io_A_Valid_2_delay_5_45;
  reg                 io_A_Valid_2_delay_6_44;
  reg                 io_A_Valid_2_delay_7_43;
  reg                 io_A_Valid_2_delay_8_42;
  reg                 io_A_Valid_2_delay_9_41;
  reg                 io_A_Valid_2_delay_10_40;
  reg                 io_A_Valid_2_delay_11_39;
  reg                 io_A_Valid_2_delay_12_38;
  reg                 io_A_Valid_2_delay_13_37;
  reg                 io_A_Valid_2_delay_14_36;
  reg                 io_A_Valid_2_delay_15_35;
  reg                 io_A_Valid_2_delay_16_34;
  reg                 io_A_Valid_2_delay_17_33;
  reg                 io_A_Valid_2_delay_18_32;
  reg                 io_A_Valid_2_delay_19_31;
  reg                 io_A_Valid_2_delay_20_30;
  reg                 io_A_Valid_2_delay_21_29;
  reg                 io_A_Valid_2_delay_22_28;
  reg                 io_A_Valid_2_delay_23_27;
  reg                 io_A_Valid_2_delay_24_26;
  reg                 io_A_Valid_2_delay_25_25;
  reg                 io_A_Valid_2_delay_26_24;
  reg                 io_A_Valid_2_delay_27_23;
  reg                 io_A_Valid_2_delay_28_22;
  reg                 io_A_Valid_2_delay_29_21;
  reg                 io_A_Valid_2_delay_30_20;
  reg                 io_A_Valid_2_delay_31_19;
  reg                 io_A_Valid_2_delay_32_18;
  reg                 io_A_Valid_2_delay_33_17;
  reg                 io_A_Valid_2_delay_34_16;
  reg                 io_A_Valid_2_delay_35_15;
  reg                 io_A_Valid_2_delay_36_14;
  reg                 io_A_Valid_2_delay_37_13;
  reg                 io_A_Valid_2_delay_38_12;
  reg                 io_A_Valid_2_delay_39_11;
  reg                 io_A_Valid_2_delay_40_10;
  reg                 io_A_Valid_2_delay_41_9;
  reg                 io_A_Valid_2_delay_42_8;
  reg                 io_A_Valid_2_delay_43_7;
  reg                 io_A_Valid_2_delay_44_6;
  reg                 io_A_Valid_2_delay_45_5;
  reg                 io_A_Valid_2_delay_46_4;
  reg                 io_A_Valid_2_delay_47_3;
  reg                 io_A_Valid_2_delay_48_2;
  reg                 io_A_Valid_2_delay_49_1;
  reg                 io_A_Valid_2_delay_50;
  reg                 io_B_Valid_50_delay_1_1;
  reg                 io_B_Valid_50_delay_2;
  reg                 io_A_Valid_2_delay_1_50;
  reg                 io_A_Valid_2_delay_2_49;
  reg                 io_A_Valid_2_delay_3_48;
  reg                 io_A_Valid_2_delay_4_47;
  reg                 io_A_Valid_2_delay_5_46;
  reg                 io_A_Valid_2_delay_6_45;
  reg                 io_A_Valid_2_delay_7_44;
  reg                 io_A_Valid_2_delay_8_43;
  reg                 io_A_Valid_2_delay_9_42;
  reg                 io_A_Valid_2_delay_10_41;
  reg                 io_A_Valid_2_delay_11_40;
  reg                 io_A_Valid_2_delay_12_39;
  reg                 io_A_Valid_2_delay_13_38;
  reg                 io_A_Valid_2_delay_14_37;
  reg                 io_A_Valid_2_delay_15_36;
  reg                 io_A_Valid_2_delay_16_35;
  reg                 io_A_Valid_2_delay_17_34;
  reg                 io_A_Valid_2_delay_18_33;
  reg                 io_A_Valid_2_delay_19_32;
  reg                 io_A_Valid_2_delay_20_31;
  reg                 io_A_Valid_2_delay_21_30;
  reg                 io_A_Valid_2_delay_22_29;
  reg                 io_A_Valid_2_delay_23_28;
  reg                 io_A_Valid_2_delay_24_27;
  reg                 io_A_Valid_2_delay_25_26;
  reg                 io_A_Valid_2_delay_26_25;
  reg                 io_A_Valid_2_delay_27_24;
  reg                 io_A_Valid_2_delay_28_23;
  reg                 io_A_Valid_2_delay_29_22;
  reg                 io_A_Valid_2_delay_30_21;
  reg                 io_A_Valid_2_delay_31_20;
  reg                 io_A_Valid_2_delay_32_19;
  reg                 io_A_Valid_2_delay_33_18;
  reg                 io_A_Valid_2_delay_34_17;
  reg                 io_A_Valid_2_delay_35_16;
  reg                 io_A_Valid_2_delay_36_15;
  reg                 io_A_Valid_2_delay_37_14;
  reg                 io_A_Valid_2_delay_38_13;
  reg                 io_A_Valid_2_delay_39_12;
  reg                 io_A_Valid_2_delay_40_11;
  reg                 io_A_Valid_2_delay_41_10;
  reg                 io_A_Valid_2_delay_42_9;
  reg                 io_A_Valid_2_delay_43_8;
  reg                 io_A_Valid_2_delay_44_7;
  reg                 io_A_Valid_2_delay_45_6;
  reg                 io_A_Valid_2_delay_46_5;
  reg                 io_A_Valid_2_delay_47_4;
  reg                 io_A_Valid_2_delay_48_3;
  reg                 io_A_Valid_2_delay_49_2;
  reg                 io_A_Valid_2_delay_50_1;
  reg                 io_A_Valid_2_delay_51;
  reg                 io_B_Valid_51_delay_1_1;
  reg                 io_B_Valid_51_delay_2;
  reg                 io_A_Valid_2_delay_1_51;
  reg                 io_A_Valid_2_delay_2_50;
  reg                 io_A_Valid_2_delay_3_49;
  reg                 io_A_Valid_2_delay_4_48;
  reg                 io_A_Valid_2_delay_5_47;
  reg                 io_A_Valid_2_delay_6_46;
  reg                 io_A_Valid_2_delay_7_45;
  reg                 io_A_Valid_2_delay_8_44;
  reg                 io_A_Valid_2_delay_9_43;
  reg                 io_A_Valid_2_delay_10_42;
  reg                 io_A_Valid_2_delay_11_41;
  reg                 io_A_Valid_2_delay_12_40;
  reg                 io_A_Valid_2_delay_13_39;
  reg                 io_A_Valid_2_delay_14_38;
  reg                 io_A_Valid_2_delay_15_37;
  reg                 io_A_Valid_2_delay_16_36;
  reg                 io_A_Valid_2_delay_17_35;
  reg                 io_A_Valid_2_delay_18_34;
  reg                 io_A_Valid_2_delay_19_33;
  reg                 io_A_Valid_2_delay_20_32;
  reg                 io_A_Valid_2_delay_21_31;
  reg                 io_A_Valid_2_delay_22_30;
  reg                 io_A_Valid_2_delay_23_29;
  reg                 io_A_Valid_2_delay_24_28;
  reg                 io_A_Valid_2_delay_25_27;
  reg                 io_A_Valid_2_delay_26_26;
  reg                 io_A_Valid_2_delay_27_25;
  reg                 io_A_Valid_2_delay_28_24;
  reg                 io_A_Valid_2_delay_29_23;
  reg                 io_A_Valid_2_delay_30_22;
  reg                 io_A_Valid_2_delay_31_21;
  reg                 io_A_Valid_2_delay_32_20;
  reg                 io_A_Valid_2_delay_33_19;
  reg                 io_A_Valid_2_delay_34_18;
  reg                 io_A_Valid_2_delay_35_17;
  reg                 io_A_Valid_2_delay_36_16;
  reg                 io_A_Valid_2_delay_37_15;
  reg                 io_A_Valid_2_delay_38_14;
  reg                 io_A_Valid_2_delay_39_13;
  reg                 io_A_Valid_2_delay_40_12;
  reg                 io_A_Valid_2_delay_41_11;
  reg                 io_A_Valid_2_delay_42_10;
  reg                 io_A_Valid_2_delay_43_9;
  reg                 io_A_Valid_2_delay_44_8;
  reg                 io_A_Valid_2_delay_45_7;
  reg                 io_A_Valid_2_delay_46_6;
  reg                 io_A_Valid_2_delay_47_5;
  reg                 io_A_Valid_2_delay_48_4;
  reg                 io_A_Valid_2_delay_49_3;
  reg                 io_A_Valid_2_delay_50_2;
  reg                 io_A_Valid_2_delay_51_1;
  reg                 io_A_Valid_2_delay_52;
  reg                 io_B_Valid_52_delay_1_1;
  reg                 io_B_Valid_52_delay_2;
  reg                 io_A_Valid_2_delay_1_52;
  reg                 io_A_Valid_2_delay_2_51;
  reg                 io_A_Valid_2_delay_3_50;
  reg                 io_A_Valid_2_delay_4_49;
  reg                 io_A_Valid_2_delay_5_48;
  reg                 io_A_Valid_2_delay_6_47;
  reg                 io_A_Valid_2_delay_7_46;
  reg                 io_A_Valid_2_delay_8_45;
  reg                 io_A_Valid_2_delay_9_44;
  reg                 io_A_Valid_2_delay_10_43;
  reg                 io_A_Valid_2_delay_11_42;
  reg                 io_A_Valid_2_delay_12_41;
  reg                 io_A_Valid_2_delay_13_40;
  reg                 io_A_Valid_2_delay_14_39;
  reg                 io_A_Valid_2_delay_15_38;
  reg                 io_A_Valid_2_delay_16_37;
  reg                 io_A_Valid_2_delay_17_36;
  reg                 io_A_Valid_2_delay_18_35;
  reg                 io_A_Valid_2_delay_19_34;
  reg                 io_A_Valid_2_delay_20_33;
  reg                 io_A_Valid_2_delay_21_32;
  reg                 io_A_Valid_2_delay_22_31;
  reg                 io_A_Valid_2_delay_23_30;
  reg                 io_A_Valid_2_delay_24_29;
  reg                 io_A_Valid_2_delay_25_28;
  reg                 io_A_Valid_2_delay_26_27;
  reg                 io_A_Valid_2_delay_27_26;
  reg                 io_A_Valid_2_delay_28_25;
  reg                 io_A_Valid_2_delay_29_24;
  reg                 io_A_Valid_2_delay_30_23;
  reg                 io_A_Valid_2_delay_31_22;
  reg                 io_A_Valid_2_delay_32_21;
  reg                 io_A_Valid_2_delay_33_20;
  reg                 io_A_Valid_2_delay_34_19;
  reg                 io_A_Valid_2_delay_35_18;
  reg                 io_A_Valid_2_delay_36_17;
  reg                 io_A_Valid_2_delay_37_16;
  reg                 io_A_Valid_2_delay_38_15;
  reg                 io_A_Valid_2_delay_39_14;
  reg                 io_A_Valid_2_delay_40_13;
  reg                 io_A_Valid_2_delay_41_12;
  reg                 io_A_Valid_2_delay_42_11;
  reg                 io_A_Valid_2_delay_43_10;
  reg                 io_A_Valid_2_delay_44_9;
  reg                 io_A_Valid_2_delay_45_8;
  reg                 io_A_Valid_2_delay_46_7;
  reg                 io_A_Valid_2_delay_47_6;
  reg                 io_A_Valid_2_delay_48_5;
  reg                 io_A_Valid_2_delay_49_4;
  reg                 io_A_Valid_2_delay_50_3;
  reg                 io_A_Valid_2_delay_51_2;
  reg                 io_A_Valid_2_delay_52_1;
  reg                 io_A_Valid_2_delay_53;
  reg                 io_B_Valid_53_delay_1_1;
  reg                 io_B_Valid_53_delay_2;
  reg                 io_A_Valid_2_delay_1_53;
  reg                 io_A_Valid_2_delay_2_52;
  reg                 io_A_Valid_2_delay_3_51;
  reg                 io_A_Valid_2_delay_4_50;
  reg                 io_A_Valid_2_delay_5_49;
  reg                 io_A_Valid_2_delay_6_48;
  reg                 io_A_Valid_2_delay_7_47;
  reg                 io_A_Valid_2_delay_8_46;
  reg                 io_A_Valid_2_delay_9_45;
  reg                 io_A_Valid_2_delay_10_44;
  reg                 io_A_Valid_2_delay_11_43;
  reg                 io_A_Valid_2_delay_12_42;
  reg                 io_A_Valid_2_delay_13_41;
  reg                 io_A_Valid_2_delay_14_40;
  reg                 io_A_Valid_2_delay_15_39;
  reg                 io_A_Valid_2_delay_16_38;
  reg                 io_A_Valid_2_delay_17_37;
  reg                 io_A_Valid_2_delay_18_36;
  reg                 io_A_Valid_2_delay_19_35;
  reg                 io_A_Valid_2_delay_20_34;
  reg                 io_A_Valid_2_delay_21_33;
  reg                 io_A_Valid_2_delay_22_32;
  reg                 io_A_Valid_2_delay_23_31;
  reg                 io_A_Valid_2_delay_24_30;
  reg                 io_A_Valid_2_delay_25_29;
  reg                 io_A_Valid_2_delay_26_28;
  reg                 io_A_Valid_2_delay_27_27;
  reg                 io_A_Valid_2_delay_28_26;
  reg                 io_A_Valid_2_delay_29_25;
  reg                 io_A_Valid_2_delay_30_24;
  reg                 io_A_Valid_2_delay_31_23;
  reg                 io_A_Valid_2_delay_32_22;
  reg                 io_A_Valid_2_delay_33_21;
  reg                 io_A_Valid_2_delay_34_20;
  reg                 io_A_Valid_2_delay_35_19;
  reg                 io_A_Valid_2_delay_36_18;
  reg                 io_A_Valid_2_delay_37_17;
  reg                 io_A_Valid_2_delay_38_16;
  reg                 io_A_Valid_2_delay_39_15;
  reg                 io_A_Valid_2_delay_40_14;
  reg                 io_A_Valid_2_delay_41_13;
  reg                 io_A_Valid_2_delay_42_12;
  reg                 io_A_Valid_2_delay_43_11;
  reg                 io_A_Valid_2_delay_44_10;
  reg                 io_A_Valid_2_delay_45_9;
  reg                 io_A_Valid_2_delay_46_8;
  reg                 io_A_Valid_2_delay_47_7;
  reg                 io_A_Valid_2_delay_48_6;
  reg                 io_A_Valid_2_delay_49_5;
  reg                 io_A_Valid_2_delay_50_4;
  reg                 io_A_Valid_2_delay_51_3;
  reg                 io_A_Valid_2_delay_52_2;
  reg                 io_A_Valid_2_delay_53_1;
  reg                 io_A_Valid_2_delay_54;
  reg                 io_B_Valid_54_delay_1_1;
  reg                 io_B_Valid_54_delay_2;
  reg                 io_A_Valid_2_delay_1_54;
  reg                 io_A_Valid_2_delay_2_53;
  reg                 io_A_Valid_2_delay_3_52;
  reg                 io_A_Valid_2_delay_4_51;
  reg                 io_A_Valid_2_delay_5_50;
  reg                 io_A_Valid_2_delay_6_49;
  reg                 io_A_Valid_2_delay_7_48;
  reg                 io_A_Valid_2_delay_8_47;
  reg                 io_A_Valid_2_delay_9_46;
  reg                 io_A_Valid_2_delay_10_45;
  reg                 io_A_Valid_2_delay_11_44;
  reg                 io_A_Valid_2_delay_12_43;
  reg                 io_A_Valid_2_delay_13_42;
  reg                 io_A_Valid_2_delay_14_41;
  reg                 io_A_Valid_2_delay_15_40;
  reg                 io_A_Valid_2_delay_16_39;
  reg                 io_A_Valid_2_delay_17_38;
  reg                 io_A_Valid_2_delay_18_37;
  reg                 io_A_Valid_2_delay_19_36;
  reg                 io_A_Valid_2_delay_20_35;
  reg                 io_A_Valid_2_delay_21_34;
  reg                 io_A_Valid_2_delay_22_33;
  reg                 io_A_Valid_2_delay_23_32;
  reg                 io_A_Valid_2_delay_24_31;
  reg                 io_A_Valid_2_delay_25_30;
  reg                 io_A_Valid_2_delay_26_29;
  reg                 io_A_Valid_2_delay_27_28;
  reg                 io_A_Valid_2_delay_28_27;
  reg                 io_A_Valid_2_delay_29_26;
  reg                 io_A_Valid_2_delay_30_25;
  reg                 io_A_Valid_2_delay_31_24;
  reg                 io_A_Valid_2_delay_32_23;
  reg                 io_A_Valid_2_delay_33_22;
  reg                 io_A_Valid_2_delay_34_21;
  reg                 io_A_Valid_2_delay_35_20;
  reg                 io_A_Valid_2_delay_36_19;
  reg                 io_A_Valid_2_delay_37_18;
  reg                 io_A_Valid_2_delay_38_17;
  reg                 io_A_Valid_2_delay_39_16;
  reg                 io_A_Valid_2_delay_40_15;
  reg                 io_A_Valid_2_delay_41_14;
  reg                 io_A_Valid_2_delay_42_13;
  reg                 io_A_Valid_2_delay_43_12;
  reg                 io_A_Valid_2_delay_44_11;
  reg                 io_A_Valid_2_delay_45_10;
  reg                 io_A_Valid_2_delay_46_9;
  reg                 io_A_Valid_2_delay_47_8;
  reg                 io_A_Valid_2_delay_48_7;
  reg                 io_A_Valid_2_delay_49_6;
  reg                 io_A_Valid_2_delay_50_5;
  reg                 io_A_Valid_2_delay_51_4;
  reg                 io_A_Valid_2_delay_52_3;
  reg                 io_A_Valid_2_delay_53_2;
  reg                 io_A_Valid_2_delay_54_1;
  reg                 io_A_Valid_2_delay_55;
  reg                 io_B_Valid_55_delay_1_1;
  reg                 io_B_Valid_55_delay_2;
  reg                 io_A_Valid_2_delay_1_55;
  reg                 io_A_Valid_2_delay_2_54;
  reg                 io_A_Valid_2_delay_3_53;
  reg                 io_A_Valid_2_delay_4_52;
  reg                 io_A_Valid_2_delay_5_51;
  reg                 io_A_Valid_2_delay_6_50;
  reg                 io_A_Valid_2_delay_7_49;
  reg                 io_A_Valid_2_delay_8_48;
  reg                 io_A_Valid_2_delay_9_47;
  reg                 io_A_Valid_2_delay_10_46;
  reg                 io_A_Valid_2_delay_11_45;
  reg                 io_A_Valid_2_delay_12_44;
  reg                 io_A_Valid_2_delay_13_43;
  reg                 io_A_Valid_2_delay_14_42;
  reg                 io_A_Valid_2_delay_15_41;
  reg                 io_A_Valid_2_delay_16_40;
  reg                 io_A_Valid_2_delay_17_39;
  reg                 io_A_Valid_2_delay_18_38;
  reg                 io_A_Valid_2_delay_19_37;
  reg                 io_A_Valid_2_delay_20_36;
  reg                 io_A_Valid_2_delay_21_35;
  reg                 io_A_Valid_2_delay_22_34;
  reg                 io_A_Valid_2_delay_23_33;
  reg                 io_A_Valid_2_delay_24_32;
  reg                 io_A_Valid_2_delay_25_31;
  reg                 io_A_Valid_2_delay_26_30;
  reg                 io_A_Valid_2_delay_27_29;
  reg                 io_A_Valid_2_delay_28_28;
  reg                 io_A_Valid_2_delay_29_27;
  reg                 io_A_Valid_2_delay_30_26;
  reg                 io_A_Valid_2_delay_31_25;
  reg                 io_A_Valid_2_delay_32_24;
  reg                 io_A_Valid_2_delay_33_23;
  reg                 io_A_Valid_2_delay_34_22;
  reg                 io_A_Valid_2_delay_35_21;
  reg                 io_A_Valid_2_delay_36_20;
  reg                 io_A_Valid_2_delay_37_19;
  reg                 io_A_Valid_2_delay_38_18;
  reg                 io_A_Valid_2_delay_39_17;
  reg                 io_A_Valid_2_delay_40_16;
  reg                 io_A_Valid_2_delay_41_15;
  reg                 io_A_Valid_2_delay_42_14;
  reg                 io_A_Valid_2_delay_43_13;
  reg                 io_A_Valid_2_delay_44_12;
  reg                 io_A_Valid_2_delay_45_11;
  reg                 io_A_Valid_2_delay_46_10;
  reg                 io_A_Valid_2_delay_47_9;
  reg                 io_A_Valid_2_delay_48_8;
  reg                 io_A_Valid_2_delay_49_7;
  reg                 io_A_Valid_2_delay_50_6;
  reg                 io_A_Valid_2_delay_51_5;
  reg                 io_A_Valid_2_delay_52_4;
  reg                 io_A_Valid_2_delay_53_3;
  reg                 io_A_Valid_2_delay_54_2;
  reg                 io_A_Valid_2_delay_55_1;
  reg                 io_A_Valid_2_delay_56;
  reg                 io_B_Valid_56_delay_1_1;
  reg                 io_B_Valid_56_delay_2;
  reg                 io_A_Valid_2_delay_1_56;
  reg                 io_A_Valid_2_delay_2_55;
  reg                 io_A_Valid_2_delay_3_54;
  reg                 io_A_Valid_2_delay_4_53;
  reg                 io_A_Valid_2_delay_5_52;
  reg                 io_A_Valid_2_delay_6_51;
  reg                 io_A_Valid_2_delay_7_50;
  reg                 io_A_Valid_2_delay_8_49;
  reg                 io_A_Valid_2_delay_9_48;
  reg                 io_A_Valid_2_delay_10_47;
  reg                 io_A_Valid_2_delay_11_46;
  reg                 io_A_Valid_2_delay_12_45;
  reg                 io_A_Valid_2_delay_13_44;
  reg                 io_A_Valid_2_delay_14_43;
  reg                 io_A_Valid_2_delay_15_42;
  reg                 io_A_Valid_2_delay_16_41;
  reg                 io_A_Valid_2_delay_17_40;
  reg                 io_A_Valid_2_delay_18_39;
  reg                 io_A_Valid_2_delay_19_38;
  reg                 io_A_Valid_2_delay_20_37;
  reg                 io_A_Valid_2_delay_21_36;
  reg                 io_A_Valid_2_delay_22_35;
  reg                 io_A_Valid_2_delay_23_34;
  reg                 io_A_Valid_2_delay_24_33;
  reg                 io_A_Valid_2_delay_25_32;
  reg                 io_A_Valid_2_delay_26_31;
  reg                 io_A_Valid_2_delay_27_30;
  reg                 io_A_Valid_2_delay_28_29;
  reg                 io_A_Valid_2_delay_29_28;
  reg                 io_A_Valid_2_delay_30_27;
  reg                 io_A_Valid_2_delay_31_26;
  reg                 io_A_Valid_2_delay_32_25;
  reg                 io_A_Valid_2_delay_33_24;
  reg                 io_A_Valid_2_delay_34_23;
  reg                 io_A_Valid_2_delay_35_22;
  reg                 io_A_Valid_2_delay_36_21;
  reg                 io_A_Valid_2_delay_37_20;
  reg                 io_A_Valid_2_delay_38_19;
  reg                 io_A_Valid_2_delay_39_18;
  reg                 io_A_Valid_2_delay_40_17;
  reg                 io_A_Valid_2_delay_41_16;
  reg                 io_A_Valid_2_delay_42_15;
  reg                 io_A_Valid_2_delay_43_14;
  reg                 io_A_Valid_2_delay_44_13;
  reg                 io_A_Valid_2_delay_45_12;
  reg                 io_A_Valid_2_delay_46_11;
  reg                 io_A_Valid_2_delay_47_10;
  reg                 io_A_Valid_2_delay_48_9;
  reg                 io_A_Valid_2_delay_49_8;
  reg                 io_A_Valid_2_delay_50_7;
  reg                 io_A_Valid_2_delay_51_6;
  reg                 io_A_Valid_2_delay_52_5;
  reg                 io_A_Valid_2_delay_53_4;
  reg                 io_A_Valid_2_delay_54_3;
  reg                 io_A_Valid_2_delay_55_2;
  reg                 io_A_Valid_2_delay_56_1;
  reg                 io_A_Valid_2_delay_57;
  reg                 io_B_Valid_57_delay_1_1;
  reg                 io_B_Valid_57_delay_2;
  reg                 io_A_Valid_2_delay_1_57;
  reg                 io_A_Valid_2_delay_2_56;
  reg                 io_A_Valid_2_delay_3_55;
  reg                 io_A_Valid_2_delay_4_54;
  reg                 io_A_Valid_2_delay_5_53;
  reg                 io_A_Valid_2_delay_6_52;
  reg                 io_A_Valid_2_delay_7_51;
  reg                 io_A_Valid_2_delay_8_50;
  reg                 io_A_Valid_2_delay_9_49;
  reg                 io_A_Valid_2_delay_10_48;
  reg                 io_A_Valid_2_delay_11_47;
  reg                 io_A_Valid_2_delay_12_46;
  reg                 io_A_Valid_2_delay_13_45;
  reg                 io_A_Valid_2_delay_14_44;
  reg                 io_A_Valid_2_delay_15_43;
  reg                 io_A_Valid_2_delay_16_42;
  reg                 io_A_Valid_2_delay_17_41;
  reg                 io_A_Valid_2_delay_18_40;
  reg                 io_A_Valid_2_delay_19_39;
  reg                 io_A_Valid_2_delay_20_38;
  reg                 io_A_Valid_2_delay_21_37;
  reg                 io_A_Valid_2_delay_22_36;
  reg                 io_A_Valid_2_delay_23_35;
  reg                 io_A_Valid_2_delay_24_34;
  reg                 io_A_Valid_2_delay_25_33;
  reg                 io_A_Valid_2_delay_26_32;
  reg                 io_A_Valid_2_delay_27_31;
  reg                 io_A_Valid_2_delay_28_30;
  reg                 io_A_Valid_2_delay_29_29;
  reg                 io_A_Valid_2_delay_30_28;
  reg                 io_A_Valid_2_delay_31_27;
  reg                 io_A_Valid_2_delay_32_26;
  reg                 io_A_Valid_2_delay_33_25;
  reg                 io_A_Valid_2_delay_34_24;
  reg                 io_A_Valid_2_delay_35_23;
  reg                 io_A_Valid_2_delay_36_22;
  reg                 io_A_Valid_2_delay_37_21;
  reg                 io_A_Valid_2_delay_38_20;
  reg                 io_A_Valid_2_delay_39_19;
  reg                 io_A_Valid_2_delay_40_18;
  reg                 io_A_Valid_2_delay_41_17;
  reg                 io_A_Valid_2_delay_42_16;
  reg                 io_A_Valid_2_delay_43_15;
  reg                 io_A_Valid_2_delay_44_14;
  reg                 io_A_Valid_2_delay_45_13;
  reg                 io_A_Valid_2_delay_46_12;
  reg                 io_A_Valid_2_delay_47_11;
  reg                 io_A_Valid_2_delay_48_10;
  reg                 io_A_Valid_2_delay_49_9;
  reg                 io_A_Valid_2_delay_50_8;
  reg                 io_A_Valid_2_delay_51_7;
  reg                 io_A_Valid_2_delay_52_6;
  reg                 io_A_Valid_2_delay_53_5;
  reg                 io_A_Valid_2_delay_54_4;
  reg                 io_A_Valid_2_delay_55_3;
  reg                 io_A_Valid_2_delay_56_2;
  reg                 io_A_Valid_2_delay_57_1;
  reg                 io_A_Valid_2_delay_58;
  reg                 io_B_Valid_58_delay_1_1;
  reg                 io_B_Valid_58_delay_2;
  reg                 io_A_Valid_2_delay_1_58;
  reg                 io_A_Valid_2_delay_2_57;
  reg                 io_A_Valid_2_delay_3_56;
  reg                 io_A_Valid_2_delay_4_55;
  reg                 io_A_Valid_2_delay_5_54;
  reg                 io_A_Valid_2_delay_6_53;
  reg                 io_A_Valid_2_delay_7_52;
  reg                 io_A_Valid_2_delay_8_51;
  reg                 io_A_Valid_2_delay_9_50;
  reg                 io_A_Valid_2_delay_10_49;
  reg                 io_A_Valid_2_delay_11_48;
  reg                 io_A_Valid_2_delay_12_47;
  reg                 io_A_Valid_2_delay_13_46;
  reg                 io_A_Valid_2_delay_14_45;
  reg                 io_A_Valid_2_delay_15_44;
  reg                 io_A_Valid_2_delay_16_43;
  reg                 io_A_Valid_2_delay_17_42;
  reg                 io_A_Valid_2_delay_18_41;
  reg                 io_A_Valid_2_delay_19_40;
  reg                 io_A_Valid_2_delay_20_39;
  reg                 io_A_Valid_2_delay_21_38;
  reg                 io_A_Valid_2_delay_22_37;
  reg                 io_A_Valid_2_delay_23_36;
  reg                 io_A_Valid_2_delay_24_35;
  reg                 io_A_Valid_2_delay_25_34;
  reg                 io_A_Valid_2_delay_26_33;
  reg                 io_A_Valid_2_delay_27_32;
  reg                 io_A_Valid_2_delay_28_31;
  reg                 io_A_Valid_2_delay_29_30;
  reg                 io_A_Valid_2_delay_30_29;
  reg                 io_A_Valid_2_delay_31_28;
  reg                 io_A_Valid_2_delay_32_27;
  reg                 io_A_Valid_2_delay_33_26;
  reg                 io_A_Valid_2_delay_34_25;
  reg                 io_A_Valid_2_delay_35_24;
  reg                 io_A_Valid_2_delay_36_23;
  reg                 io_A_Valid_2_delay_37_22;
  reg                 io_A_Valid_2_delay_38_21;
  reg                 io_A_Valid_2_delay_39_20;
  reg                 io_A_Valid_2_delay_40_19;
  reg                 io_A_Valid_2_delay_41_18;
  reg                 io_A_Valid_2_delay_42_17;
  reg                 io_A_Valid_2_delay_43_16;
  reg                 io_A_Valid_2_delay_44_15;
  reg                 io_A_Valid_2_delay_45_14;
  reg                 io_A_Valid_2_delay_46_13;
  reg                 io_A_Valid_2_delay_47_12;
  reg                 io_A_Valid_2_delay_48_11;
  reg                 io_A_Valid_2_delay_49_10;
  reg                 io_A_Valid_2_delay_50_9;
  reg                 io_A_Valid_2_delay_51_8;
  reg                 io_A_Valid_2_delay_52_7;
  reg                 io_A_Valid_2_delay_53_6;
  reg                 io_A_Valid_2_delay_54_5;
  reg                 io_A_Valid_2_delay_55_4;
  reg                 io_A_Valid_2_delay_56_3;
  reg                 io_A_Valid_2_delay_57_2;
  reg                 io_A_Valid_2_delay_58_1;
  reg                 io_A_Valid_2_delay_59;
  reg                 io_B_Valid_59_delay_1_1;
  reg                 io_B_Valid_59_delay_2;
  reg                 io_A_Valid_2_delay_1_59;
  reg                 io_A_Valid_2_delay_2_58;
  reg                 io_A_Valid_2_delay_3_57;
  reg                 io_A_Valid_2_delay_4_56;
  reg                 io_A_Valid_2_delay_5_55;
  reg                 io_A_Valid_2_delay_6_54;
  reg                 io_A_Valid_2_delay_7_53;
  reg                 io_A_Valid_2_delay_8_52;
  reg                 io_A_Valid_2_delay_9_51;
  reg                 io_A_Valid_2_delay_10_50;
  reg                 io_A_Valid_2_delay_11_49;
  reg                 io_A_Valid_2_delay_12_48;
  reg                 io_A_Valid_2_delay_13_47;
  reg                 io_A_Valid_2_delay_14_46;
  reg                 io_A_Valid_2_delay_15_45;
  reg                 io_A_Valid_2_delay_16_44;
  reg                 io_A_Valid_2_delay_17_43;
  reg                 io_A_Valid_2_delay_18_42;
  reg                 io_A_Valid_2_delay_19_41;
  reg                 io_A_Valid_2_delay_20_40;
  reg                 io_A_Valid_2_delay_21_39;
  reg                 io_A_Valid_2_delay_22_38;
  reg                 io_A_Valid_2_delay_23_37;
  reg                 io_A_Valid_2_delay_24_36;
  reg                 io_A_Valid_2_delay_25_35;
  reg                 io_A_Valid_2_delay_26_34;
  reg                 io_A_Valid_2_delay_27_33;
  reg                 io_A_Valid_2_delay_28_32;
  reg                 io_A_Valid_2_delay_29_31;
  reg                 io_A_Valid_2_delay_30_30;
  reg                 io_A_Valid_2_delay_31_29;
  reg                 io_A_Valid_2_delay_32_28;
  reg                 io_A_Valid_2_delay_33_27;
  reg                 io_A_Valid_2_delay_34_26;
  reg                 io_A_Valid_2_delay_35_25;
  reg                 io_A_Valid_2_delay_36_24;
  reg                 io_A_Valid_2_delay_37_23;
  reg                 io_A_Valid_2_delay_38_22;
  reg                 io_A_Valid_2_delay_39_21;
  reg                 io_A_Valid_2_delay_40_20;
  reg                 io_A_Valid_2_delay_41_19;
  reg                 io_A_Valid_2_delay_42_18;
  reg                 io_A_Valid_2_delay_43_17;
  reg                 io_A_Valid_2_delay_44_16;
  reg                 io_A_Valid_2_delay_45_15;
  reg                 io_A_Valid_2_delay_46_14;
  reg                 io_A_Valid_2_delay_47_13;
  reg                 io_A_Valid_2_delay_48_12;
  reg                 io_A_Valid_2_delay_49_11;
  reg                 io_A_Valid_2_delay_50_10;
  reg                 io_A_Valid_2_delay_51_9;
  reg                 io_A_Valid_2_delay_52_8;
  reg                 io_A_Valid_2_delay_53_7;
  reg                 io_A_Valid_2_delay_54_6;
  reg                 io_A_Valid_2_delay_55_5;
  reg                 io_A_Valid_2_delay_56_4;
  reg                 io_A_Valid_2_delay_57_3;
  reg                 io_A_Valid_2_delay_58_2;
  reg                 io_A_Valid_2_delay_59_1;
  reg                 io_A_Valid_2_delay_60;
  reg                 io_B_Valid_60_delay_1_1;
  reg                 io_B_Valid_60_delay_2;
  reg                 io_A_Valid_2_delay_1_60;
  reg                 io_A_Valid_2_delay_2_59;
  reg                 io_A_Valid_2_delay_3_58;
  reg                 io_A_Valid_2_delay_4_57;
  reg                 io_A_Valid_2_delay_5_56;
  reg                 io_A_Valid_2_delay_6_55;
  reg                 io_A_Valid_2_delay_7_54;
  reg                 io_A_Valid_2_delay_8_53;
  reg                 io_A_Valid_2_delay_9_52;
  reg                 io_A_Valid_2_delay_10_51;
  reg                 io_A_Valid_2_delay_11_50;
  reg                 io_A_Valid_2_delay_12_49;
  reg                 io_A_Valid_2_delay_13_48;
  reg                 io_A_Valid_2_delay_14_47;
  reg                 io_A_Valid_2_delay_15_46;
  reg                 io_A_Valid_2_delay_16_45;
  reg                 io_A_Valid_2_delay_17_44;
  reg                 io_A_Valid_2_delay_18_43;
  reg                 io_A_Valid_2_delay_19_42;
  reg                 io_A_Valid_2_delay_20_41;
  reg                 io_A_Valid_2_delay_21_40;
  reg                 io_A_Valid_2_delay_22_39;
  reg                 io_A_Valid_2_delay_23_38;
  reg                 io_A_Valid_2_delay_24_37;
  reg                 io_A_Valid_2_delay_25_36;
  reg                 io_A_Valid_2_delay_26_35;
  reg                 io_A_Valid_2_delay_27_34;
  reg                 io_A_Valid_2_delay_28_33;
  reg                 io_A_Valid_2_delay_29_32;
  reg                 io_A_Valid_2_delay_30_31;
  reg                 io_A_Valid_2_delay_31_30;
  reg                 io_A_Valid_2_delay_32_29;
  reg                 io_A_Valid_2_delay_33_28;
  reg                 io_A_Valid_2_delay_34_27;
  reg                 io_A_Valid_2_delay_35_26;
  reg                 io_A_Valid_2_delay_36_25;
  reg                 io_A_Valid_2_delay_37_24;
  reg                 io_A_Valid_2_delay_38_23;
  reg                 io_A_Valid_2_delay_39_22;
  reg                 io_A_Valid_2_delay_40_21;
  reg                 io_A_Valid_2_delay_41_20;
  reg                 io_A_Valid_2_delay_42_19;
  reg                 io_A_Valid_2_delay_43_18;
  reg                 io_A_Valid_2_delay_44_17;
  reg                 io_A_Valid_2_delay_45_16;
  reg                 io_A_Valid_2_delay_46_15;
  reg                 io_A_Valid_2_delay_47_14;
  reg                 io_A_Valid_2_delay_48_13;
  reg                 io_A_Valid_2_delay_49_12;
  reg                 io_A_Valid_2_delay_50_11;
  reg                 io_A_Valid_2_delay_51_10;
  reg                 io_A_Valid_2_delay_52_9;
  reg                 io_A_Valid_2_delay_53_8;
  reg                 io_A_Valid_2_delay_54_7;
  reg                 io_A_Valid_2_delay_55_6;
  reg                 io_A_Valid_2_delay_56_5;
  reg                 io_A_Valid_2_delay_57_4;
  reg                 io_A_Valid_2_delay_58_3;
  reg                 io_A_Valid_2_delay_59_2;
  reg                 io_A_Valid_2_delay_60_1;
  reg                 io_A_Valid_2_delay_61;
  reg                 io_B_Valid_61_delay_1_1;
  reg                 io_B_Valid_61_delay_2;
  reg                 io_A_Valid_2_delay_1_61;
  reg                 io_A_Valid_2_delay_2_60;
  reg                 io_A_Valid_2_delay_3_59;
  reg                 io_A_Valid_2_delay_4_58;
  reg                 io_A_Valid_2_delay_5_57;
  reg                 io_A_Valid_2_delay_6_56;
  reg                 io_A_Valid_2_delay_7_55;
  reg                 io_A_Valid_2_delay_8_54;
  reg                 io_A_Valid_2_delay_9_53;
  reg                 io_A_Valid_2_delay_10_52;
  reg                 io_A_Valid_2_delay_11_51;
  reg                 io_A_Valid_2_delay_12_50;
  reg                 io_A_Valid_2_delay_13_49;
  reg                 io_A_Valid_2_delay_14_48;
  reg                 io_A_Valid_2_delay_15_47;
  reg                 io_A_Valid_2_delay_16_46;
  reg                 io_A_Valid_2_delay_17_45;
  reg                 io_A_Valid_2_delay_18_44;
  reg                 io_A_Valid_2_delay_19_43;
  reg                 io_A_Valid_2_delay_20_42;
  reg                 io_A_Valid_2_delay_21_41;
  reg                 io_A_Valid_2_delay_22_40;
  reg                 io_A_Valid_2_delay_23_39;
  reg                 io_A_Valid_2_delay_24_38;
  reg                 io_A_Valid_2_delay_25_37;
  reg                 io_A_Valid_2_delay_26_36;
  reg                 io_A_Valid_2_delay_27_35;
  reg                 io_A_Valid_2_delay_28_34;
  reg                 io_A_Valid_2_delay_29_33;
  reg                 io_A_Valid_2_delay_30_32;
  reg                 io_A_Valid_2_delay_31_31;
  reg                 io_A_Valid_2_delay_32_30;
  reg                 io_A_Valid_2_delay_33_29;
  reg                 io_A_Valid_2_delay_34_28;
  reg                 io_A_Valid_2_delay_35_27;
  reg                 io_A_Valid_2_delay_36_26;
  reg                 io_A_Valid_2_delay_37_25;
  reg                 io_A_Valid_2_delay_38_24;
  reg                 io_A_Valid_2_delay_39_23;
  reg                 io_A_Valid_2_delay_40_22;
  reg                 io_A_Valid_2_delay_41_21;
  reg                 io_A_Valid_2_delay_42_20;
  reg                 io_A_Valid_2_delay_43_19;
  reg                 io_A_Valid_2_delay_44_18;
  reg                 io_A_Valid_2_delay_45_17;
  reg                 io_A_Valid_2_delay_46_16;
  reg                 io_A_Valid_2_delay_47_15;
  reg                 io_A_Valid_2_delay_48_14;
  reg                 io_A_Valid_2_delay_49_13;
  reg                 io_A_Valid_2_delay_50_12;
  reg                 io_A_Valid_2_delay_51_11;
  reg                 io_A_Valid_2_delay_52_10;
  reg                 io_A_Valid_2_delay_53_9;
  reg                 io_A_Valid_2_delay_54_8;
  reg                 io_A_Valid_2_delay_55_7;
  reg                 io_A_Valid_2_delay_56_6;
  reg                 io_A_Valid_2_delay_57_5;
  reg                 io_A_Valid_2_delay_58_4;
  reg                 io_A_Valid_2_delay_59_3;
  reg                 io_A_Valid_2_delay_60_2;
  reg                 io_A_Valid_2_delay_61_1;
  reg                 io_A_Valid_2_delay_62;
  reg                 io_B_Valid_62_delay_1_1;
  reg                 io_B_Valid_62_delay_2;
  reg                 io_A_Valid_2_delay_1_62;
  reg                 io_A_Valid_2_delay_2_61;
  reg                 io_A_Valid_2_delay_3_60;
  reg                 io_A_Valid_2_delay_4_59;
  reg                 io_A_Valid_2_delay_5_58;
  reg                 io_A_Valid_2_delay_6_57;
  reg                 io_A_Valid_2_delay_7_56;
  reg                 io_A_Valid_2_delay_8_55;
  reg                 io_A_Valid_2_delay_9_54;
  reg                 io_A_Valid_2_delay_10_53;
  reg                 io_A_Valid_2_delay_11_52;
  reg                 io_A_Valid_2_delay_12_51;
  reg                 io_A_Valid_2_delay_13_50;
  reg                 io_A_Valid_2_delay_14_49;
  reg                 io_A_Valid_2_delay_15_48;
  reg                 io_A_Valid_2_delay_16_47;
  reg                 io_A_Valid_2_delay_17_46;
  reg                 io_A_Valid_2_delay_18_45;
  reg                 io_A_Valid_2_delay_19_44;
  reg                 io_A_Valid_2_delay_20_43;
  reg                 io_A_Valid_2_delay_21_42;
  reg                 io_A_Valid_2_delay_22_41;
  reg                 io_A_Valid_2_delay_23_40;
  reg                 io_A_Valid_2_delay_24_39;
  reg                 io_A_Valid_2_delay_25_38;
  reg                 io_A_Valid_2_delay_26_37;
  reg                 io_A_Valid_2_delay_27_36;
  reg                 io_A_Valid_2_delay_28_35;
  reg                 io_A_Valid_2_delay_29_34;
  reg                 io_A_Valid_2_delay_30_33;
  reg                 io_A_Valid_2_delay_31_32;
  reg                 io_A_Valid_2_delay_32_31;
  reg                 io_A_Valid_2_delay_33_30;
  reg                 io_A_Valid_2_delay_34_29;
  reg                 io_A_Valid_2_delay_35_28;
  reg                 io_A_Valid_2_delay_36_27;
  reg                 io_A_Valid_2_delay_37_26;
  reg                 io_A_Valid_2_delay_38_25;
  reg                 io_A_Valid_2_delay_39_24;
  reg                 io_A_Valid_2_delay_40_23;
  reg                 io_A_Valid_2_delay_41_22;
  reg                 io_A_Valid_2_delay_42_21;
  reg                 io_A_Valid_2_delay_43_20;
  reg                 io_A_Valid_2_delay_44_19;
  reg                 io_A_Valid_2_delay_45_18;
  reg                 io_A_Valid_2_delay_46_17;
  reg                 io_A_Valid_2_delay_47_16;
  reg                 io_A_Valid_2_delay_48_15;
  reg                 io_A_Valid_2_delay_49_14;
  reg                 io_A_Valid_2_delay_50_13;
  reg                 io_A_Valid_2_delay_51_12;
  reg                 io_A_Valid_2_delay_52_11;
  reg                 io_A_Valid_2_delay_53_10;
  reg                 io_A_Valid_2_delay_54_9;
  reg                 io_A_Valid_2_delay_55_8;
  reg                 io_A_Valid_2_delay_56_7;
  reg                 io_A_Valid_2_delay_57_6;
  reg                 io_A_Valid_2_delay_58_5;
  reg                 io_A_Valid_2_delay_59_4;
  reg                 io_A_Valid_2_delay_60_3;
  reg                 io_A_Valid_2_delay_61_2;
  reg                 io_A_Valid_2_delay_62_1;
  reg                 io_A_Valid_2_delay_63;
  reg                 io_B_Valid_63_delay_1_1;
  reg                 io_B_Valid_63_delay_2;
  reg        [15:0]   io_signCount_regNextWhen_3;
  reg                 io_B_Valid_0_delay_1_2;
  reg                 io_B_Valid_0_delay_2_1;
  reg                 io_B_Valid_0_delay_3;
  reg                 io_A_Valid_3_delay_1;
  reg                 io_B_Valid_1_delay_1_2;
  reg                 io_B_Valid_1_delay_2_1;
  reg                 io_B_Valid_1_delay_3;
  reg                 io_A_Valid_3_delay_1_1;
  reg                 io_A_Valid_3_delay_2;
  reg                 io_B_Valid_2_delay_1_2;
  reg                 io_B_Valid_2_delay_2_1;
  reg                 io_B_Valid_2_delay_3;
  reg                 io_A_Valid_3_delay_1_2;
  reg                 io_A_Valid_3_delay_2_1;
  reg                 io_A_Valid_3_delay_3;
  reg                 io_B_Valid_3_delay_1_2;
  reg                 io_B_Valid_3_delay_2_1;
  reg                 io_B_Valid_3_delay_3;
  reg                 io_A_Valid_3_delay_1_3;
  reg                 io_A_Valid_3_delay_2_2;
  reg                 io_A_Valid_3_delay_3_1;
  reg                 io_A_Valid_3_delay_4;
  reg                 io_B_Valid_4_delay_1_2;
  reg                 io_B_Valid_4_delay_2_1;
  reg                 io_B_Valid_4_delay_3;
  reg                 io_A_Valid_3_delay_1_4;
  reg                 io_A_Valid_3_delay_2_3;
  reg                 io_A_Valid_3_delay_3_2;
  reg                 io_A_Valid_3_delay_4_1;
  reg                 io_A_Valid_3_delay_5;
  reg                 io_B_Valid_5_delay_1_2;
  reg                 io_B_Valid_5_delay_2_1;
  reg                 io_B_Valid_5_delay_3;
  reg                 io_A_Valid_3_delay_1_5;
  reg                 io_A_Valid_3_delay_2_4;
  reg                 io_A_Valid_3_delay_3_3;
  reg                 io_A_Valid_3_delay_4_2;
  reg                 io_A_Valid_3_delay_5_1;
  reg                 io_A_Valid_3_delay_6;
  reg                 io_B_Valid_6_delay_1_2;
  reg                 io_B_Valid_6_delay_2_1;
  reg                 io_B_Valid_6_delay_3;
  reg                 io_A_Valid_3_delay_1_6;
  reg                 io_A_Valid_3_delay_2_5;
  reg                 io_A_Valid_3_delay_3_4;
  reg                 io_A_Valid_3_delay_4_3;
  reg                 io_A_Valid_3_delay_5_2;
  reg                 io_A_Valid_3_delay_6_1;
  reg                 io_A_Valid_3_delay_7;
  reg                 io_B_Valid_7_delay_1_2;
  reg                 io_B_Valid_7_delay_2_1;
  reg                 io_B_Valid_7_delay_3;
  reg                 io_A_Valid_3_delay_1_7;
  reg                 io_A_Valid_3_delay_2_6;
  reg                 io_A_Valid_3_delay_3_5;
  reg                 io_A_Valid_3_delay_4_4;
  reg                 io_A_Valid_3_delay_5_3;
  reg                 io_A_Valid_3_delay_6_2;
  reg                 io_A_Valid_3_delay_7_1;
  reg                 io_A_Valid_3_delay_8;
  reg                 io_B_Valid_8_delay_1_2;
  reg                 io_B_Valid_8_delay_2_1;
  reg                 io_B_Valid_8_delay_3;
  reg                 io_A_Valid_3_delay_1_8;
  reg                 io_A_Valid_3_delay_2_7;
  reg                 io_A_Valid_3_delay_3_6;
  reg                 io_A_Valid_3_delay_4_5;
  reg                 io_A_Valid_3_delay_5_4;
  reg                 io_A_Valid_3_delay_6_3;
  reg                 io_A_Valid_3_delay_7_2;
  reg                 io_A_Valid_3_delay_8_1;
  reg                 io_A_Valid_3_delay_9;
  reg                 io_B_Valid_9_delay_1_2;
  reg                 io_B_Valid_9_delay_2_1;
  reg                 io_B_Valid_9_delay_3;
  reg                 io_A_Valid_3_delay_1_9;
  reg                 io_A_Valid_3_delay_2_8;
  reg                 io_A_Valid_3_delay_3_7;
  reg                 io_A_Valid_3_delay_4_6;
  reg                 io_A_Valid_3_delay_5_5;
  reg                 io_A_Valid_3_delay_6_4;
  reg                 io_A_Valid_3_delay_7_3;
  reg                 io_A_Valid_3_delay_8_2;
  reg                 io_A_Valid_3_delay_9_1;
  reg                 io_A_Valid_3_delay_10;
  reg                 io_B_Valid_10_delay_1_2;
  reg                 io_B_Valid_10_delay_2_1;
  reg                 io_B_Valid_10_delay_3;
  reg                 io_A_Valid_3_delay_1_10;
  reg                 io_A_Valid_3_delay_2_9;
  reg                 io_A_Valid_3_delay_3_8;
  reg                 io_A_Valid_3_delay_4_7;
  reg                 io_A_Valid_3_delay_5_6;
  reg                 io_A_Valid_3_delay_6_5;
  reg                 io_A_Valid_3_delay_7_4;
  reg                 io_A_Valid_3_delay_8_3;
  reg                 io_A_Valid_3_delay_9_2;
  reg                 io_A_Valid_3_delay_10_1;
  reg                 io_A_Valid_3_delay_11;
  reg                 io_B_Valid_11_delay_1_2;
  reg                 io_B_Valid_11_delay_2_1;
  reg                 io_B_Valid_11_delay_3;
  reg                 io_A_Valid_3_delay_1_11;
  reg                 io_A_Valid_3_delay_2_10;
  reg                 io_A_Valid_3_delay_3_9;
  reg                 io_A_Valid_3_delay_4_8;
  reg                 io_A_Valid_3_delay_5_7;
  reg                 io_A_Valid_3_delay_6_6;
  reg                 io_A_Valid_3_delay_7_5;
  reg                 io_A_Valid_3_delay_8_4;
  reg                 io_A_Valid_3_delay_9_3;
  reg                 io_A_Valid_3_delay_10_2;
  reg                 io_A_Valid_3_delay_11_1;
  reg                 io_A_Valid_3_delay_12;
  reg                 io_B_Valid_12_delay_1_2;
  reg                 io_B_Valid_12_delay_2_1;
  reg                 io_B_Valid_12_delay_3;
  reg                 io_A_Valid_3_delay_1_12;
  reg                 io_A_Valid_3_delay_2_11;
  reg                 io_A_Valid_3_delay_3_10;
  reg                 io_A_Valid_3_delay_4_9;
  reg                 io_A_Valid_3_delay_5_8;
  reg                 io_A_Valid_3_delay_6_7;
  reg                 io_A_Valid_3_delay_7_6;
  reg                 io_A_Valid_3_delay_8_5;
  reg                 io_A_Valid_3_delay_9_4;
  reg                 io_A_Valid_3_delay_10_3;
  reg                 io_A_Valid_3_delay_11_2;
  reg                 io_A_Valid_3_delay_12_1;
  reg                 io_A_Valid_3_delay_13;
  reg                 io_B_Valid_13_delay_1_2;
  reg                 io_B_Valid_13_delay_2_1;
  reg                 io_B_Valid_13_delay_3;
  reg                 io_A_Valid_3_delay_1_13;
  reg                 io_A_Valid_3_delay_2_12;
  reg                 io_A_Valid_3_delay_3_11;
  reg                 io_A_Valid_3_delay_4_10;
  reg                 io_A_Valid_3_delay_5_9;
  reg                 io_A_Valid_3_delay_6_8;
  reg                 io_A_Valid_3_delay_7_7;
  reg                 io_A_Valid_3_delay_8_6;
  reg                 io_A_Valid_3_delay_9_5;
  reg                 io_A_Valid_3_delay_10_4;
  reg                 io_A_Valid_3_delay_11_3;
  reg                 io_A_Valid_3_delay_12_2;
  reg                 io_A_Valid_3_delay_13_1;
  reg                 io_A_Valid_3_delay_14;
  reg                 io_B_Valid_14_delay_1_2;
  reg                 io_B_Valid_14_delay_2_1;
  reg                 io_B_Valid_14_delay_3;
  reg                 io_A_Valid_3_delay_1_14;
  reg                 io_A_Valid_3_delay_2_13;
  reg                 io_A_Valid_3_delay_3_12;
  reg                 io_A_Valid_3_delay_4_11;
  reg                 io_A_Valid_3_delay_5_10;
  reg                 io_A_Valid_3_delay_6_9;
  reg                 io_A_Valid_3_delay_7_8;
  reg                 io_A_Valid_3_delay_8_7;
  reg                 io_A_Valid_3_delay_9_6;
  reg                 io_A_Valid_3_delay_10_5;
  reg                 io_A_Valid_3_delay_11_4;
  reg                 io_A_Valid_3_delay_12_3;
  reg                 io_A_Valid_3_delay_13_2;
  reg                 io_A_Valid_3_delay_14_1;
  reg                 io_A_Valid_3_delay_15;
  reg                 io_B_Valid_15_delay_1_2;
  reg                 io_B_Valid_15_delay_2_1;
  reg                 io_B_Valid_15_delay_3;
  reg                 io_A_Valid_3_delay_1_15;
  reg                 io_A_Valid_3_delay_2_14;
  reg                 io_A_Valid_3_delay_3_13;
  reg                 io_A_Valid_3_delay_4_12;
  reg                 io_A_Valid_3_delay_5_11;
  reg                 io_A_Valid_3_delay_6_10;
  reg                 io_A_Valid_3_delay_7_9;
  reg                 io_A_Valid_3_delay_8_8;
  reg                 io_A_Valid_3_delay_9_7;
  reg                 io_A_Valid_3_delay_10_6;
  reg                 io_A_Valid_3_delay_11_5;
  reg                 io_A_Valid_3_delay_12_4;
  reg                 io_A_Valid_3_delay_13_3;
  reg                 io_A_Valid_3_delay_14_2;
  reg                 io_A_Valid_3_delay_15_1;
  reg                 io_A_Valid_3_delay_16;
  reg                 io_B_Valid_16_delay_1_2;
  reg                 io_B_Valid_16_delay_2_1;
  reg                 io_B_Valid_16_delay_3;
  reg                 io_A_Valid_3_delay_1_16;
  reg                 io_A_Valid_3_delay_2_15;
  reg                 io_A_Valid_3_delay_3_14;
  reg                 io_A_Valid_3_delay_4_13;
  reg                 io_A_Valid_3_delay_5_12;
  reg                 io_A_Valid_3_delay_6_11;
  reg                 io_A_Valid_3_delay_7_10;
  reg                 io_A_Valid_3_delay_8_9;
  reg                 io_A_Valid_3_delay_9_8;
  reg                 io_A_Valid_3_delay_10_7;
  reg                 io_A_Valid_3_delay_11_6;
  reg                 io_A_Valid_3_delay_12_5;
  reg                 io_A_Valid_3_delay_13_4;
  reg                 io_A_Valid_3_delay_14_3;
  reg                 io_A_Valid_3_delay_15_2;
  reg                 io_A_Valid_3_delay_16_1;
  reg                 io_A_Valid_3_delay_17;
  reg                 io_B_Valid_17_delay_1_2;
  reg                 io_B_Valid_17_delay_2_1;
  reg                 io_B_Valid_17_delay_3;
  reg                 io_A_Valid_3_delay_1_17;
  reg                 io_A_Valid_3_delay_2_16;
  reg                 io_A_Valid_3_delay_3_15;
  reg                 io_A_Valid_3_delay_4_14;
  reg                 io_A_Valid_3_delay_5_13;
  reg                 io_A_Valid_3_delay_6_12;
  reg                 io_A_Valid_3_delay_7_11;
  reg                 io_A_Valid_3_delay_8_10;
  reg                 io_A_Valid_3_delay_9_9;
  reg                 io_A_Valid_3_delay_10_8;
  reg                 io_A_Valid_3_delay_11_7;
  reg                 io_A_Valid_3_delay_12_6;
  reg                 io_A_Valid_3_delay_13_5;
  reg                 io_A_Valid_3_delay_14_4;
  reg                 io_A_Valid_3_delay_15_3;
  reg                 io_A_Valid_3_delay_16_2;
  reg                 io_A_Valid_3_delay_17_1;
  reg                 io_A_Valid_3_delay_18;
  reg                 io_B_Valid_18_delay_1_2;
  reg                 io_B_Valid_18_delay_2_1;
  reg                 io_B_Valid_18_delay_3;
  reg                 io_A_Valid_3_delay_1_18;
  reg                 io_A_Valid_3_delay_2_17;
  reg                 io_A_Valid_3_delay_3_16;
  reg                 io_A_Valid_3_delay_4_15;
  reg                 io_A_Valid_3_delay_5_14;
  reg                 io_A_Valid_3_delay_6_13;
  reg                 io_A_Valid_3_delay_7_12;
  reg                 io_A_Valid_3_delay_8_11;
  reg                 io_A_Valid_3_delay_9_10;
  reg                 io_A_Valid_3_delay_10_9;
  reg                 io_A_Valid_3_delay_11_8;
  reg                 io_A_Valid_3_delay_12_7;
  reg                 io_A_Valid_3_delay_13_6;
  reg                 io_A_Valid_3_delay_14_5;
  reg                 io_A_Valid_3_delay_15_4;
  reg                 io_A_Valid_3_delay_16_3;
  reg                 io_A_Valid_3_delay_17_2;
  reg                 io_A_Valid_3_delay_18_1;
  reg                 io_A_Valid_3_delay_19;
  reg                 io_B_Valid_19_delay_1_2;
  reg                 io_B_Valid_19_delay_2_1;
  reg                 io_B_Valid_19_delay_3;
  reg                 io_A_Valid_3_delay_1_19;
  reg                 io_A_Valid_3_delay_2_18;
  reg                 io_A_Valid_3_delay_3_17;
  reg                 io_A_Valid_3_delay_4_16;
  reg                 io_A_Valid_3_delay_5_15;
  reg                 io_A_Valid_3_delay_6_14;
  reg                 io_A_Valid_3_delay_7_13;
  reg                 io_A_Valid_3_delay_8_12;
  reg                 io_A_Valid_3_delay_9_11;
  reg                 io_A_Valid_3_delay_10_10;
  reg                 io_A_Valid_3_delay_11_9;
  reg                 io_A_Valid_3_delay_12_8;
  reg                 io_A_Valid_3_delay_13_7;
  reg                 io_A_Valid_3_delay_14_6;
  reg                 io_A_Valid_3_delay_15_5;
  reg                 io_A_Valid_3_delay_16_4;
  reg                 io_A_Valid_3_delay_17_3;
  reg                 io_A_Valid_3_delay_18_2;
  reg                 io_A_Valid_3_delay_19_1;
  reg                 io_A_Valid_3_delay_20;
  reg                 io_B_Valid_20_delay_1_2;
  reg                 io_B_Valid_20_delay_2_1;
  reg                 io_B_Valid_20_delay_3;
  reg                 io_A_Valid_3_delay_1_20;
  reg                 io_A_Valid_3_delay_2_19;
  reg                 io_A_Valid_3_delay_3_18;
  reg                 io_A_Valid_3_delay_4_17;
  reg                 io_A_Valid_3_delay_5_16;
  reg                 io_A_Valid_3_delay_6_15;
  reg                 io_A_Valid_3_delay_7_14;
  reg                 io_A_Valid_3_delay_8_13;
  reg                 io_A_Valid_3_delay_9_12;
  reg                 io_A_Valid_3_delay_10_11;
  reg                 io_A_Valid_3_delay_11_10;
  reg                 io_A_Valid_3_delay_12_9;
  reg                 io_A_Valid_3_delay_13_8;
  reg                 io_A_Valid_3_delay_14_7;
  reg                 io_A_Valid_3_delay_15_6;
  reg                 io_A_Valid_3_delay_16_5;
  reg                 io_A_Valid_3_delay_17_4;
  reg                 io_A_Valid_3_delay_18_3;
  reg                 io_A_Valid_3_delay_19_2;
  reg                 io_A_Valid_3_delay_20_1;
  reg                 io_A_Valid_3_delay_21;
  reg                 io_B_Valid_21_delay_1_2;
  reg                 io_B_Valid_21_delay_2_1;
  reg                 io_B_Valid_21_delay_3;
  reg                 io_A_Valid_3_delay_1_21;
  reg                 io_A_Valid_3_delay_2_20;
  reg                 io_A_Valid_3_delay_3_19;
  reg                 io_A_Valid_3_delay_4_18;
  reg                 io_A_Valid_3_delay_5_17;
  reg                 io_A_Valid_3_delay_6_16;
  reg                 io_A_Valid_3_delay_7_15;
  reg                 io_A_Valid_3_delay_8_14;
  reg                 io_A_Valid_3_delay_9_13;
  reg                 io_A_Valid_3_delay_10_12;
  reg                 io_A_Valid_3_delay_11_11;
  reg                 io_A_Valid_3_delay_12_10;
  reg                 io_A_Valid_3_delay_13_9;
  reg                 io_A_Valid_3_delay_14_8;
  reg                 io_A_Valid_3_delay_15_7;
  reg                 io_A_Valid_3_delay_16_6;
  reg                 io_A_Valid_3_delay_17_5;
  reg                 io_A_Valid_3_delay_18_4;
  reg                 io_A_Valid_3_delay_19_3;
  reg                 io_A_Valid_3_delay_20_2;
  reg                 io_A_Valid_3_delay_21_1;
  reg                 io_A_Valid_3_delay_22;
  reg                 io_B_Valid_22_delay_1_2;
  reg                 io_B_Valid_22_delay_2_1;
  reg                 io_B_Valid_22_delay_3;
  reg                 io_A_Valid_3_delay_1_22;
  reg                 io_A_Valid_3_delay_2_21;
  reg                 io_A_Valid_3_delay_3_20;
  reg                 io_A_Valid_3_delay_4_19;
  reg                 io_A_Valid_3_delay_5_18;
  reg                 io_A_Valid_3_delay_6_17;
  reg                 io_A_Valid_3_delay_7_16;
  reg                 io_A_Valid_3_delay_8_15;
  reg                 io_A_Valid_3_delay_9_14;
  reg                 io_A_Valid_3_delay_10_13;
  reg                 io_A_Valid_3_delay_11_12;
  reg                 io_A_Valid_3_delay_12_11;
  reg                 io_A_Valid_3_delay_13_10;
  reg                 io_A_Valid_3_delay_14_9;
  reg                 io_A_Valid_3_delay_15_8;
  reg                 io_A_Valid_3_delay_16_7;
  reg                 io_A_Valid_3_delay_17_6;
  reg                 io_A_Valid_3_delay_18_5;
  reg                 io_A_Valid_3_delay_19_4;
  reg                 io_A_Valid_3_delay_20_3;
  reg                 io_A_Valid_3_delay_21_2;
  reg                 io_A_Valid_3_delay_22_1;
  reg                 io_A_Valid_3_delay_23;
  reg                 io_B_Valid_23_delay_1_2;
  reg                 io_B_Valid_23_delay_2_1;
  reg                 io_B_Valid_23_delay_3;
  reg                 io_A_Valid_3_delay_1_23;
  reg                 io_A_Valid_3_delay_2_22;
  reg                 io_A_Valid_3_delay_3_21;
  reg                 io_A_Valid_3_delay_4_20;
  reg                 io_A_Valid_3_delay_5_19;
  reg                 io_A_Valid_3_delay_6_18;
  reg                 io_A_Valid_3_delay_7_17;
  reg                 io_A_Valid_3_delay_8_16;
  reg                 io_A_Valid_3_delay_9_15;
  reg                 io_A_Valid_3_delay_10_14;
  reg                 io_A_Valid_3_delay_11_13;
  reg                 io_A_Valid_3_delay_12_12;
  reg                 io_A_Valid_3_delay_13_11;
  reg                 io_A_Valid_3_delay_14_10;
  reg                 io_A_Valid_3_delay_15_9;
  reg                 io_A_Valid_3_delay_16_8;
  reg                 io_A_Valid_3_delay_17_7;
  reg                 io_A_Valid_3_delay_18_6;
  reg                 io_A_Valid_3_delay_19_5;
  reg                 io_A_Valid_3_delay_20_4;
  reg                 io_A_Valid_3_delay_21_3;
  reg                 io_A_Valid_3_delay_22_2;
  reg                 io_A_Valid_3_delay_23_1;
  reg                 io_A_Valid_3_delay_24;
  reg                 io_B_Valid_24_delay_1_2;
  reg                 io_B_Valid_24_delay_2_1;
  reg                 io_B_Valid_24_delay_3;
  reg                 io_A_Valid_3_delay_1_24;
  reg                 io_A_Valid_3_delay_2_23;
  reg                 io_A_Valid_3_delay_3_22;
  reg                 io_A_Valid_3_delay_4_21;
  reg                 io_A_Valid_3_delay_5_20;
  reg                 io_A_Valid_3_delay_6_19;
  reg                 io_A_Valid_3_delay_7_18;
  reg                 io_A_Valid_3_delay_8_17;
  reg                 io_A_Valid_3_delay_9_16;
  reg                 io_A_Valid_3_delay_10_15;
  reg                 io_A_Valid_3_delay_11_14;
  reg                 io_A_Valid_3_delay_12_13;
  reg                 io_A_Valid_3_delay_13_12;
  reg                 io_A_Valid_3_delay_14_11;
  reg                 io_A_Valid_3_delay_15_10;
  reg                 io_A_Valid_3_delay_16_9;
  reg                 io_A_Valid_3_delay_17_8;
  reg                 io_A_Valid_3_delay_18_7;
  reg                 io_A_Valid_3_delay_19_6;
  reg                 io_A_Valid_3_delay_20_5;
  reg                 io_A_Valid_3_delay_21_4;
  reg                 io_A_Valid_3_delay_22_3;
  reg                 io_A_Valid_3_delay_23_2;
  reg                 io_A_Valid_3_delay_24_1;
  reg                 io_A_Valid_3_delay_25;
  reg                 io_B_Valid_25_delay_1_2;
  reg                 io_B_Valid_25_delay_2_1;
  reg                 io_B_Valid_25_delay_3;
  reg                 io_A_Valid_3_delay_1_25;
  reg                 io_A_Valid_3_delay_2_24;
  reg                 io_A_Valid_3_delay_3_23;
  reg                 io_A_Valid_3_delay_4_22;
  reg                 io_A_Valid_3_delay_5_21;
  reg                 io_A_Valid_3_delay_6_20;
  reg                 io_A_Valid_3_delay_7_19;
  reg                 io_A_Valid_3_delay_8_18;
  reg                 io_A_Valid_3_delay_9_17;
  reg                 io_A_Valid_3_delay_10_16;
  reg                 io_A_Valid_3_delay_11_15;
  reg                 io_A_Valid_3_delay_12_14;
  reg                 io_A_Valid_3_delay_13_13;
  reg                 io_A_Valid_3_delay_14_12;
  reg                 io_A_Valid_3_delay_15_11;
  reg                 io_A_Valid_3_delay_16_10;
  reg                 io_A_Valid_3_delay_17_9;
  reg                 io_A_Valid_3_delay_18_8;
  reg                 io_A_Valid_3_delay_19_7;
  reg                 io_A_Valid_3_delay_20_6;
  reg                 io_A_Valid_3_delay_21_5;
  reg                 io_A_Valid_3_delay_22_4;
  reg                 io_A_Valid_3_delay_23_3;
  reg                 io_A_Valid_3_delay_24_2;
  reg                 io_A_Valid_3_delay_25_1;
  reg                 io_A_Valid_3_delay_26;
  reg                 io_B_Valid_26_delay_1_2;
  reg                 io_B_Valid_26_delay_2_1;
  reg                 io_B_Valid_26_delay_3;
  reg                 io_A_Valid_3_delay_1_26;
  reg                 io_A_Valid_3_delay_2_25;
  reg                 io_A_Valid_3_delay_3_24;
  reg                 io_A_Valid_3_delay_4_23;
  reg                 io_A_Valid_3_delay_5_22;
  reg                 io_A_Valid_3_delay_6_21;
  reg                 io_A_Valid_3_delay_7_20;
  reg                 io_A_Valid_3_delay_8_19;
  reg                 io_A_Valid_3_delay_9_18;
  reg                 io_A_Valid_3_delay_10_17;
  reg                 io_A_Valid_3_delay_11_16;
  reg                 io_A_Valid_3_delay_12_15;
  reg                 io_A_Valid_3_delay_13_14;
  reg                 io_A_Valid_3_delay_14_13;
  reg                 io_A_Valid_3_delay_15_12;
  reg                 io_A_Valid_3_delay_16_11;
  reg                 io_A_Valid_3_delay_17_10;
  reg                 io_A_Valid_3_delay_18_9;
  reg                 io_A_Valid_3_delay_19_8;
  reg                 io_A_Valid_3_delay_20_7;
  reg                 io_A_Valid_3_delay_21_6;
  reg                 io_A_Valid_3_delay_22_5;
  reg                 io_A_Valid_3_delay_23_4;
  reg                 io_A_Valid_3_delay_24_3;
  reg                 io_A_Valid_3_delay_25_2;
  reg                 io_A_Valid_3_delay_26_1;
  reg                 io_A_Valid_3_delay_27;
  reg                 io_B_Valid_27_delay_1_2;
  reg                 io_B_Valid_27_delay_2_1;
  reg                 io_B_Valid_27_delay_3;
  reg                 io_A_Valid_3_delay_1_27;
  reg                 io_A_Valid_3_delay_2_26;
  reg                 io_A_Valid_3_delay_3_25;
  reg                 io_A_Valid_3_delay_4_24;
  reg                 io_A_Valid_3_delay_5_23;
  reg                 io_A_Valid_3_delay_6_22;
  reg                 io_A_Valid_3_delay_7_21;
  reg                 io_A_Valid_3_delay_8_20;
  reg                 io_A_Valid_3_delay_9_19;
  reg                 io_A_Valid_3_delay_10_18;
  reg                 io_A_Valid_3_delay_11_17;
  reg                 io_A_Valid_3_delay_12_16;
  reg                 io_A_Valid_3_delay_13_15;
  reg                 io_A_Valid_3_delay_14_14;
  reg                 io_A_Valid_3_delay_15_13;
  reg                 io_A_Valid_3_delay_16_12;
  reg                 io_A_Valid_3_delay_17_11;
  reg                 io_A_Valid_3_delay_18_10;
  reg                 io_A_Valid_3_delay_19_9;
  reg                 io_A_Valid_3_delay_20_8;
  reg                 io_A_Valid_3_delay_21_7;
  reg                 io_A_Valid_3_delay_22_6;
  reg                 io_A_Valid_3_delay_23_5;
  reg                 io_A_Valid_3_delay_24_4;
  reg                 io_A_Valid_3_delay_25_3;
  reg                 io_A_Valid_3_delay_26_2;
  reg                 io_A_Valid_3_delay_27_1;
  reg                 io_A_Valid_3_delay_28;
  reg                 io_B_Valid_28_delay_1_2;
  reg                 io_B_Valid_28_delay_2_1;
  reg                 io_B_Valid_28_delay_3;
  reg                 io_A_Valid_3_delay_1_28;
  reg                 io_A_Valid_3_delay_2_27;
  reg                 io_A_Valid_3_delay_3_26;
  reg                 io_A_Valid_3_delay_4_25;
  reg                 io_A_Valid_3_delay_5_24;
  reg                 io_A_Valid_3_delay_6_23;
  reg                 io_A_Valid_3_delay_7_22;
  reg                 io_A_Valid_3_delay_8_21;
  reg                 io_A_Valid_3_delay_9_20;
  reg                 io_A_Valid_3_delay_10_19;
  reg                 io_A_Valid_3_delay_11_18;
  reg                 io_A_Valid_3_delay_12_17;
  reg                 io_A_Valid_3_delay_13_16;
  reg                 io_A_Valid_3_delay_14_15;
  reg                 io_A_Valid_3_delay_15_14;
  reg                 io_A_Valid_3_delay_16_13;
  reg                 io_A_Valid_3_delay_17_12;
  reg                 io_A_Valid_3_delay_18_11;
  reg                 io_A_Valid_3_delay_19_10;
  reg                 io_A_Valid_3_delay_20_9;
  reg                 io_A_Valid_3_delay_21_8;
  reg                 io_A_Valid_3_delay_22_7;
  reg                 io_A_Valid_3_delay_23_6;
  reg                 io_A_Valid_3_delay_24_5;
  reg                 io_A_Valid_3_delay_25_4;
  reg                 io_A_Valid_3_delay_26_3;
  reg                 io_A_Valid_3_delay_27_2;
  reg                 io_A_Valid_3_delay_28_1;
  reg                 io_A_Valid_3_delay_29;
  reg                 io_B_Valid_29_delay_1_2;
  reg                 io_B_Valid_29_delay_2_1;
  reg                 io_B_Valid_29_delay_3;
  reg                 io_A_Valid_3_delay_1_29;
  reg                 io_A_Valid_3_delay_2_28;
  reg                 io_A_Valid_3_delay_3_27;
  reg                 io_A_Valid_3_delay_4_26;
  reg                 io_A_Valid_3_delay_5_25;
  reg                 io_A_Valid_3_delay_6_24;
  reg                 io_A_Valid_3_delay_7_23;
  reg                 io_A_Valid_3_delay_8_22;
  reg                 io_A_Valid_3_delay_9_21;
  reg                 io_A_Valid_3_delay_10_20;
  reg                 io_A_Valid_3_delay_11_19;
  reg                 io_A_Valid_3_delay_12_18;
  reg                 io_A_Valid_3_delay_13_17;
  reg                 io_A_Valid_3_delay_14_16;
  reg                 io_A_Valid_3_delay_15_15;
  reg                 io_A_Valid_3_delay_16_14;
  reg                 io_A_Valid_3_delay_17_13;
  reg                 io_A_Valid_3_delay_18_12;
  reg                 io_A_Valid_3_delay_19_11;
  reg                 io_A_Valid_3_delay_20_10;
  reg                 io_A_Valid_3_delay_21_9;
  reg                 io_A_Valid_3_delay_22_8;
  reg                 io_A_Valid_3_delay_23_7;
  reg                 io_A_Valid_3_delay_24_6;
  reg                 io_A_Valid_3_delay_25_5;
  reg                 io_A_Valid_3_delay_26_4;
  reg                 io_A_Valid_3_delay_27_3;
  reg                 io_A_Valid_3_delay_28_2;
  reg                 io_A_Valid_3_delay_29_1;
  reg                 io_A_Valid_3_delay_30;
  reg                 io_B_Valid_30_delay_1_2;
  reg                 io_B_Valid_30_delay_2_1;
  reg                 io_B_Valid_30_delay_3;
  reg                 io_A_Valid_3_delay_1_30;
  reg                 io_A_Valid_3_delay_2_29;
  reg                 io_A_Valid_3_delay_3_28;
  reg                 io_A_Valid_3_delay_4_27;
  reg                 io_A_Valid_3_delay_5_26;
  reg                 io_A_Valid_3_delay_6_25;
  reg                 io_A_Valid_3_delay_7_24;
  reg                 io_A_Valid_3_delay_8_23;
  reg                 io_A_Valid_3_delay_9_22;
  reg                 io_A_Valid_3_delay_10_21;
  reg                 io_A_Valid_3_delay_11_20;
  reg                 io_A_Valid_3_delay_12_19;
  reg                 io_A_Valid_3_delay_13_18;
  reg                 io_A_Valid_3_delay_14_17;
  reg                 io_A_Valid_3_delay_15_16;
  reg                 io_A_Valid_3_delay_16_15;
  reg                 io_A_Valid_3_delay_17_14;
  reg                 io_A_Valid_3_delay_18_13;
  reg                 io_A_Valid_3_delay_19_12;
  reg                 io_A_Valid_3_delay_20_11;
  reg                 io_A_Valid_3_delay_21_10;
  reg                 io_A_Valid_3_delay_22_9;
  reg                 io_A_Valid_3_delay_23_8;
  reg                 io_A_Valid_3_delay_24_7;
  reg                 io_A_Valid_3_delay_25_6;
  reg                 io_A_Valid_3_delay_26_5;
  reg                 io_A_Valid_3_delay_27_4;
  reg                 io_A_Valid_3_delay_28_3;
  reg                 io_A_Valid_3_delay_29_2;
  reg                 io_A_Valid_3_delay_30_1;
  reg                 io_A_Valid_3_delay_31;
  reg                 io_B_Valid_31_delay_1_2;
  reg                 io_B_Valid_31_delay_2_1;
  reg                 io_B_Valid_31_delay_3;
  reg                 io_A_Valid_3_delay_1_31;
  reg                 io_A_Valid_3_delay_2_30;
  reg                 io_A_Valid_3_delay_3_29;
  reg                 io_A_Valid_3_delay_4_28;
  reg                 io_A_Valid_3_delay_5_27;
  reg                 io_A_Valid_3_delay_6_26;
  reg                 io_A_Valid_3_delay_7_25;
  reg                 io_A_Valid_3_delay_8_24;
  reg                 io_A_Valid_3_delay_9_23;
  reg                 io_A_Valid_3_delay_10_22;
  reg                 io_A_Valid_3_delay_11_21;
  reg                 io_A_Valid_3_delay_12_20;
  reg                 io_A_Valid_3_delay_13_19;
  reg                 io_A_Valid_3_delay_14_18;
  reg                 io_A_Valid_3_delay_15_17;
  reg                 io_A_Valid_3_delay_16_16;
  reg                 io_A_Valid_3_delay_17_15;
  reg                 io_A_Valid_3_delay_18_14;
  reg                 io_A_Valid_3_delay_19_13;
  reg                 io_A_Valid_3_delay_20_12;
  reg                 io_A_Valid_3_delay_21_11;
  reg                 io_A_Valid_3_delay_22_10;
  reg                 io_A_Valid_3_delay_23_9;
  reg                 io_A_Valid_3_delay_24_8;
  reg                 io_A_Valid_3_delay_25_7;
  reg                 io_A_Valid_3_delay_26_6;
  reg                 io_A_Valid_3_delay_27_5;
  reg                 io_A_Valid_3_delay_28_4;
  reg                 io_A_Valid_3_delay_29_3;
  reg                 io_A_Valid_3_delay_30_2;
  reg                 io_A_Valid_3_delay_31_1;
  reg                 io_A_Valid_3_delay_32;
  reg                 io_B_Valid_32_delay_1_2;
  reg                 io_B_Valid_32_delay_2_1;
  reg                 io_B_Valid_32_delay_3;
  reg                 io_A_Valid_3_delay_1_32;
  reg                 io_A_Valid_3_delay_2_31;
  reg                 io_A_Valid_3_delay_3_30;
  reg                 io_A_Valid_3_delay_4_29;
  reg                 io_A_Valid_3_delay_5_28;
  reg                 io_A_Valid_3_delay_6_27;
  reg                 io_A_Valid_3_delay_7_26;
  reg                 io_A_Valid_3_delay_8_25;
  reg                 io_A_Valid_3_delay_9_24;
  reg                 io_A_Valid_3_delay_10_23;
  reg                 io_A_Valid_3_delay_11_22;
  reg                 io_A_Valid_3_delay_12_21;
  reg                 io_A_Valid_3_delay_13_20;
  reg                 io_A_Valid_3_delay_14_19;
  reg                 io_A_Valid_3_delay_15_18;
  reg                 io_A_Valid_3_delay_16_17;
  reg                 io_A_Valid_3_delay_17_16;
  reg                 io_A_Valid_3_delay_18_15;
  reg                 io_A_Valid_3_delay_19_14;
  reg                 io_A_Valid_3_delay_20_13;
  reg                 io_A_Valid_3_delay_21_12;
  reg                 io_A_Valid_3_delay_22_11;
  reg                 io_A_Valid_3_delay_23_10;
  reg                 io_A_Valid_3_delay_24_9;
  reg                 io_A_Valid_3_delay_25_8;
  reg                 io_A_Valid_3_delay_26_7;
  reg                 io_A_Valid_3_delay_27_6;
  reg                 io_A_Valid_3_delay_28_5;
  reg                 io_A_Valid_3_delay_29_4;
  reg                 io_A_Valid_3_delay_30_3;
  reg                 io_A_Valid_3_delay_31_2;
  reg                 io_A_Valid_3_delay_32_1;
  reg                 io_A_Valid_3_delay_33;
  reg                 io_B_Valid_33_delay_1_2;
  reg                 io_B_Valid_33_delay_2_1;
  reg                 io_B_Valid_33_delay_3;
  reg                 io_A_Valid_3_delay_1_33;
  reg                 io_A_Valid_3_delay_2_32;
  reg                 io_A_Valid_3_delay_3_31;
  reg                 io_A_Valid_3_delay_4_30;
  reg                 io_A_Valid_3_delay_5_29;
  reg                 io_A_Valid_3_delay_6_28;
  reg                 io_A_Valid_3_delay_7_27;
  reg                 io_A_Valid_3_delay_8_26;
  reg                 io_A_Valid_3_delay_9_25;
  reg                 io_A_Valid_3_delay_10_24;
  reg                 io_A_Valid_3_delay_11_23;
  reg                 io_A_Valid_3_delay_12_22;
  reg                 io_A_Valid_3_delay_13_21;
  reg                 io_A_Valid_3_delay_14_20;
  reg                 io_A_Valid_3_delay_15_19;
  reg                 io_A_Valid_3_delay_16_18;
  reg                 io_A_Valid_3_delay_17_17;
  reg                 io_A_Valid_3_delay_18_16;
  reg                 io_A_Valid_3_delay_19_15;
  reg                 io_A_Valid_3_delay_20_14;
  reg                 io_A_Valid_3_delay_21_13;
  reg                 io_A_Valid_3_delay_22_12;
  reg                 io_A_Valid_3_delay_23_11;
  reg                 io_A_Valid_3_delay_24_10;
  reg                 io_A_Valid_3_delay_25_9;
  reg                 io_A_Valid_3_delay_26_8;
  reg                 io_A_Valid_3_delay_27_7;
  reg                 io_A_Valid_3_delay_28_6;
  reg                 io_A_Valid_3_delay_29_5;
  reg                 io_A_Valid_3_delay_30_4;
  reg                 io_A_Valid_3_delay_31_3;
  reg                 io_A_Valid_3_delay_32_2;
  reg                 io_A_Valid_3_delay_33_1;
  reg                 io_A_Valid_3_delay_34;
  reg                 io_B_Valid_34_delay_1_2;
  reg                 io_B_Valid_34_delay_2_1;
  reg                 io_B_Valid_34_delay_3;
  reg                 io_A_Valid_3_delay_1_34;
  reg                 io_A_Valid_3_delay_2_33;
  reg                 io_A_Valid_3_delay_3_32;
  reg                 io_A_Valid_3_delay_4_31;
  reg                 io_A_Valid_3_delay_5_30;
  reg                 io_A_Valid_3_delay_6_29;
  reg                 io_A_Valid_3_delay_7_28;
  reg                 io_A_Valid_3_delay_8_27;
  reg                 io_A_Valid_3_delay_9_26;
  reg                 io_A_Valid_3_delay_10_25;
  reg                 io_A_Valid_3_delay_11_24;
  reg                 io_A_Valid_3_delay_12_23;
  reg                 io_A_Valid_3_delay_13_22;
  reg                 io_A_Valid_3_delay_14_21;
  reg                 io_A_Valid_3_delay_15_20;
  reg                 io_A_Valid_3_delay_16_19;
  reg                 io_A_Valid_3_delay_17_18;
  reg                 io_A_Valid_3_delay_18_17;
  reg                 io_A_Valid_3_delay_19_16;
  reg                 io_A_Valid_3_delay_20_15;
  reg                 io_A_Valid_3_delay_21_14;
  reg                 io_A_Valid_3_delay_22_13;
  reg                 io_A_Valid_3_delay_23_12;
  reg                 io_A_Valid_3_delay_24_11;
  reg                 io_A_Valid_3_delay_25_10;
  reg                 io_A_Valid_3_delay_26_9;
  reg                 io_A_Valid_3_delay_27_8;
  reg                 io_A_Valid_3_delay_28_7;
  reg                 io_A_Valid_3_delay_29_6;
  reg                 io_A_Valid_3_delay_30_5;
  reg                 io_A_Valid_3_delay_31_4;
  reg                 io_A_Valid_3_delay_32_3;
  reg                 io_A_Valid_3_delay_33_2;
  reg                 io_A_Valid_3_delay_34_1;
  reg                 io_A_Valid_3_delay_35;
  reg                 io_B_Valid_35_delay_1_2;
  reg                 io_B_Valid_35_delay_2_1;
  reg                 io_B_Valid_35_delay_3;
  reg                 io_A_Valid_3_delay_1_35;
  reg                 io_A_Valid_3_delay_2_34;
  reg                 io_A_Valid_3_delay_3_33;
  reg                 io_A_Valid_3_delay_4_32;
  reg                 io_A_Valid_3_delay_5_31;
  reg                 io_A_Valid_3_delay_6_30;
  reg                 io_A_Valid_3_delay_7_29;
  reg                 io_A_Valid_3_delay_8_28;
  reg                 io_A_Valid_3_delay_9_27;
  reg                 io_A_Valid_3_delay_10_26;
  reg                 io_A_Valid_3_delay_11_25;
  reg                 io_A_Valid_3_delay_12_24;
  reg                 io_A_Valid_3_delay_13_23;
  reg                 io_A_Valid_3_delay_14_22;
  reg                 io_A_Valid_3_delay_15_21;
  reg                 io_A_Valid_3_delay_16_20;
  reg                 io_A_Valid_3_delay_17_19;
  reg                 io_A_Valid_3_delay_18_18;
  reg                 io_A_Valid_3_delay_19_17;
  reg                 io_A_Valid_3_delay_20_16;
  reg                 io_A_Valid_3_delay_21_15;
  reg                 io_A_Valid_3_delay_22_14;
  reg                 io_A_Valid_3_delay_23_13;
  reg                 io_A_Valid_3_delay_24_12;
  reg                 io_A_Valid_3_delay_25_11;
  reg                 io_A_Valid_3_delay_26_10;
  reg                 io_A_Valid_3_delay_27_9;
  reg                 io_A_Valid_3_delay_28_8;
  reg                 io_A_Valid_3_delay_29_7;
  reg                 io_A_Valid_3_delay_30_6;
  reg                 io_A_Valid_3_delay_31_5;
  reg                 io_A_Valid_3_delay_32_4;
  reg                 io_A_Valid_3_delay_33_3;
  reg                 io_A_Valid_3_delay_34_2;
  reg                 io_A_Valid_3_delay_35_1;
  reg                 io_A_Valid_3_delay_36;
  reg                 io_B_Valid_36_delay_1_2;
  reg                 io_B_Valid_36_delay_2_1;
  reg                 io_B_Valid_36_delay_3;
  reg                 io_A_Valid_3_delay_1_36;
  reg                 io_A_Valid_3_delay_2_35;
  reg                 io_A_Valid_3_delay_3_34;
  reg                 io_A_Valid_3_delay_4_33;
  reg                 io_A_Valid_3_delay_5_32;
  reg                 io_A_Valid_3_delay_6_31;
  reg                 io_A_Valid_3_delay_7_30;
  reg                 io_A_Valid_3_delay_8_29;
  reg                 io_A_Valid_3_delay_9_28;
  reg                 io_A_Valid_3_delay_10_27;
  reg                 io_A_Valid_3_delay_11_26;
  reg                 io_A_Valid_3_delay_12_25;
  reg                 io_A_Valid_3_delay_13_24;
  reg                 io_A_Valid_3_delay_14_23;
  reg                 io_A_Valid_3_delay_15_22;
  reg                 io_A_Valid_3_delay_16_21;
  reg                 io_A_Valid_3_delay_17_20;
  reg                 io_A_Valid_3_delay_18_19;
  reg                 io_A_Valid_3_delay_19_18;
  reg                 io_A_Valid_3_delay_20_17;
  reg                 io_A_Valid_3_delay_21_16;
  reg                 io_A_Valid_3_delay_22_15;
  reg                 io_A_Valid_3_delay_23_14;
  reg                 io_A_Valid_3_delay_24_13;
  reg                 io_A_Valid_3_delay_25_12;
  reg                 io_A_Valid_3_delay_26_11;
  reg                 io_A_Valid_3_delay_27_10;
  reg                 io_A_Valid_3_delay_28_9;
  reg                 io_A_Valid_3_delay_29_8;
  reg                 io_A_Valid_3_delay_30_7;
  reg                 io_A_Valid_3_delay_31_6;
  reg                 io_A_Valid_3_delay_32_5;
  reg                 io_A_Valid_3_delay_33_4;
  reg                 io_A_Valid_3_delay_34_3;
  reg                 io_A_Valid_3_delay_35_2;
  reg                 io_A_Valid_3_delay_36_1;
  reg                 io_A_Valid_3_delay_37;
  reg                 io_B_Valid_37_delay_1_2;
  reg                 io_B_Valid_37_delay_2_1;
  reg                 io_B_Valid_37_delay_3;
  reg                 io_A_Valid_3_delay_1_37;
  reg                 io_A_Valid_3_delay_2_36;
  reg                 io_A_Valid_3_delay_3_35;
  reg                 io_A_Valid_3_delay_4_34;
  reg                 io_A_Valid_3_delay_5_33;
  reg                 io_A_Valid_3_delay_6_32;
  reg                 io_A_Valid_3_delay_7_31;
  reg                 io_A_Valid_3_delay_8_30;
  reg                 io_A_Valid_3_delay_9_29;
  reg                 io_A_Valid_3_delay_10_28;
  reg                 io_A_Valid_3_delay_11_27;
  reg                 io_A_Valid_3_delay_12_26;
  reg                 io_A_Valid_3_delay_13_25;
  reg                 io_A_Valid_3_delay_14_24;
  reg                 io_A_Valid_3_delay_15_23;
  reg                 io_A_Valid_3_delay_16_22;
  reg                 io_A_Valid_3_delay_17_21;
  reg                 io_A_Valid_3_delay_18_20;
  reg                 io_A_Valid_3_delay_19_19;
  reg                 io_A_Valid_3_delay_20_18;
  reg                 io_A_Valid_3_delay_21_17;
  reg                 io_A_Valid_3_delay_22_16;
  reg                 io_A_Valid_3_delay_23_15;
  reg                 io_A_Valid_3_delay_24_14;
  reg                 io_A_Valid_3_delay_25_13;
  reg                 io_A_Valid_3_delay_26_12;
  reg                 io_A_Valid_3_delay_27_11;
  reg                 io_A_Valid_3_delay_28_10;
  reg                 io_A_Valid_3_delay_29_9;
  reg                 io_A_Valid_3_delay_30_8;
  reg                 io_A_Valid_3_delay_31_7;
  reg                 io_A_Valid_3_delay_32_6;
  reg                 io_A_Valid_3_delay_33_5;
  reg                 io_A_Valid_3_delay_34_4;
  reg                 io_A_Valid_3_delay_35_3;
  reg                 io_A_Valid_3_delay_36_2;
  reg                 io_A_Valid_3_delay_37_1;
  reg                 io_A_Valid_3_delay_38;
  reg                 io_B_Valid_38_delay_1_2;
  reg                 io_B_Valid_38_delay_2_1;
  reg                 io_B_Valid_38_delay_3;
  reg                 io_A_Valid_3_delay_1_38;
  reg                 io_A_Valid_3_delay_2_37;
  reg                 io_A_Valid_3_delay_3_36;
  reg                 io_A_Valid_3_delay_4_35;
  reg                 io_A_Valid_3_delay_5_34;
  reg                 io_A_Valid_3_delay_6_33;
  reg                 io_A_Valid_3_delay_7_32;
  reg                 io_A_Valid_3_delay_8_31;
  reg                 io_A_Valid_3_delay_9_30;
  reg                 io_A_Valid_3_delay_10_29;
  reg                 io_A_Valid_3_delay_11_28;
  reg                 io_A_Valid_3_delay_12_27;
  reg                 io_A_Valid_3_delay_13_26;
  reg                 io_A_Valid_3_delay_14_25;
  reg                 io_A_Valid_3_delay_15_24;
  reg                 io_A_Valid_3_delay_16_23;
  reg                 io_A_Valid_3_delay_17_22;
  reg                 io_A_Valid_3_delay_18_21;
  reg                 io_A_Valid_3_delay_19_20;
  reg                 io_A_Valid_3_delay_20_19;
  reg                 io_A_Valid_3_delay_21_18;
  reg                 io_A_Valid_3_delay_22_17;
  reg                 io_A_Valid_3_delay_23_16;
  reg                 io_A_Valid_3_delay_24_15;
  reg                 io_A_Valid_3_delay_25_14;
  reg                 io_A_Valid_3_delay_26_13;
  reg                 io_A_Valid_3_delay_27_12;
  reg                 io_A_Valid_3_delay_28_11;
  reg                 io_A_Valid_3_delay_29_10;
  reg                 io_A_Valid_3_delay_30_9;
  reg                 io_A_Valid_3_delay_31_8;
  reg                 io_A_Valid_3_delay_32_7;
  reg                 io_A_Valid_3_delay_33_6;
  reg                 io_A_Valid_3_delay_34_5;
  reg                 io_A_Valid_3_delay_35_4;
  reg                 io_A_Valid_3_delay_36_3;
  reg                 io_A_Valid_3_delay_37_2;
  reg                 io_A_Valid_3_delay_38_1;
  reg                 io_A_Valid_3_delay_39;
  reg                 io_B_Valid_39_delay_1_2;
  reg                 io_B_Valid_39_delay_2_1;
  reg                 io_B_Valid_39_delay_3;
  reg                 io_A_Valid_3_delay_1_39;
  reg                 io_A_Valid_3_delay_2_38;
  reg                 io_A_Valid_3_delay_3_37;
  reg                 io_A_Valid_3_delay_4_36;
  reg                 io_A_Valid_3_delay_5_35;
  reg                 io_A_Valid_3_delay_6_34;
  reg                 io_A_Valid_3_delay_7_33;
  reg                 io_A_Valid_3_delay_8_32;
  reg                 io_A_Valid_3_delay_9_31;
  reg                 io_A_Valid_3_delay_10_30;
  reg                 io_A_Valid_3_delay_11_29;
  reg                 io_A_Valid_3_delay_12_28;
  reg                 io_A_Valid_3_delay_13_27;
  reg                 io_A_Valid_3_delay_14_26;
  reg                 io_A_Valid_3_delay_15_25;
  reg                 io_A_Valid_3_delay_16_24;
  reg                 io_A_Valid_3_delay_17_23;
  reg                 io_A_Valid_3_delay_18_22;
  reg                 io_A_Valid_3_delay_19_21;
  reg                 io_A_Valid_3_delay_20_20;
  reg                 io_A_Valid_3_delay_21_19;
  reg                 io_A_Valid_3_delay_22_18;
  reg                 io_A_Valid_3_delay_23_17;
  reg                 io_A_Valid_3_delay_24_16;
  reg                 io_A_Valid_3_delay_25_15;
  reg                 io_A_Valid_3_delay_26_14;
  reg                 io_A_Valid_3_delay_27_13;
  reg                 io_A_Valid_3_delay_28_12;
  reg                 io_A_Valid_3_delay_29_11;
  reg                 io_A_Valid_3_delay_30_10;
  reg                 io_A_Valid_3_delay_31_9;
  reg                 io_A_Valid_3_delay_32_8;
  reg                 io_A_Valid_3_delay_33_7;
  reg                 io_A_Valid_3_delay_34_6;
  reg                 io_A_Valid_3_delay_35_5;
  reg                 io_A_Valid_3_delay_36_4;
  reg                 io_A_Valid_3_delay_37_3;
  reg                 io_A_Valid_3_delay_38_2;
  reg                 io_A_Valid_3_delay_39_1;
  reg                 io_A_Valid_3_delay_40;
  reg                 io_B_Valid_40_delay_1_2;
  reg                 io_B_Valid_40_delay_2_1;
  reg                 io_B_Valid_40_delay_3;
  reg                 io_A_Valid_3_delay_1_40;
  reg                 io_A_Valid_3_delay_2_39;
  reg                 io_A_Valid_3_delay_3_38;
  reg                 io_A_Valid_3_delay_4_37;
  reg                 io_A_Valid_3_delay_5_36;
  reg                 io_A_Valid_3_delay_6_35;
  reg                 io_A_Valid_3_delay_7_34;
  reg                 io_A_Valid_3_delay_8_33;
  reg                 io_A_Valid_3_delay_9_32;
  reg                 io_A_Valid_3_delay_10_31;
  reg                 io_A_Valid_3_delay_11_30;
  reg                 io_A_Valid_3_delay_12_29;
  reg                 io_A_Valid_3_delay_13_28;
  reg                 io_A_Valid_3_delay_14_27;
  reg                 io_A_Valid_3_delay_15_26;
  reg                 io_A_Valid_3_delay_16_25;
  reg                 io_A_Valid_3_delay_17_24;
  reg                 io_A_Valid_3_delay_18_23;
  reg                 io_A_Valid_3_delay_19_22;
  reg                 io_A_Valid_3_delay_20_21;
  reg                 io_A_Valid_3_delay_21_20;
  reg                 io_A_Valid_3_delay_22_19;
  reg                 io_A_Valid_3_delay_23_18;
  reg                 io_A_Valid_3_delay_24_17;
  reg                 io_A_Valid_3_delay_25_16;
  reg                 io_A_Valid_3_delay_26_15;
  reg                 io_A_Valid_3_delay_27_14;
  reg                 io_A_Valid_3_delay_28_13;
  reg                 io_A_Valid_3_delay_29_12;
  reg                 io_A_Valid_3_delay_30_11;
  reg                 io_A_Valid_3_delay_31_10;
  reg                 io_A_Valid_3_delay_32_9;
  reg                 io_A_Valid_3_delay_33_8;
  reg                 io_A_Valid_3_delay_34_7;
  reg                 io_A_Valid_3_delay_35_6;
  reg                 io_A_Valid_3_delay_36_5;
  reg                 io_A_Valid_3_delay_37_4;
  reg                 io_A_Valid_3_delay_38_3;
  reg                 io_A_Valid_3_delay_39_2;
  reg                 io_A_Valid_3_delay_40_1;
  reg                 io_A_Valid_3_delay_41;
  reg                 io_B_Valid_41_delay_1_2;
  reg                 io_B_Valid_41_delay_2_1;
  reg                 io_B_Valid_41_delay_3;
  reg                 io_A_Valid_3_delay_1_41;
  reg                 io_A_Valid_3_delay_2_40;
  reg                 io_A_Valid_3_delay_3_39;
  reg                 io_A_Valid_3_delay_4_38;
  reg                 io_A_Valid_3_delay_5_37;
  reg                 io_A_Valid_3_delay_6_36;
  reg                 io_A_Valid_3_delay_7_35;
  reg                 io_A_Valid_3_delay_8_34;
  reg                 io_A_Valid_3_delay_9_33;
  reg                 io_A_Valid_3_delay_10_32;
  reg                 io_A_Valid_3_delay_11_31;
  reg                 io_A_Valid_3_delay_12_30;
  reg                 io_A_Valid_3_delay_13_29;
  reg                 io_A_Valid_3_delay_14_28;
  reg                 io_A_Valid_3_delay_15_27;
  reg                 io_A_Valid_3_delay_16_26;
  reg                 io_A_Valid_3_delay_17_25;
  reg                 io_A_Valid_3_delay_18_24;
  reg                 io_A_Valid_3_delay_19_23;
  reg                 io_A_Valid_3_delay_20_22;
  reg                 io_A_Valid_3_delay_21_21;
  reg                 io_A_Valid_3_delay_22_20;
  reg                 io_A_Valid_3_delay_23_19;
  reg                 io_A_Valid_3_delay_24_18;
  reg                 io_A_Valid_3_delay_25_17;
  reg                 io_A_Valid_3_delay_26_16;
  reg                 io_A_Valid_3_delay_27_15;
  reg                 io_A_Valid_3_delay_28_14;
  reg                 io_A_Valid_3_delay_29_13;
  reg                 io_A_Valid_3_delay_30_12;
  reg                 io_A_Valid_3_delay_31_11;
  reg                 io_A_Valid_3_delay_32_10;
  reg                 io_A_Valid_3_delay_33_9;
  reg                 io_A_Valid_3_delay_34_8;
  reg                 io_A_Valid_3_delay_35_7;
  reg                 io_A_Valid_3_delay_36_6;
  reg                 io_A_Valid_3_delay_37_5;
  reg                 io_A_Valid_3_delay_38_4;
  reg                 io_A_Valid_3_delay_39_3;
  reg                 io_A_Valid_3_delay_40_2;
  reg                 io_A_Valid_3_delay_41_1;
  reg                 io_A_Valid_3_delay_42;
  reg                 io_B_Valid_42_delay_1_2;
  reg                 io_B_Valid_42_delay_2_1;
  reg                 io_B_Valid_42_delay_3;
  reg                 io_A_Valid_3_delay_1_42;
  reg                 io_A_Valid_3_delay_2_41;
  reg                 io_A_Valid_3_delay_3_40;
  reg                 io_A_Valid_3_delay_4_39;
  reg                 io_A_Valid_3_delay_5_38;
  reg                 io_A_Valid_3_delay_6_37;
  reg                 io_A_Valid_3_delay_7_36;
  reg                 io_A_Valid_3_delay_8_35;
  reg                 io_A_Valid_3_delay_9_34;
  reg                 io_A_Valid_3_delay_10_33;
  reg                 io_A_Valid_3_delay_11_32;
  reg                 io_A_Valid_3_delay_12_31;
  reg                 io_A_Valid_3_delay_13_30;
  reg                 io_A_Valid_3_delay_14_29;
  reg                 io_A_Valid_3_delay_15_28;
  reg                 io_A_Valid_3_delay_16_27;
  reg                 io_A_Valid_3_delay_17_26;
  reg                 io_A_Valid_3_delay_18_25;
  reg                 io_A_Valid_3_delay_19_24;
  reg                 io_A_Valid_3_delay_20_23;
  reg                 io_A_Valid_3_delay_21_22;
  reg                 io_A_Valid_3_delay_22_21;
  reg                 io_A_Valid_3_delay_23_20;
  reg                 io_A_Valid_3_delay_24_19;
  reg                 io_A_Valid_3_delay_25_18;
  reg                 io_A_Valid_3_delay_26_17;
  reg                 io_A_Valid_3_delay_27_16;
  reg                 io_A_Valid_3_delay_28_15;
  reg                 io_A_Valid_3_delay_29_14;
  reg                 io_A_Valid_3_delay_30_13;
  reg                 io_A_Valid_3_delay_31_12;
  reg                 io_A_Valid_3_delay_32_11;
  reg                 io_A_Valid_3_delay_33_10;
  reg                 io_A_Valid_3_delay_34_9;
  reg                 io_A_Valid_3_delay_35_8;
  reg                 io_A_Valid_3_delay_36_7;
  reg                 io_A_Valid_3_delay_37_6;
  reg                 io_A_Valid_3_delay_38_5;
  reg                 io_A_Valid_3_delay_39_4;
  reg                 io_A_Valid_3_delay_40_3;
  reg                 io_A_Valid_3_delay_41_2;
  reg                 io_A_Valid_3_delay_42_1;
  reg                 io_A_Valid_3_delay_43;
  reg                 io_B_Valid_43_delay_1_2;
  reg                 io_B_Valid_43_delay_2_1;
  reg                 io_B_Valid_43_delay_3;
  reg                 io_A_Valid_3_delay_1_43;
  reg                 io_A_Valid_3_delay_2_42;
  reg                 io_A_Valid_3_delay_3_41;
  reg                 io_A_Valid_3_delay_4_40;
  reg                 io_A_Valid_3_delay_5_39;
  reg                 io_A_Valid_3_delay_6_38;
  reg                 io_A_Valid_3_delay_7_37;
  reg                 io_A_Valid_3_delay_8_36;
  reg                 io_A_Valid_3_delay_9_35;
  reg                 io_A_Valid_3_delay_10_34;
  reg                 io_A_Valid_3_delay_11_33;
  reg                 io_A_Valid_3_delay_12_32;
  reg                 io_A_Valid_3_delay_13_31;
  reg                 io_A_Valid_3_delay_14_30;
  reg                 io_A_Valid_3_delay_15_29;
  reg                 io_A_Valid_3_delay_16_28;
  reg                 io_A_Valid_3_delay_17_27;
  reg                 io_A_Valid_3_delay_18_26;
  reg                 io_A_Valid_3_delay_19_25;
  reg                 io_A_Valid_3_delay_20_24;
  reg                 io_A_Valid_3_delay_21_23;
  reg                 io_A_Valid_3_delay_22_22;
  reg                 io_A_Valid_3_delay_23_21;
  reg                 io_A_Valid_3_delay_24_20;
  reg                 io_A_Valid_3_delay_25_19;
  reg                 io_A_Valid_3_delay_26_18;
  reg                 io_A_Valid_3_delay_27_17;
  reg                 io_A_Valid_3_delay_28_16;
  reg                 io_A_Valid_3_delay_29_15;
  reg                 io_A_Valid_3_delay_30_14;
  reg                 io_A_Valid_3_delay_31_13;
  reg                 io_A_Valid_3_delay_32_12;
  reg                 io_A_Valid_3_delay_33_11;
  reg                 io_A_Valid_3_delay_34_10;
  reg                 io_A_Valid_3_delay_35_9;
  reg                 io_A_Valid_3_delay_36_8;
  reg                 io_A_Valid_3_delay_37_7;
  reg                 io_A_Valid_3_delay_38_6;
  reg                 io_A_Valid_3_delay_39_5;
  reg                 io_A_Valid_3_delay_40_4;
  reg                 io_A_Valid_3_delay_41_3;
  reg                 io_A_Valid_3_delay_42_2;
  reg                 io_A_Valid_3_delay_43_1;
  reg                 io_A_Valid_3_delay_44;
  reg                 io_B_Valid_44_delay_1_2;
  reg                 io_B_Valid_44_delay_2_1;
  reg                 io_B_Valid_44_delay_3;
  reg                 io_A_Valid_3_delay_1_44;
  reg                 io_A_Valid_3_delay_2_43;
  reg                 io_A_Valid_3_delay_3_42;
  reg                 io_A_Valid_3_delay_4_41;
  reg                 io_A_Valid_3_delay_5_40;
  reg                 io_A_Valid_3_delay_6_39;
  reg                 io_A_Valid_3_delay_7_38;
  reg                 io_A_Valid_3_delay_8_37;
  reg                 io_A_Valid_3_delay_9_36;
  reg                 io_A_Valid_3_delay_10_35;
  reg                 io_A_Valid_3_delay_11_34;
  reg                 io_A_Valid_3_delay_12_33;
  reg                 io_A_Valid_3_delay_13_32;
  reg                 io_A_Valid_3_delay_14_31;
  reg                 io_A_Valid_3_delay_15_30;
  reg                 io_A_Valid_3_delay_16_29;
  reg                 io_A_Valid_3_delay_17_28;
  reg                 io_A_Valid_3_delay_18_27;
  reg                 io_A_Valid_3_delay_19_26;
  reg                 io_A_Valid_3_delay_20_25;
  reg                 io_A_Valid_3_delay_21_24;
  reg                 io_A_Valid_3_delay_22_23;
  reg                 io_A_Valid_3_delay_23_22;
  reg                 io_A_Valid_3_delay_24_21;
  reg                 io_A_Valid_3_delay_25_20;
  reg                 io_A_Valid_3_delay_26_19;
  reg                 io_A_Valid_3_delay_27_18;
  reg                 io_A_Valid_3_delay_28_17;
  reg                 io_A_Valid_3_delay_29_16;
  reg                 io_A_Valid_3_delay_30_15;
  reg                 io_A_Valid_3_delay_31_14;
  reg                 io_A_Valid_3_delay_32_13;
  reg                 io_A_Valid_3_delay_33_12;
  reg                 io_A_Valid_3_delay_34_11;
  reg                 io_A_Valid_3_delay_35_10;
  reg                 io_A_Valid_3_delay_36_9;
  reg                 io_A_Valid_3_delay_37_8;
  reg                 io_A_Valid_3_delay_38_7;
  reg                 io_A_Valid_3_delay_39_6;
  reg                 io_A_Valid_3_delay_40_5;
  reg                 io_A_Valid_3_delay_41_4;
  reg                 io_A_Valid_3_delay_42_3;
  reg                 io_A_Valid_3_delay_43_2;
  reg                 io_A_Valid_3_delay_44_1;
  reg                 io_A_Valid_3_delay_45;
  reg                 io_B_Valid_45_delay_1_2;
  reg                 io_B_Valid_45_delay_2_1;
  reg                 io_B_Valid_45_delay_3;
  reg                 io_A_Valid_3_delay_1_45;
  reg                 io_A_Valid_3_delay_2_44;
  reg                 io_A_Valid_3_delay_3_43;
  reg                 io_A_Valid_3_delay_4_42;
  reg                 io_A_Valid_3_delay_5_41;
  reg                 io_A_Valid_3_delay_6_40;
  reg                 io_A_Valid_3_delay_7_39;
  reg                 io_A_Valid_3_delay_8_38;
  reg                 io_A_Valid_3_delay_9_37;
  reg                 io_A_Valid_3_delay_10_36;
  reg                 io_A_Valid_3_delay_11_35;
  reg                 io_A_Valid_3_delay_12_34;
  reg                 io_A_Valid_3_delay_13_33;
  reg                 io_A_Valid_3_delay_14_32;
  reg                 io_A_Valid_3_delay_15_31;
  reg                 io_A_Valid_3_delay_16_30;
  reg                 io_A_Valid_3_delay_17_29;
  reg                 io_A_Valid_3_delay_18_28;
  reg                 io_A_Valid_3_delay_19_27;
  reg                 io_A_Valid_3_delay_20_26;
  reg                 io_A_Valid_3_delay_21_25;
  reg                 io_A_Valid_3_delay_22_24;
  reg                 io_A_Valid_3_delay_23_23;
  reg                 io_A_Valid_3_delay_24_22;
  reg                 io_A_Valid_3_delay_25_21;
  reg                 io_A_Valid_3_delay_26_20;
  reg                 io_A_Valid_3_delay_27_19;
  reg                 io_A_Valid_3_delay_28_18;
  reg                 io_A_Valid_3_delay_29_17;
  reg                 io_A_Valid_3_delay_30_16;
  reg                 io_A_Valid_3_delay_31_15;
  reg                 io_A_Valid_3_delay_32_14;
  reg                 io_A_Valid_3_delay_33_13;
  reg                 io_A_Valid_3_delay_34_12;
  reg                 io_A_Valid_3_delay_35_11;
  reg                 io_A_Valid_3_delay_36_10;
  reg                 io_A_Valid_3_delay_37_9;
  reg                 io_A_Valid_3_delay_38_8;
  reg                 io_A_Valid_3_delay_39_7;
  reg                 io_A_Valid_3_delay_40_6;
  reg                 io_A_Valid_3_delay_41_5;
  reg                 io_A_Valid_3_delay_42_4;
  reg                 io_A_Valid_3_delay_43_3;
  reg                 io_A_Valid_3_delay_44_2;
  reg                 io_A_Valid_3_delay_45_1;
  reg                 io_A_Valid_3_delay_46;
  reg                 io_B_Valid_46_delay_1_2;
  reg                 io_B_Valid_46_delay_2_1;
  reg                 io_B_Valid_46_delay_3;
  reg                 io_A_Valid_3_delay_1_46;
  reg                 io_A_Valid_3_delay_2_45;
  reg                 io_A_Valid_3_delay_3_44;
  reg                 io_A_Valid_3_delay_4_43;
  reg                 io_A_Valid_3_delay_5_42;
  reg                 io_A_Valid_3_delay_6_41;
  reg                 io_A_Valid_3_delay_7_40;
  reg                 io_A_Valid_3_delay_8_39;
  reg                 io_A_Valid_3_delay_9_38;
  reg                 io_A_Valid_3_delay_10_37;
  reg                 io_A_Valid_3_delay_11_36;
  reg                 io_A_Valid_3_delay_12_35;
  reg                 io_A_Valid_3_delay_13_34;
  reg                 io_A_Valid_3_delay_14_33;
  reg                 io_A_Valid_3_delay_15_32;
  reg                 io_A_Valid_3_delay_16_31;
  reg                 io_A_Valid_3_delay_17_30;
  reg                 io_A_Valid_3_delay_18_29;
  reg                 io_A_Valid_3_delay_19_28;
  reg                 io_A_Valid_3_delay_20_27;
  reg                 io_A_Valid_3_delay_21_26;
  reg                 io_A_Valid_3_delay_22_25;
  reg                 io_A_Valid_3_delay_23_24;
  reg                 io_A_Valid_3_delay_24_23;
  reg                 io_A_Valid_3_delay_25_22;
  reg                 io_A_Valid_3_delay_26_21;
  reg                 io_A_Valid_3_delay_27_20;
  reg                 io_A_Valid_3_delay_28_19;
  reg                 io_A_Valid_3_delay_29_18;
  reg                 io_A_Valid_3_delay_30_17;
  reg                 io_A_Valid_3_delay_31_16;
  reg                 io_A_Valid_3_delay_32_15;
  reg                 io_A_Valid_3_delay_33_14;
  reg                 io_A_Valid_3_delay_34_13;
  reg                 io_A_Valid_3_delay_35_12;
  reg                 io_A_Valid_3_delay_36_11;
  reg                 io_A_Valid_3_delay_37_10;
  reg                 io_A_Valid_3_delay_38_9;
  reg                 io_A_Valid_3_delay_39_8;
  reg                 io_A_Valid_3_delay_40_7;
  reg                 io_A_Valid_3_delay_41_6;
  reg                 io_A_Valid_3_delay_42_5;
  reg                 io_A_Valid_3_delay_43_4;
  reg                 io_A_Valid_3_delay_44_3;
  reg                 io_A_Valid_3_delay_45_2;
  reg                 io_A_Valid_3_delay_46_1;
  reg                 io_A_Valid_3_delay_47;
  reg                 io_B_Valid_47_delay_1_2;
  reg                 io_B_Valid_47_delay_2_1;
  reg                 io_B_Valid_47_delay_3;
  reg                 io_A_Valid_3_delay_1_47;
  reg                 io_A_Valid_3_delay_2_46;
  reg                 io_A_Valid_3_delay_3_45;
  reg                 io_A_Valid_3_delay_4_44;
  reg                 io_A_Valid_3_delay_5_43;
  reg                 io_A_Valid_3_delay_6_42;
  reg                 io_A_Valid_3_delay_7_41;
  reg                 io_A_Valid_3_delay_8_40;
  reg                 io_A_Valid_3_delay_9_39;
  reg                 io_A_Valid_3_delay_10_38;
  reg                 io_A_Valid_3_delay_11_37;
  reg                 io_A_Valid_3_delay_12_36;
  reg                 io_A_Valid_3_delay_13_35;
  reg                 io_A_Valid_3_delay_14_34;
  reg                 io_A_Valid_3_delay_15_33;
  reg                 io_A_Valid_3_delay_16_32;
  reg                 io_A_Valid_3_delay_17_31;
  reg                 io_A_Valid_3_delay_18_30;
  reg                 io_A_Valid_3_delay_19_29;
  reg                 io_A_Valid_3_delay_20_28;
  reg                 io_A_Valid_3_delay_21_27;
  reg                 io_A_Valid_3_delay_22_26;
  reg                 io_A_Valid_3_delay_23_25;
  reg                 io_A_Valid_3_delay_24_24;
  reg                 io_A_Valid_3_delay_25_23;
  reg                 io_A_Valid_3_delay_26_22;
  reg                 io_A_Valid_3_delay_27_21;
  reg                 io_A_Valid_3_delay_28_20;
  reg                 io_A_Valid_3_delay_29_19;
  reg                 io_A_Valid_3_delay_30_18;
  reg                 io_A_Valid_3_delay_31_17;
  reg                 io_A_Valid_3_delay_32_16;
  reg                 io_A_Valid_3_delay_33_15;
  reg                 io_A_Valid_3_delay_34_14;
  reg                 io_A_Valid_3_delay_35_13;
  reg                 io_A_Valid_3_delay_36_12;
  reg                 io_A_Valid_3_delay_37_11;
  reg                 io_A_Valid_3_delay_38_10;
  reg                 io_A_Valid_3_delay_39_9;
  reg                 io_A_Valid_3_delay_40_8;
  reg                 io_A_Valid_3_delay_41_7;
  reg                 io_A_Valid_3_delay_42_6;
  reg                 io_A_Valid_3_delay_43_5;
  reg                 io_A_Valid_3_delay_44_4;
  reg                 io_A_Valid_3_delay_45_3;
  reg                 io_A_Valid_3_delay_46_2;
  reg                 io_A_Valid_3_delay_47_1;
  reg                 io_A_Valid_3_delay_48;
  reg                 io_B_Valid_48_delay_1_2;
  reg                 io_B_Valid_48_delay_2_1;
  reg                 io_B_Valid_48_delay_3;
  reg                 io_A_Valid_3_delay_1_48;
  reg                 io_A_Valid_3_delay_2_47;
  reg                 io_A_Valid_3_delay_3_46;
  reg                 io_A_Valid_3_delay_4_45;
  reg                 io_A_Valid_3_delay_5_44;
  reg                 io_A_Valid_3_delay_6_43;
  reg                 io_A_Valid_3_delay_7_42;
  reg                 io_A_Valid_3_delay_8_41;
  reg                 io_A_Valid_3_delay_9_40;
  reg                 io_A_Valid_3_delay_10_39;
  reg                 io_A_Valid_3_delay_11_38;
  reg                 io_A_Valid_3_delay_12_37;
  reg                 io_A_Valid_3_delay_13_36;
  reg                 io_A_Valid_3_delay_14_35;
  reg                 io_A_Valid_3_delay_15_34;
  reg                 io_A_Valid_3_delay_16_33;
  reg                 io_A_Valid_3_delay_17_32;
  reg                 io_A_Valid_3_delay_18_31;
  reg                 io_A_Valid_3_delay_19_30;
  reg                 io_A_Valid_3_delay_20_29;
  reg                 io_A_Valid_3_delay_21_28;
  reg                 io_A_Valid_3_delay_22_27;
  reg                 io_A_Valid_3_delay_23_26;
  reg                 io_A_Valid_3_delay_24_25;
  reg                 io_A_Valid_3_delay_25_24;
  reg                 io_A_Valid_3_delay_26_23;
  reg                 io_A_Valid_3_delay_27_22;
  reg                 io_A_Valid_3_delay_28_21;
  reg                 io_A_Valid_3_delay_29_20;
  reg                 io_A_Valid_3_delay_30_19;
  reg                 io_A_Valid_3_delay_31_18;
  reg                 io_A_Valid_3_delay_32_17;
  reg                 io_A_Valid_3_delay_33_16;
  reg                 io_A_Valid_3_delay_34_15;
  reg                 io_A_Valid_3_delay_35_14;
  reg                 io_A_Valid_3_delay_36_13;
  reg                 io_A_Valid_3_delay_37_12;
  reg                 io_A_Valid_3_delay_38_11;
  reg                 io_A_Valid_3_delay_39_10;
  reg                 io_A_Valid_3_delay_40_9;
  reg                 io_A_Valid_3_delay_41_8;
  reg                 io_A_Valid_3_delay_42_7;
  reg                 io_A_Valid_3_delay_43_6;
  reg                 io_A_Valid_3_delay_44_5;
  reg                 io_A_Valid_3_delay_45_4;
  reg                 io_A_Valid_3_delay_46_3;
  reg                 io_A_Valid_3_delay_47_2;
  reg                 io_A_Valid_3_delay_48_1;
  reg                 io_A_Valid_3_delay_49;
  reg                 io_B_Valid_49_delay_1_2;
  reg                 io_B_Valid_49_delay_2_1;
  reg                 io_B_Valid_49_delay_3;
  reg                 io_A_Valid_3_delay_1_49;
  reg                 io_A_Valid_3_delay_2_48;
  reg                 io_A_Valid_3_delay_3_47;
  reg                 io_A_Valid_3_delay_4_46;
  reg                 io_A_Valid_3_delay_5_45;
  reg                 io_A_Valid_3_delay_6_44;
  reg                 io_A_Valid_3_delay_7_43;
  reg                 io_A_Valid_3_delay_8_42;
  reg                 io_A_Valid_3_delay_9_41;
  reg                 io_A_Valid_3_delay_10_40;
  reg                 io_A_Valid_3_delay_11_39;
  reg                 io_A_Valid_3_delay_12_38;
  reg                 io_A_Valid_3_delay_13_37;
  reg                 io_A_Valid_3_delay_14_36;
  reg                 io_A_Valid_3_delay_15_35;
  reg                 io_A_Valid_3_delay_16_34;
  reg                 io_A_Valid_3_delay_17_33;
  reg                 io_A_Valid_3_delay_18_32;
  reg                 io_A_Valid_3_delay_19_31;
  reg                 io_A_Valid_3_delay_20_30;
  reg                 io_A_Valid_3_delay_21_29;
  reg                 io_A_Valid_3_delay_22_28;
  reg                 io_A_Valid_3_delay_23_27;
  reg                 io_A_Valid_3_delay_24_26;
  reg                 io_A_Valid_3_delay_25_25;
  reg                 io_A_Valid_3_delay_26_24;
  reg                 io_A_Valid_3_delay_27_23;
  reg                 io_A_Valid_3_delay_28_22;
  reg                 io_A_Valid_3_delay_29_21;
  reg                 io_A_Valid_3_delay_30_20;
  reg                 io_A_Valid_3_delay_31_19;
  reg                 io_A_Valid_3_delay_32_18;
  reg                 io_A_Valid_3_delay_33_17;
  reg                 io_A_Valid_3_delay_34_16;
  reg                 io_A_Valid_3_delay_35_15;
  reg                 io_A_Valid_3_delay_36_14;
  reg                 io_A_Valid_3_delay_37_13;
  reg                 io_A_Valid_3_delay_38_12;
  reg                 io_A_Valid_3_delay_39_11;
  reg                 io_A_Valid_3_delay_40_10;
  reg                 io_A_Valid_3_delay_41_9;
  reg                 io_A_Valid_3_delay_42_8;
  reg                 io_A_Valid_3_delay_43_7;
  reg                 io_A_Valid_3_delay_44_6;
  reg                 io_A_Valid_3_delay_45_5;
  reg                 io_A_Valid_3_delay_46_4;
  reg                 io_A_Valid_3_delay_47_3;
  reg                 io_A_Valid_3_delay_48_2;
  reg                 io_A_Valid_3_delay_49_1;
  reg                 io_A_Valid_3_delay_50;
  reg                 io_B_Valid_50_delay_1_2;
  reg                 io_B_Valid_50_delay_2_1;
  reg                 io_B_Valid_50_delay_3;
  reg                 io_A_Valid_3_delay_1_50;
  reg                 io_A_Valid_3_delay_2_49;
  reg                 io_A_Valid_3_delay_3_48;
  reg                 io_A_Valid_3_delay_4_47;
  reg                 io_A_Valid_3_delay_5_46;
  reg                 io_A_Valid_3_delay_6_45;
  reg                 io_A_Valid_3_delay_7_44;
  reg                 io_A_Valid_3_delay_8_43;
  reg                 io_A_Valid_3_delay_9_42;
  reg                 io_A_Valid_3_delay_10_41;
  reg                 io_A_Valid_3_delay_11_40;
  reg                 io_A_Valid_3_delay_12_39;
  reg                 io_A_Valid_3_delay_13_38;
  reg                 io_A_Valid_3_delay_14_37;
  reg                 io_A_Valid_3_delay_15_36;
  reg                 io_A_Valid_3_delay_16_35;
  reg                 io_A_Valid_3_delay_17_34;
  reg                 io_A_Valid_3_delay_18_33;
  reg                 io_A_Valid_3_delay_19_32;
  reg                 io_A_Valid_3_delay_20_31;
  reg                 io_A_Valid_3_delay_21_30;
  reg                 io_A_Valid_3_delay_22_29;
  reg                 io_A_Valid_3_delay_23_28;
  reg                 io_A_Valid_3_delay_24_27;
  reg                 io_A_Valid_3_delay_25_26;
  reg                 io_A_Valid_3_delay_26_25;
  reg                 io_A_Valid_3_delay_27_24;
  reg                 io_A_Valid_3_delay_28_23;
  reg                 io_A_Valid_3_delay_29_22;
  reg                 io_A_Valid_3_delay_30_21;
  reg                 io_A_Valid_3_delay_31_20;
  reg                 io_A_Valid_3_delay_32_19;
  reg                 io_A_Valid_3_delay_33_18;
  reg                 io_A_Valid_3_delay_34_17;
  reg                 io_A_Valid_3_delay_35_16;
  reg                 io_A_Valid_3_delay_36_15;
  reg                 io_A_Valid_3_delay_37_14;
  reg                 io_A_Valid_3_delay_38_13;
  reg                 io_A_Valid_3_delay_39_12;
  reg                 io_A_Valid_3_delay_40_11;
  reg                 io_A_Valid_3_delay_41_10;
  reg                 io_A_Valid_3_delay_42_9;
  reg                 io_A_Valid_3_delay_43_8;
  reg                 io_A_Valid_3_delay_44_7;
  reg                 io_A_Valid_3_delay_45_6;
  reg                 io_A_Valid_3_delay_46_5;
  reg                 io_A_Valid_3_delay_47_4;
  reg                 io_A_Valid_3_delay_48_3;
  reg                 io_A_Valid_3_delay_49_2;
  reg                 io_A_Valid_3_delay_50_1;
  reg                 io_A_Valid_3_delay_51;
  reg                 io_B_Valid_51_delay_1_2;
  reg                 io_B_Valid_51_delay_2_1;
  reg                 io_B_Valid_51_delay_3;
  reg                 io_A_Valid_3_delay_1_51;
  reg                 io_A_Valid_3_delay_2_50;
  reg                 io_A_Valid_3_delay_3_49;
  reg                 io_A_Valid_3_delay_4_48;
  reg                 io_A_Valid_3_delay_5_47;
  reg                 io_A_Valid_3_delay_6_46;
  reg                 io_A_Valid_3_delay_7_45;
  reg                 io_A_Valid_3_delay_8_44;
  reg                 io_A_Valid_3_delay_9_43;
  reg                 io_A_Valid_3_delay_10_42;
  reg                 io_A_Valid_3_delay_11_41;
  reg                 io_A_Valid_3_delay_12_40;
  reg                 io_A_Valid_3_delay_13_39;
  reg                 io_A_Valid_3_delay_14_38;
  reg                 io_A_Valid_3_delay_15_37;
  reg                 io_A_Valid_3_delay_16_36;
  reg                 io_A_Valid_3_delay_17_35;
  reg                 io_A_Valid_3_delay_18_34;
  reg                 io_A_Valid_3_delay_19_33;
  reg                 io_A_Valid_3_delay_20_32;
  reg                 io_A_Valid_3_delay_21_31;
  reg                 io_A_Valid_3_delay_22_30;
  reg                 io_A_Valid_3_delay_23_29;
  reg                 io_A_Valid_3_delay_24_28;
  reg                 io_A_Valid_3_delay_25_27;
  reg                 io_A_Valid_3_delay_26_26;
  reg                 io_A_Valid_3_delay_27_25;
  reg                 io_A_Valid_3_delay_28_24;
  reg                 io_A_Valid_3_delay_29_23;
  reg                 io_A_Valid_3_delay_30_22;
  reg                 io_A_Valid_3_delay_31_21;
  reg                 io_A_Valid_3_delay_32_20;
  reg                 io_A_Valid_3_delay_33_19;
  reg                 io_A_Valid_3_delay_34_18;
  reg                 io_A_Valid_3_delay_35_17;
  reg                 io_A_Valid_3_delay_36_16;
  reg                 io_A_Valid_3_delay_37_15;
  reg                 io_A_Valid_3_delay_38_14;
  reg                 io_A_Valid_3_delay_39_13;
  reg                 io_A_Valid_3_delay_40_12;
  reg                 io_A_Valid_3_delay_41_11;
  reg                 io_A_Valid_3_delay_42_10;
  reg                 io_A_Valid_3_delay_43_9;
  reg                 io_A_Valid_3_delay_44_8;
  reg                 io_A_Valid_3_delay_45_7;
  reg                 io_A_Valid_3_delay_46_6;
  reg                 io_A_Valid_3_delay_47_5;
  reg                 io_A_Valid_3_delay_48_4;
  reg                 io_A_Valid_3_delay_49_3;
  reg                 io_A_Valid_3_delay_50_2;
  reg                 io_A_Valid_3_delay_51_1;
  reg                 io_A_Valid_3_delay_52;
  reg                 io_B_Valid_52_delay_1_2;
  reg                 io_B_Valid_52_delay_2_1;
  reg                 io_B_Valid_52_delay_3;
  reg                 io_A_Valid_3_delay_1_52;
  reg                 io_A_Valid_3_delay_2_51;
  reg                 io_A_Valid_3_delay_3_50;
  reg                 io_A_Valid_3_delay_4_49;
  reg                 io_A_Valid_3_delay_5_48;
  reg                 io_A_Valid_3_delay_6_47;
  reg                 io_A_Valid_3_delay_7_46;
  reg                 io_A_Valid_3_delay_8_45;
  reg                 io_A_Valid_3_delay_9_44;
  reg                 io_A_Valid_3_delay_10_43;
  reg                 io_A_Valid_3_delay_11_42;
  reg                 io_A_Valid_3_delay_12_41;
  reg                 io_A_Valid_3_delay_13_40;
  reg                 io_A_Valid_3_delay_14_39;
  reg                 io_A_Valid_3_delay_15_38;
  reg                 io_A_Valid_3_delay_16_37;
  reg                 io_A_Valid_3_delay_17_36;
  reg                 io_A_Valid_3_delay_18_35;
  reg                 io_A_Valid_3_delay_19_34;
  reg                 io_A_Valid_3_delay_20_33;
  reg                 io_A_Valid_3_delay_21_32;
  reg                 io_A_Valid_3_delay_22_31;
  reg                 io_A_Valid_3_delay_23_30;
  reg                 io_A_Valid_3_delay_24_29;
  reg                 io_A_Valid_3_delay_25_28;
  reg                 io_A_Valid_3_delay_26_27;
  reg                 io_A_Valid_3_delay_27_26;
  reg                 io_A_Valid_3_delay_28_25;
  reg                 io_A_Valid_3_delay_29_24;
  reg                 io_A_Valid_3_delay_30_23;
  reg                 io_A_Valid_3_delay_31_22;
  reg                 io_A_Valid_3_delay_32_21;
  reg                 io_A_Valid_3_delay_33_20;
  reg                 io_A_Valid_3_delay_34_19;
  reg                 io_A_Valid_3_delay_35_18;
  reg                 io_A_Valid_3_delay_36_17;
  reg                 io_A_Valid_3_delay_37_16;
  reg                 io_A_Valid_3_delay_38_15;
  reg                 io_A_Valid_3_delay_39_14;
  reg                 io_A_Valid_3_delay_40_13;
  reg                 io_A_Valid_3_delay_41_12;
  reg                 io_A_Valid_3_delay_42_11;
  reg                 io_A_Valid_3_delay_43_10;
  reg                 io_A_Valid_3_delay_44_9;
  reg                 io_A_Valid_3_delay_45_8;
  reg                 io_A_Valid_3_delay_46_7;
  reg                 io_A_Valid_3_delay_47_6;
  reg                 io_A_Valid_3_delay_48_5;
  reg                 io_A_Valid_3_delay_49_4;
  reg                 io_A_Valid_3_delay_50_3;
  reg                 io_A_Valid_3_delay_51_2;
  reg                 io_A_Valid_3_delay_52_1;
  reg                 io_A_Valid_3_delay_53;
  reg                 io_B_Valid_53_delay_1_2;
  reg                 io_B_Valid_53_delay_2_1;
  reg                 io_B_Valid_53_delay_3;
  reg                 io_A_Valid_3_delay_1_53;
  reg                 io_A_Valid_3_delay_2_52;
  reg                 io_A_Valid_3_delay_3_51;
  reg                 io_A_Valid_3_delay_4_50;
  reg                 io_A_Valid_3_delay_5_49;
  reg                 io_A_Valid_3_delay_6_48;
  reg                 io_A_Valid_3_delay_7_47;
  reg                 io_A_Valid_3_delay_8_46;
  reg                 io_A_Valid_3_delay_9_45;
  reg                 io_A_Valid_3_delay_10_44;
  reg                 io_A_Valid_3_delay_11_43;
  reg                 io_A_Valid_3_delay_12_42;
  reg                 io_A_Valid_3_delay_13_41;
  reg                 io_A_Valid_3_delay_14_40;
  reg                 io_A_Valid_3_delay_15_39;
  reg                 io_A_Valid_3_delay_16_38;
  reg                 io_A_Valid_3_delay_17_37;
  reg                 io_A_Valid_3_delay_18_36;
  reg                 io_A_Valid_3_delay_19_35;
  reg                 io_A_Valid_3_delay_20_34;
  reg                 io_A_Valid_3_delay_21_33;
  reg                 io_A_Valid_3_delay_22_32;
  reg                 io_A_Valid_3_delay_23_31;
  reg                 io_A_Valid_3_delay_24_30;
  reg                 io_A_Valid_3_delay_25_29;
  reg                 io_A_Valid_3_delay_26_28;
  reg                 io_A_Valid_3_delay_27_27;
  reg                 io_A_Valid_3_delay_28_26;
  reg                 io_A_Valid_3_delay_29_25;
  reg                 io_A_Valid_3_delay_30_24;
  reg                 io_A_Valid_3_delay_31_23;
  reg                 io_A_Valid_3_delay_32_22;
  reg                 io_A_Valid_3_delay_33_21;
  reg                 io_A_Valid_3_delay_34_20;
  reg                 io_A_Valid_3_delay_35_19;
  reg                 io_A_Valid_3_delay_36_18;
  reg                 io_A_Valid_3_delay_37_17;
  reg                 io_A_Valid_3_delay_38_16;
  reg                 io_A_Valid_3_delay_39_15;
  reg                 io_A_Valid_3_delay_40_14;
  reg                 io_A_Valid_3_delay_41_13;
  reg                 io_A_Valid_3_delay_42_12;
  reg                 io_A_Valid_3_delay_43_11;
  reg                 io_A_Valid_3_delay_44_10;
  reg                 io_A_Valid_3_delay_45_9;
  reg                 io_A_Valid_3_delay_46_8;
  reg                 io_A_Valid_3_delay_47_7;
  reg                 io_A_Valid_3_delay_48_6;
  reg                 io_A_Valid_3_delay_49_5;
  reg                 io_A_Valid_3_delay_50_4;
  reg                 io_A_Valid_3_delay_51_3;
  reg                 io_A_Valid_3_delay_52_2;
  reg                 io_A_Valid_3_delay_53_1;
  reg                 io_A_Valid_3_delay_54;
  reg                 io_B_Valid_54_delay_1_2;
  reg                 io_B_Valid_54_delay_2_1;
  reg                 io_B_Valid_54_delay_3;
  reg                 io_A_Valid_3_delay_1_54;
  reg                 io_A_Valid_3_delay_2_53;
  reg                 io_A_Valid_3_delay_3_52;
  reg                 io_A_Valid_3_delay_4_51;
  reg                 io_A_Valid_3_delay_5_50;
  reg                 io_A_Valid_3_delay_6_49;
  reg                 io_A_Valid_3_delay_7_48;
  reg                 io_A_Valid_3_delay_8_47;
  reg                 io_A_Valid_3_delay_9_46;
  reg                 io_A_Valid_3_delay_10_45;
  reg                 io_A_Valid_3_delay_11_44;
  reg                 io_A_Valid_3_delay_12_43;
  reg                 io_A_Valid_3_delay_13_42;
  reg                 io_A_Valid_3_delay_14_41;
  reg                 io_A_Valid_3_delay_15_40;
  reg                 io_A_Valid_3_delay_16_39;
  reg                 io_A_Valid_3_delay_17_38;
  reg                 io_A_Valid_3_delay_18_37;
  reg                 io_A_Valid_3_delay_19_36;
  reg                 io_A_Valid_3_delay_20_35;
  reg                 io_A_Valid_3_delay_21_34;
  reg                 io_A_Valid_3_delay_22_33;
  reg                 io_A_Valid_3_delay_23_32;
  reg                 io_A_Valid_3_delay_24_31;
  reg                 io_A_Valid_3_delay_25_30;
  reg                 io_A_Valid_3_delay_26_29;
  reg                 io_A_Valid_3_delay_27_28;
  reg                 io_A_Valid_3_delay_28_27;
  reg                 io_A_Valid_3_delay_29_26;
  reg                 io_A_Valid_3_delay_30_25;
  reg                 io_A_Valid_3_delay_31_24;
  reg                 io_A_Valid_3_delay_32_23;
  reg                 io_A_Valid_3_delay_33_22;
  reg                 io_A_Valid_3_delay_34_21;
  reg                 io_A_Valid_3_delay_35_20;
  reg                 io_A_Valid_3_delay_36_19;
  reg                 io_A_Valid_3_delay_37_18;
  reg                 io_A_Valid_3_delay_38_17;
  reg                 io_A_Valid_3_delay_39_16;
  reg                 io_A_Valid_3_delay_40_15;
  reg                 io_A_Valid_3_delay_41_14;
  reg                 io_A_Valid_3_delay_42_13;
  reg                 io_A_Valid_3_delay_43_12;
  reg                 io_A_Valid_3_delay_44_11;
  reg                 io_A_Valid_3_delay_45_10;
  reg                 io_A_Valid_3_delay_46_9;
  reg                 io_A_Valid_3_delay_47_8;
  reg                 io_A_Valid_3_delay_48_7;
  reg                 io_A_Valid_3_delay_49_6;
  reg                 io_A_Valid_3_delay_50_5;
  reg                 io_A_Valid_3_delay_51_4;
  reg                 io_A_Valid_3_delay_52_3;
  reg                 io_A_Valid_3_delay_53_2;
  reg                 io_A_Valid_3_delay_54_1;
  reg                 io_A_Valid_3_delay_55;
  reg                 io_B_Valid_55_delay_1_2;
  reg                 io_B_Valid_55_delay_2_1;
  reg                 io_B_Valid_55_delay_3;
  reg                 io_A_Valid_3_delay_1_55;
  reg                 io_A_Valid_3_delay_2_54;
  reg                 io_A_Valid_3_delay_3_53;
  reg                 io_A_Valid_3_delay_4_52;
  reg                 io_A_Valid_3_delay_5_51;
  reg                 io_A_Valid_3_delay_6_50;
  reg                 io_A_Valid_3_delay_7_49;
  reg                 io_A_Valid_3_delay_8_48;
  reg                 io_A_Valid_3_delay_9_47;
  reg                 io_A_Valid_3_delay_10_46;
  reg                 io_A_Valid_3_delay_11_45;
  reg                 io_A_Valid_3_delay_12_44;
  reg                 io_A_Valid_3_delay_13_43;
  reg                 io_A_Valid_3_delay_14_42;
  reg                 io_A_Valid_3_delay_15_41;
  reg                 io_A_Valid_3_delay_16_40;
  reg                 io_A_Valid_3_delay_17_39;
  reg                 io_A_Valid_3_delay_18_38;
  reg                 io_A_Valid_3_delay_19_37;
  reg                 io_A_Valid_3_delay_20_36;
  reg                 io_A_Valid_3_delay_21_35;
  reg                 io_A_Valid_3_delay_22_34;
  reg                 io_A_Valid_3_delay_23_33;
  reg                 io_A_Valid_3_delay_24_32;
  reg                 io_A_Valid_3_delay_25_31;
  reg                 io_A_Valid_3_delay_26_30;
  reg                 io_A_Valid_3_delay_27_29;
  reg                 io_A_Valid_3_delay_28_28;
  reg                 io_A_Valid_3_delay_29_27;
  reg                 io_A_Valid_3_delay_30_26;
  reg                 io_A_Valid_3_delay_31_25;
  reg                 io_A_Valid_3_delay_32_24;
  reg                 io_A_Valid_3_delay_33_23;
  reg                 io_A_Valid_3_delay_34_22;
  reg                 io_A_Valid_3_delay_35_21;
  reg                 io_A_Valid_3_delay_36_20;
  reg                 io_A_Valid_3_delay_37_19;
  reg                 io_A_Valid_3_delay_38_18;
  reg                 io_A_Valid_3_delay_39_17;
  reg                 io_A_Valid_3_delay_40_16;
  reg                 io_A_Valid_3_delay_41_15;
  reg                 io_A_Valid_3_delay_42_14;
  reg                 io_A_Valid_3_delay_43_13;
  reg                 io_A_Valid_3_delay_44_12;
  reg                 io_A_Valid_3_delay_45_11;
  reg                 io_A_Valid_3_delay_46_10;
  reg                 io_A_Valid_3_delay_47_9;
  reg                 io_A_Valid_3_delay_48_8;
  reg                 io_A_Valid_3_delay_49_7;
  reg                 io_A_Valid_3_delay_50_6;
  reg                 io_A_Valid_3_delay_51_5;
  reg                 io_A_Valid_3_delay_52_4;
  reg                 io_A_Valid_3_delay_53_3;
  reg                 io_A_Valid_3_delay_54_2;
  reg                 io_A_Valid_3_delay_55_1;
  reg                 io_A_Valid_3_delay_56;
  reg                 io_B_Valid_56_delay_1_2;
  reg                 io_B_Valid_56_delay_2_1;
  reg                 io_B_Valid_56_delay_3;
  reg                 io_A_Valid_3_delay_1_56;
  reg                 io_A_Valid_3_delay_2_55;
  reg                 io_A_Valid_3_delay_3_54;
  reg                 io_A_Valid_3_delay_4_53;
  reg                 io_A_Valid_3_delay_5_52;
  reg                 io_A_Valid_3_delay_6_51;
  reg                 io_A_Valid_3_delay_7_50;
  reg                 io_A_Valid_3_delay_8_49;
  reg                 io_A_Valid_3_delay_9_48;
  reg                 io_A_Valid_3_delay_10_47;
  reg                 io_A_Valid_3_delay_11_46;
  reg                 io_A_Valid_3_delay_12_45;
  reg                 io_A_Valid_3_delay_13_44;
  reg                 io_A_Valid_3_delay_14_43;
  reg                 io_A_Valid_3_delay_15_42;
  reg                 io_A_Valid_3_delay_16_41;
  reg                 io_A_Valid_3_delay_17_40;
  reg                 io_A_Valid_3_delay_18_39;
  reg                 io_A_Valid_3_delay_19_38;
  reg                 io_A_Valid_3_delay_20_37;
  reg                 io_A_Valid_3_delay_21_36;
  reg                 io_A_Valid_3_delay_22_35;
  reg                 io_A_Valid_3_delay_23_34;
  reg                 io_A_Valid_3_delay_24_33;
  reg                 io_A_Valid_3_delay_25_32;
  reg                 io_A_Valid_3_delay_26_31;
  reg                 io_A_Valid_3_delay_27_30;
  reg                 io_A_Valid_3_delay_28_29;
  reg                 io_A_Valid_3_delay_29_28;
  reg                 io_A_Valid_3_delay_30_27;
  reg                 io_A_Valid_3_delay_31_26;
  reg                 io_A_Valid_3_delay_32_25;
  reg                 io_A_Valid_3_delay_33_24;
  reg                 io_A_Valid_3_delay_34_23;
  reg                 io_A_Valid_3_delay_35_22;
  reg                 io_A_Valid_3_delay_36_21;
  reg                 io_A_Valid_3_delay_37_20;
  reg                 io_A_Valid_3_delay_38_19;
  reg                 io_A_Valid_3_delay_39_18;
  reg                 io_A_Valid_3_delay_40_17;
  reg                 io_A_Valid_3_delay_41_16;
  reg                 io_A_Valid_3_delay_42_15;
  reg                 io_A_Valid_3_delay_43_14;
  reg                 io_A_Valid_3_delay_44_13;
  reg                 io_A_Valid_3_delay_45_12;
  reg                 io_A_Valid_3_delay_46_11;
  reg                 io_A_Valid_3_delay_47_10;
  reg                 io_A_Valid_3_delay_48_9;
  reg                 io_A_Valid_3_delay_49_8;
  reg                 io_A_Valid_3_delay_50_7;
  reg                 io_A_Valid_3_delay_51_6;
  reg                 io_A_Valid_3_delay_52_5;
  reg                 io_A_Valid_3_delay_53_4;
  reg                 io_A_Valid_3_delay_54_3;
  reg                 io_A_Valid_3_delay_55_2;
  reg                 io_A_Valid_3_delay_56_1;
  reg                 io_A_Valid_3_delay_57;
  reg                 io_B_Valid_57_delay_1_2;
  reg                 io_B_Valid_57_delay_2_1;
  reg                 io_B_Valid_57_delay_3;
  reg                 io_A_Valid_3_delay_1_57;
  reg                 io_A_Valid_3_delay_2_56;
  reg                 io_A_Valid_3_delay_3_55;
  reg                 io_A_Valid_3_delay_4_54;
  reg                 io_A_Valid_3_delay_5_53;
  reg                 io_A_Valid_3_delay_6_52;
  reg                 io_A_Valid_3_delay_7_51;
  reg                 io_A_Valid_3_delay_8_50;
  reg                 io_A_Valid_3_delay_9_49;
  reg                 io_A_Valid_3_delay_10_48;
  reg                 io_A_Valid_3_delay_11_47;
  reg                 io_A_Valid_3_delay_12_46;
  reg                 io_A_Valid_3_delay_13_45;
  reg                 io_A_Valid_3_delay_14_44;
  reg                 io_A_Valid_3_delay_15_43;
  reg                 io_A_Valid_3_delay_16_42;
  reg                 io_A_Valid_3_delay_17_41;
  reg                 io_A_Valid_3_delay_18_40;
  reg                 io_A_Valid_3_delay_19_39;
  reg                 io_A_Valid_3_delay_20_38;
  reg                 io_A_Valid_3_delay_21_37;
  reg                 io_A_Valid_3_delay_22_36;
  reg                 io_A_Valid_3_delay_23_35;
  reg                 io_A_Valid_3_delay_24_34;
  reg                 io_A_Valid_3_delay_25_33;
  reg                 io_A_Valid_3_delay_26_32;
  reg                 io_A_Valid_3_delay_27_31;
  reg                 io_A_Valid_3_delay_28_30;
  reg                 io_A_Valid_3_delay_29_29;
  reg                 io_A_Valid_3_delay_30_28;
  reg                 io_A_Valid_3_delay_31_27;
  reg                 io_A_Valid_3_delay_32_26;
  reg                 io_A_Valid_3_delay_33_25;
  reg                 io_A_Valid_3_delay_34_24;
  reg                 io_A_Valid_3_delay_35_23;
  reg                 io_A_Valid_3_delay_36_22;
  reg                 io_A_Valid_3_delay_37_21;
  reg                 io_A_Valid_3_delay_38_20;
  reg                 io_A_Valid_3_delay_39_19;
  reg                 io_A_Valid_3_delay_40_18;
  reg                 io_A_Valid_3_delay_41_17;
  reg                 io_A_Valid_3_delay_42_16;
  reg                 io_A_Valid_3_delay_43_15;
  reg                 io_A_Valid_3_delay_44_14;
  reg                 io_A_Valid_3_delay_45_13;
  reg                 io_A_Valid_3_delay_46_12;
  reg                 io_A_Valid_3_delay_47_11;
  reg                 io_A_Valid_3_delay_48_10;
  reg                 io_A_Valid_3_delay_49_9;
  reg                 io_A_Valid_3_delay_50_8;
  reg                 io_A_Valid_3_delay_51_7;
  reg                 io_A_Valid_3_delay_52_6;
  reg                 io_A_Valid_3_delay_53_5;
  reg                 io_A_Valid_3_delay_54_4;
  reg                 io_A_Valid_3_delay_55_3;
  reg                 io_A_Valid_3_delay_56_2;
  reg                 io_A_Valid_3_delay_57_1;
  reg                 io_A_Valid_3_delay_58;
  reg                 io_B_Valid_58_delay_1_2;
  reg                 io_B_Valid_58_delay_2_1;
  reg                 io_B_Valid_58_delay_3;
  reg                 io_A_Valid_3_delay_1_58;
  reg                 io_A_Valid_3_delay_2_57;
  reg                 io_A_Valid_3_delay_3_56;
  reg                 io_A_Valid_3_delay_4_55;
  reg                 io_A_Valid_3_delay_5_54;
  reg                 io_A_Valid_3_delay_6_53;
  reg                 io_A_Valid_3_delay_7_52;
  reg                 io_A_Valid_3_delay_8_51;
  reg                 io_A_Valid_3_delay_9_50;
  reg                 io_A_Valid_3_delay_10_49;
  reg                 io_A_Valid_3_delay_11_48;
  reg                 io_A_Valid_3_delay_12_47;
  reg                 io_A_Valid_3_delay_13_46;
  reg                 io_A_Valid_3_delay_14_45;
  reg                 io_A_Valid_3_delay_15_44;
  reg                 io_A_Valid_3_delay_16_43;
  reg                 io_A_Valid_3_delay_17_42;
  reg                 io_A_Valid_3_delay_18_41;
  reg                 io_A_Valid_3_delay_19_40;
  reg                 io_A_Valid_3_delay_20_39;
  reg                 io_A_Valid_3_delay_21_38;
  reg                 io_A_Valid_3_delay_22_37;
  reg                 io_A_Valid_3_delay_23_36;
  reg                 io_A_Valid_3_delay_24_35;
  reg                 io_A_Valid_3_delay_25_34;
  reg                 io_A_Valid_3_delay_26_33;
  reg                 io_A_Valid_3_delay_27_32;
  reg                 io_A_Valid_3_delay_28_31;
  reg                 io_A_Valid_3_delay_29_30;
  reg                 io_A_Valid_3_delay_30_29;
  reg                 io_A_Valid_3_delay_31_28;
  reg                 io_A_Valid_3_delay_32_27;
  reg                 io_A_Valid_3_delay_33_26;
  reg                 io_A_Valid_3_delay_34_25;
  reg                 io_A_Valid_3_delay_35_24;
  reg                 io_A_Valid_3_delay_36_23;
  reg                 io_A_Valid_3_delay_37_22;
  reg                 io_A_Valid_3_delay_38_21;
  reg                 io_A_Valid_3_delay_39_20;
  reg                 io_A_Valid_3_delay_40_19;
  reg                 io_A_Valid_3_delay_41_18;
  reg                 io_A_Valid_3_delay_42_17;
  reg                 io_A_Valid_3_delay_43_16;
  reg                 io_A_Valid_3_delay_44_15;
  reg                 io_A_Valid_3_delay_45_14;
  reg                 io_A_Valid_3_delay_46_13;
  reg                 io_A_Valid_3_delay_47_12;
  reg                 io_A_Valid_3_delay_48_11;
  reg                 io_A_Valid_3_delay_49_10;
  reg                 io_A_Valid_3_delay_50_9;
  reg                 io_A_Valid_3_delay_51_8;
  reg                 io_A_Valid_3_delay_52_7;
  reg                 io_A_Valid_3_delay_53_6;
  reg                 io_A_Valid_3_delay_54_5;
  reg                 io_A_Valid_3_delay_55_4;
  reg                 io_A_Valid_3_delay_56_3;
  reg                 io_A_Valid_3_delay_57_2;
  reg                 io_A_Valid_3_delay_58_1;
  reg                 io_A_Valid_3_delay_59;
  reg                 io_B_Valid_59_delay_1_2;
  reg                 io_B_Valid_59_delay_2_1;
  reg                 io_B_Valid_59_delay_3;
  reg                 io_A_Valid_3_delay_1_59;
  reg                 io_A_Valid_3_delay_2_58;
  reg                 io_A_Valid_3_delay_3_57;
  reg                 io_A_Valid_3_delay_4_56;
  reg                 io_A_Valid_3_delay_5_55;
  reg                 io_A_Valid_3_delay_6_54;
  reg                 io_A_Valid_3_delay_7_53;
  reg                 io_A_Valid_3_delay_8_52;
  reg                 io_A_Valid_3_delay_9_51;
  reg                 io_A_Valid_3_delay_10_50;
  reg                 io_A_Valid_3_delay_11_49;
  reg                 io_A_Valid_3_delay_12_48;
  reg                 io_A_Valid_3_delay_13_47;
  reg                 io_A_Valid_3_delay_14_46;
  reg                 io_A_Valid_3_delay_15_45;
  reg                 io_A_Valid_3_delay_16_44;
  reg                 io_A_Valid_3_delay_17_43;
  reg                 io_A_Valid_3_delay_18_42;
  reg                 io_A_Valid_3_delay_19_41;
  reg                 io_A_Valid_3_delay_20_40;
  reg                 io_A_Valid_3_delay_21_39;
  reg                 io_A_Valid_3_delay_22_38;
  reg                 io_A_Valid_3_delay_23_37;
  reg                 io_A_Valid_3_delay_24_36;
  reg                 io_A_Valid_3_delay_25_35;
  reg                 io_A_Valid_3_delay_26_34;
  reg                 io_A_Valid_3_delay_27_33;
  reg                 io_A_Valid_3_delay_28_32;
  reg                 io_A_Valid_3_delay_29_31;
  reg                 io_A_Valid_3_delay_30_30;
  reg                 io_A_Valid_3_delay_31_29;
  reg                 io_A_Valid_3_delay_32_28;
  reg                 io_A_Valid_3_delay_33_27;
  reg                 io_A_Valid_3_delay_34_26;
  reg                 io_A_Valid_3_delay_35_25;
  reg                 io_A_Valid_3_delay_36_24;
  reg                 io_A_Valid_3_delay_37_23;
  reg                 io_A_Valid_3_delay_38_22;
  reg                 io_A_Valid_3_delay_39_21;
  reg                 io_A_Valid_3_delay_40_20;
  reg                 io_A_Valid_3_delay_41_19;
  reg                 io_A_Valid_3_delay_42_18;
  reg                 io_A_Valid_3_delay_43_17;
  reg                 io_A_Valid_3_delay_44_16;
  reg                 io_A_Valid_3_delay_45_15;
  reg                 io_A_Valid_3_delay_46_14;
  reg                 io_A_Valid_3_delay_47_13;
  reg                 io_A_Valid_3_delay_48_12;
  reg                 io_A_Valid_3_delay_49_11;
  reg                 io_A_Valid_3_delay_50_10;
  reg                 io_A_Valid_3_delay_51_9;
  reg                 io_A_Valid_3_delay_52_8;
  reg                 io_A_Valid_3_delay_53_7;
  reg                 io_A_Valid_3_delay_54_6;
  reg                 io_A_Valid_3_delay_55_5;
  reg                 io_A_Valid_3_delay_56_4;
  reg                 io_A_Valid_3_delay_57_3;
  reg                 io_A_Valid_3_delay_58_2;
  reg                 io_A_Valid_3_delay_59_1;
  reg                 io_A_Valid_3_delay_60;
  reg                 io_B_Valid_60_delay_1_2;
  reg                 io_B_Valid_60_delay_2_1;
  reg                 io_B_Valid_60_delay_3;
  reg                 io_A_Valid_3_delay_1_60;
  reg                 io_A_Valid_3_delay_2_59;
  reg                 io_A_Valid_3_delay_3_58;
  reg                 io_A_Valid_3_delay_4_57;
  reg                 io_A_Valid_3_delay_5_56;
  reg                 io_A_Valid_3_delay_6_55;
  reg                 io_A_Valid_3_delay_7_54;
  reg                 io_A_Valid_3_delay_8_53;
  reg                 io_A_Valid_3_delay_9_52;
  reg                 io_A_Valid_3_delay_10_51;
  reg                 io_A_Valid_3_delay_11_50;
  reg                 io_A_Valid_3_delay_12_49;
  reg                 io_A_Valid_3_delay_13_48;
  reg                 io_A_Valid_3_delay_14_47;
  reg                 io_A_Valid_3_delay_15_46;
  reg                 io_A_Valid_3_delay_16_45;
  reg                 io_A_Valid_3_delay_17_44;
  reg                 io_A_Valid_3_delay_18_43;
  reg                 io_A_Valid_3_delay_19_42;
  reg                 io_A_Valid_3_delay_20_41;
  reg                 io_A_Valid_3_delay_21_40;
  reg                 io_A_Valid_3_delay_22_39;
  reg                 io_A_Valid_3_delay_23_38;
  reg                 io_A_Valid_3_delay_24_37;
  reg                 io_A_Valid_3_delay_25_36;
  reg                 io_A_Valid_3_delay_26_35;
  reg                 io_A_Valid_3_delay_27_34;
  reg                 io_A_Valid_3_delay_28_33;
  reg                 io_A_Valid_3_delay_29_32;
  reg                 io_A_Valid_3_delay_30_31;
  reg                 io_A_Valid_3_delay_31_30;
  reg                 io_A_Valid_3_delay_32_29;
  reg                 io_A_Valid_3_delay_33_28;
  reg                 io_A_Valid_3_delay_34_27;
  reg                 io_A_Valid_3_delay_35_26;
  reg                 io_A_Valid_3_delay_36_25;
  reg                 io_A_Valid_3_delay_37_24;
  reg                 io_A_Valid_3_delay_38_23;
  reg                 io_A_Valid_3_delay_39_22;
  reg                 io_A_Valid_3_delay_40_21;
  reg                 io_A_Valid_3_delay_41_20;
  reg                 io_A_Valid_3_delay_42_19;
  reg                 io_A_Valid_3_delay_43_18;
  reg                 io_A_Valid_3_delay_44_17;
  reg                 io_A_Valid_3_delay_45_16;
  reg                 io_A_Valid_3_delay_46_15;
  reg                 io_A_Valid_3_delay_47_14;
  reg                 io_A_Valid_3_delay_48_13;
  reg                 io_A_Valid_3_delay_49_12;
  reg                 io_A_Valid_3_delay_50_11;
  reg                 io_A_Valid_3_delay_51_10;
  reg                 io_A_Valid_3_delay_52_9;
  reg                 io_A_Valid_3_delay_53_8;
  reg                 io_A_Valid_3_delay_54_7;
  reg                 io_A_Valid_3_delay_55_6;
  reg                 io_A_Valid_3_delay_56_5;
  reg                 io_A_Valid_3_delay_57_4;
  reg                 io_A_Valid_3_delay_58_3;
  reg                 io_A_Valid_3_delay_59_2;
  reg                 io_A_Valid_3_delay_60_1;
  reg                 io_A_Valid_3_delay_61;
  reg                 io_B_Valid_61_delay_1_2;
  reg                 io_B_Valid_61_delay_2_1;
  reg                 io_B_Valid_61_delay_3;
  reg                 io_A_Valid_3_delay_1_61;
  reg                 io_A_Valid_3_delay_2_60;
  reg                 io_A_Valid_3_delay_3_59;
  reg                 io_A_Valid_3_delay_4_58;
  reg                 io_A_Valid_3_delay_5_57;
  reg                 io_A_Valid_3_delay_6_56;
  reg                 io_A_Valid_3_delay_7_55;
  reg                 io_A_Valid_3_delay_8_54;
  reg                 io_A_Valid_3_delay_9_53;
  reg                 io_A_Valid_3_delay_10_52;
  reg                 io_A_Valid_3_delay_11_51;
  reg                 io_A_Valid_3_delay_12_50;
  reg                 io_A_Valid_3_delay_13_49;
  reg                 io_A_Valid_3_delay_14_48;
  reg                 io_A_Valid_3_delay_15_47;
  reg                 io_A_Valid_3_delay_16_46;
  reg                 io_A_Valid_3_delay_17_45;
  reg                 io_A_Valid_3_delay_18_44;
  reg                 io_A_Valid_3_delay_19_43;
  reg                 io_A_Valid_3_delay_20_42;
  reg                 io_A_Valid_3_delay_21_41;
  reg                 io_A_Valid_3_delay_22_40;
  reg                 io_A_Valid_3_delay_23_39;
  reg                 io_A_Valid_3_delay_24_38;
  reg                 io_A_Valid_3_delay_25_37;
  reg                 io_A_Valid_3_delay_26_36;
  reg                 io_A_Valid_3_delay_27_35;
  reg                 io_A_Valid_3_delay_28_34;
  reg                 io_A_Valid_3_delay_29_33;
  reg                 io_A_Valid_3_delay_30_32;
  reg                 io_A_Valid_3_delay_31_31;
  reg                 io_A_Valid_3_delay_32_30;
  reg                 io_A_Valid_3_delay_33_29;
  reg                 io_A_Valid_3_delay_34_28;
  reg                 io_A_Valid_3_delay_35_27;
  reg                 io_A_Valid_3_delay_36_26;
  reg                 io_A_Valid_3_delay_37_25;
  reg                 io_A_Valid_3_delay_38_24;
  reg                 io_A_Valid_3_delay_39_23;
  reg                 io_A_Valid_3_delay_40_22;
  reg                 io_A_Valid_3_delay_41_21;
  reg                 io_A_Valid_3_delay_42_20;
  reg                 io_A_Valid_3_delay_43_19;
  reg                 io_A_Valid_3_delay_44_18;
  reg                 io_A_Valid_3_delay_45_17;
  reg                 io_A_Valid_3_delay_46_16;
  reg                 io_A_Valid_3_delay_47_15;
  reg                 io_A_Valid_3_delay_48_14;
  reg                 io_A_Valid_3_delay_49_13;
  reg                 io_A_Valid_3_delay_50_12;
  reg                 io_A_Valid_3_delay_51_11;
  reg                 io_A_Valid_3_delay_52_10;
  reg                 io_A_Valid_3_delay_53_9;
  reg                 io_A_Valid_3_delay_54_8;
  reg                 io_A_Valid_3_delay_55_7;
  reg                 io_A_Valid_3_delay_56_6;
  reg                 io_A_Valid_3_delay_57_5;
  reg                 io_A_Valid_3_delay_58_4;
  reg                 io_A_Valid_3_delay_59_3;
  reg                 io_A_Valid_3_delay_60_2;
  reg                 io_A_Valid_3_delay_61_1;
  reg                 io_A_Valid_3_delay_62;
  reg                 io_B_Valid_62_delay_1_2;
  reg                 io_B_Valid_62_delay_2_1;
  reg                 io_B_Valid_62_delay_3;
  reg                 io_A_Valid_3_delay_1_62;
  reg                 io_A_Valid_3_delay_2_61;
  reg                 io_A_Valid_3_delay_3_60;
  reg                 io_A_Valid_3_delay_4_59;
  reg                 io_A_Valid_3_delay_5_58;
  reg                 io_A_Valid_3_delay_6_57;
  reg                 io_A_Valid_3_delay_7_56;
  reg                 io_A_Valid_3_delay_8_55;
  reg                 io_A_Valid_3_delay_9_54;
  reg                 io_A_Valid_3_delay_10_53;
  reg                 io_A_Valid_3_delay_11_52;
  reg                 io_A_Valid_3_delay_12_51;
  reg                 io_A_Valid_3_delay_13_50;
  reg                 io_A_Valid_3_delay_14_49;
  reg                 io_A_Valid_3_delay_15_48;
  reg                 io_A_Valid_3_delay_16_47;
  reg                 io_A_Valid_3_delay_17_46;
  reg                 io_A_Valid_3_delay_18_45;
  reg                 io_A_Valid_3_delay_19_44;
  reg                 io_A_Valid_3_delay_20_43;
  reg                 io_A_Valid_3_delay_21_42;
  reg                 io_A_Valid_3_delay_22_41;
  reg                 io_A_Valid_3_delay_23_40;
  reg                 io_A_Valid_3_delay_24_39;
  reg                 io_A_Valid_3_delay_25_38;
  reg                 io_A_Valid_3_delay_26_37;
  reg                 io_A_Valid_3_delay_27_36;
  reg                 io_A_Valid_3_delay_28_35;
  reg                 io_A_Valid_3_delay_29_34;
  reg                 io_A_Valid_3_delay_30_33;
  reg                 io_A_Valid_3_delay_31_32;
  reg                 io_A_Valid_3_delay_32_31;
  reg                 io_A_Valid_3_delay_33_30;
  reg                 io_A_Valid_3_delay_34_29;
  reg                 io_A_Valid_3_delay_35_28;
  reg                 io_A_Valid_3_delay_36_27;
  reg                 io_A_Valid_3_delay_37_26;
  reg                 io_A_Valid_3_delay_38_25;
  reg                 io_A_Valid_3_delay_39_24;
  reg                 io_A_Valid_3_delay_40_23;
  reg                 io_A_Valid_3_delay_41_22;
  reg                 io_A_Valid_3_delay_42_21;
  reg                 io_A_Valid_3_delay_43_20;
  reg                 io_A_Valid_3_delay_44_19;
  reg                 io_A_Valid_3_delay_45_18;
  reg                 io_A_Valid_3_delay_46_17;
  reg                 io_A_Valid_3_delay_47_16;
  reg                 io_A_Valid_3_delay_48_15;
  reg                 io_A_Valid_3_delay_49_14;
  reg                 io_A_Valid_3_delay_50_13;
  reg                 io_A_Valid_3_delay_51_12;
  reg                 io_A_Valid_3_delay_52_11;
  reg                 io_A_Valid_3_delay_53_10;
  reg                 io_A_Valid_3_delay_54_9;
  reg                 io_A_Valid_3_delay_55_8;
  reg                 io_A_Valid_3_delay_56_7;
  reg                 io_A_Valid_3_delay_57_6;
  reg                 io_A_Valid_3_delay_58_5;
  reg                 io_A_Valid_3_delay_59_4;
  reg                 io_A_Valid_3_delay_60_3;
  reg                 io_A_Valid_3_delay_61_2;
  reg                 io_A_Valid_3_delay_62_1;
  reg                 io_A_Valid_3_delay_63;
  reg                 io_B_Valid_63_delay_1_2;
  reg                 io_B_Valid_63_delay_2_1;
  reg                 io_B_Valid_63_delay_3;
  reg        [15:0]   io_signCount_regNextWhen_4;
  reg                 io_B_Valid_0_delay_1_3;
  reg                 io_B_Valid_0_delay_2_2;
  reg                 io_B_Valid_0_delay_3_1;
  reg                 io_B_Valid_0_delay_4;
  reg                 io_A_Valid_4_delay_1;
  reg                 io_B_Valid_1_delay_1_3;
  reg                 io_B_Valid_1_delay_2_2;
  reg                 io_B_Valid_1_delay_3_1;
  reg                 io_B_Valid_1_delay_4;
  reg                 io_A_Valid_4_delay_1_1;
  reg                 io_A_Valid_4_delay_2;
  reg                 io_B_Valid_2_delay_1_3;
  reg                 io_B_Valid_2_delay_2_2;
  reg                 io_B_Valid_2_delay_3_1;
  reg                 io_B_Valid_2_delay_4;
  reg                 io_A_Valid_4_delay_1_2;
  reg                 io_A_Valid_4_delay_2_1;
  reg                 io_A_Valid_4_delay_3;
  reg                 io_B_Valid_3_delay_1_3;
  reg                 io_B_Valid_3_delay_2_2;
  reg                 io_B_Valid_3_delay_3_1;
  reg                 io_B_Valid_3_delay_4;
  reg                 io_A_Valid_4_delay_1_3;
  reg                 io_A_Valid_4_delay_2_2;
  reg                 io_A_Valid_4_delay_3_1;
  reg                 io_A_Valid_4_delay_4;
  reg                 io_B_Valid_4_delay_1_3;
  reg                 io_B_Valid_4_delay_2_2;
  reg                 io_B_Valid_4_delay_3_1;
  reg                 io_B_Valid_4_delay_4;
  reg                 io_A_Valid_4_delay_1_4;
  reg                 io_A_Valid_4_delay_2_3;
  reg                 io_A_Valid_4_delay_3_2;
  reg                 io_A_Valid_4_delay_4_1;
  reg                 io_A_Valid_4_delay_5;
  reg                 io_B_Valid_5_delay_1_3;
  reg                 io_B_Valid_5_delay_2_2;
  reg                 io_B_Valid_5_delay_3_1;
  reg                 io_B_Valid_5_delay_4;
  reg                 io_A_Valid_4_delay_1_5;
  reg                 io_A_Valid_4_delay_2_4;
  reg                 io_A_Valid_4_delay_3_3;
  reg                 io_A_Valid_4_delay_4_2;
  reg                 io_A_Valid_4_delay_5_1;
  reg                 io_A_Valid_4_delay_6;
  reg                 io_B_Valid_6_delay_1_3;
  reg                 io_B_Valid_6_delay_2_2;
  reg                 io_B_Valid_6_delay_3_1;
  reg                 io_B_Valid_6_delay_4;
  reg                 io_A_Valid_4_delay_1_6;
  reg                 io_A_Valid_4_delay_2_5;
  reg                 io_A_Valid_4_delay_3_4;
  reg                 io_A_Valid_4_delay_4_3;
  reg                 io_A_Valid_4_delay_5_2;
  reg                 io_A_Valid_4_delay_6_1;
  reg                 io_A_Valid_4_delay_7;
  reg                 io_B_Valid_7_delay_1_3;
  reg                 io_B_Valid_7_delay_2_2;
  reg                 io_B_Valid_7_delay_3_1;
  reg                 io_B_Valid_7_delay_4;
  reg                 io_A_Valid_4_delay_1_7;
  reg                 io_A_Valid_4_delay_2_6;
  reg                 io_A_Valid_4_delay_3_5;
  reg                 io_A_Valid_4_delay_4_4;
  reg                 io_A_Valid_4_delay_5_3;
  reg                 io_A_Valid_4_delay_6_2;
  reg                 io_A_Valid_4_delay_7_1;
  reg                 io_A_Valid_4_delay_8;
  reg                 io_B_Valid_8_delay_1_3;
  reg                 io_B_Valid_8_delay_2_2;
  reg                 io_B_Valid_8_delay_3_1;
  reg                 io_B_Valid_8_delay_4;
  reg                 io_A_Valid_4_delay_1_8;
  reg                 io_A_Valid_4_delay_2_7;
  reg                 io_A_Valid_4_delay_3_6;
  reg                 io_A_Valid_4_delay_4_5;
  reg                 io_A_Valid_4_delay_5_4;
  reg                 io_A_Valid_4_delay_6_3;
  reg                 io_A_Valid_4_delay_7_2;
  reg                 io_A_Valid_4_delay_8_1;
  reg                 io_A_Valid_4_delay_9;
  reg                 io_B_Valid_9_delay_1_3;
  reg                 io_B_Valid_9_delay_2_2;
  reg                 io_B_Valid_9_delay_3_1;
  reg                 io_B_Valid_9_delay_4;
  reg                 io_A_Valid_4_delay_1_9;
  reg                 io_A_Valid_4_delay_2_8;
  reg                 io_A_Valid_4_delay_3_7;
  reg                 io_A_Valid_4_delay_4_6;
  reg                 io_A_Valid_4_delay_5_5;
  reg                 io_A_Valid_4_delay_6_4;
  reg                 io_A_Valid_4_delay_7_3;
  reg                 io_A_Valid_4_delay_8_2;
  reg                 io_A_Valid_4_delay_9_1;
  reg                 io_A_Valid_4_delay_10;
  reg                 io_B_Valid_10_delay_1_3;
  reg                 io_B_Valid_10_delay_2_2;
  reg                 io_B_Valid_10_delay_3_1;
  reg                 io_B_Valid_10_delay_4;
  reg                 io_A_Valid_4_delay_1_10;
  reg                 io_A_Valid_4_delay_2_9;
  reg                 io_A_Valid_4_delay_3_8;
  reg                 io_A_Valid_4_delay_4_7;
  reg                 io_A_Valid_4_delay_5_6;
  reg                 io_A_Valid_4_delay_6_5;
  reg                 io_A_Valid_4_delay_7_4;
  reg                 io_A_Valid_4_delay_8_3;
  reg                 io_A_Valid_4_delay_9_2;
  reg                 io_A_Valid_4_delay_10_1;
  reg                 io_A_Valid_4_delay_11;
  reg                 io_B_Valid_11_delay_1_3;
  reg                 io_B_Valid_11_delay_2_2;
  reg                 io_B_Valid_11_delay_3_1;
  reg                 io_B_Valid_11_delay_4;
  reg                 io_A_Valid_4_delay_1_11;
  reg                 io_A_Valid_4_delay_2_10;
  reg                 io_A_Valid_4_delay_3_9;
  reg                 io_A_Valid_4_delay_4_8;
  reg                 io_A_Valid_4_delay_5_7;
  reg                 io_A_Valid_4_delay_6_6;
  reg                 io_A_Valid_4_delay_7_5;
  reg                 io_A_Valid_4_delay_8_4;
  reg                 io_A_Valid_4_delay_9_3;
  reg                 io_A_Valid_4_delay_10_2;
  reg                 io_A_Valid_4_delay_11_1;
  reg                 io_A_Valid_4_delay_12;
  reg                 io_B_Valid_12_delay_1_3;
  reg                 io_B_Valid_12_delay_2_2;
  reg                 io_B_Valid_12_delay_3_1;
  reg                 io_B_Valid_12_delay_4;
  reg                 io_A_Valid_4_delay_1_12;
  reg                 io_A_Valid_4_delay_2_11;
  reg                 io_A_Valid_4_delay_3_10;
  reg                 io_A_Valid_4_delay_4_9;
  reg                 io_A_Valid_4_delay_5_8;
  reg                 io_A_Valid_4_delay_6_7;
  reg                 io_A_Valid_4_delay_7_6;
  reg                 io_A_Valid_4_delay_8_5;
  reg                 io_A_Valid_4_delay_9_4;
  reg                 io_A_Valid_4_delay_10_3;
  reg                 io_A_Valid_4_delay_11_2;
  reg                 io_A_Valid_4_delay_12_1;
  reg                 io_A_Valid_4_delay_13;
  reg                 io_B_Valid_13_delay_1_3;
  reg                 io_B_Valid_13_delay_2_2;
  reg                 io_B_Valid_13_delay_3_1;
  reg                 io_B_Valid_13_delay_4;
  reg                 io_A_Valid_4_delay_1_13;
  reg                 io_A_Valid_4_delay_2_12;
  reg                 io_A_Valid_4_delay_3_11;
  reg                 io_A_Valid_4_delay_4_10;
  reg                 io_A_Valid_4_delay_5_9;
  reg                 io_A_Valid_4_delay_6_8;
  reg                 io_A_Valid_4_delay_7_7;
  reg                 io_A_Valid_4_delay_8_6;
  reg                 io_A_Valid_4_delay_9_5;
  reg                 io_A_Valid_4_delay_10_4;
  reg                 io_A_Valid_4_delay_11_3;
  reg                 io_A_Valid_4_delay_12_2;
  reg                 io_A_Valid_4_delay_13_1;
  reg                 io_A_Valid_4_delay_14;
  reg                 io_B_Valid_14_delay_1_3;
  reg                 io_B_Valid_14_delay_2_2;
  reg                 io_B_Valid_14_delay_3_1;
  reg                 io_B_Valid_14_delay_4;
  reg                 io_A_Valid_4_delay_1_14;
  reg                 io_A_Valid_4_delay_2_13;
  reg                 io_A_Valid_4_delay_3_12;
  reg                 io_A_Valid_4_delay_4_11;
  reg                 io_A_Valid_4_delay_5_10;
  reg                 io_A_Valid_4_delay_6_9;
  reg                 io_A_Valid_4_delay_7_8;
  reg                 io_A_Valid_4_delay_8_7;
  reg                 io_A_Valid_4_delay_9_6;
  reg                 io_A_Valid_4_delay_10_5;
  reg                 io_A_Valid_4_delay_11_4;
  reg                 io_A_Valid_4_delay_12_3;
  reg                 io_A_Valid_4_delay_13_2;
  reg                 io_A_Valid_4_delay_14_1;
  reg                 io_A_Valid_4_delay_15;
  reg                 io_B_Valid_15_delay_1_3;
  reg                 io_B_Valid_15_delay_2_2;
  reg                 io_B_Valid_15_delay_3_1;
  reg                 io_B_Valid_15_delay_4;
  reg                 io_A_Valid_4_delay_1_15;
  reg                 io_A_Valid_4_delay_2_14;
  reg                 io_A_Valid_4_delay_3_13;
  reg                 io_A_Valid_4_delay_4_12;
  reg                 io_A_Valid_4_delay_5_11;
  reg                 io_A_Valid_4_delay_6_10;
  reg                 io_A_Valid_4_delay_7_9;
  reg                 io_A_Valid_4_delay_8_8;
  reg                 io_A_Valid_4_delay_9_7;
  reg                 io_A_Valid_4_delay_10_6;
  reg                 io_A_Valid_4_delay_11_5;
  reg                 io_A_Valid_4_delay_12_4;
  reg                 io_A_Valid_4_delay_13_3;
  reg                 io_A_Valid_4_delay_14_2;
  reg                 io_A_Valid_4_delay_15_1;
  reg                 io_A_Valid_4_delay_16;
  reg                 io_B_Valid_16_delay_1_3;
  reg                 io_B_Valid_16_delay_2_2;
  reg                 io_B_Valid_16_delay_3_1;
  reg                 io_B_Valid_16_delay_4;
  reg                 io_A_Valid_4_delay_1_16;
  reg                 io_A_Valid_4_delay_2_15;
  reg                 io_A_Valid_4_delay_3_14;
  reg                 io_A_Valid_4_delay_4_13;
  reg                 io_A_Valid_4_delay_5_12;
  reg                 io_A_Valid_4_delay_6_11;
  reg                 io_A_Valid_4_delay_7_10;
  reg                 io_A_Valid_4_delay_8_9;
  reg                 io_A_Valid_4_delay_9_8;
  reg                 io_A_Valid_4_delay_10_7;
  reg                 io_A_Valid_4_delay_11_6;
  reg                 io_A_Valid_4_delay_12_5;
  reg                 io_A_Valid_4_delay_13_4;
  reg                 io_A_Valid_4_delay_14_3;
  reg                 io_A_Valid_4_delay_15_2;
  reg                 io_A_Valid_4_delay_16_1;
  reg                 io_A_Valid_4_delay_17;
  reg                 io_B_Valid_17_delay_1_3;
  reg                 io_B_Valid_17_delay_2_2;
  reg                 io_B_Valid_17_delay_3_1;
  reg                 io_B_Valid_17_delay_4;
  reg                 io_A_Valid_4_delay_1_17;
  reg                 io_A_Valid_4_delay_2_16;
  reg                 io_A_Valid_4_delay_3_15;
  reg                 io_A_Valid_4_delay_4_14;
  reg                 io_A_Valid_4_delay_5_13;
  reg                 io_A_Valid_4_delay_6_12;
  reg                 io_A_Valid_4_delay_7_11;
  reg                 io_A_Valid_4_delay_8_10;
  reg                 io_A_Valid_4_delay_9_9;
  reg                 io_A_Valid_4_delay_10_8;
  reg                 io_A_Valid_4_delay_11_7;
  reg                 io_A_Valid_4_delay_12_6;
  reg                 io_A_Valid_4_delay_13_5;
  reg                 io_A_Valid_4_delay_14_4;
  reg                 io_A_Valid_4_delay_15_3;
  reg                 io_A_Valid_4_delay_16_2;
  reg                 io_A_Valid_4_delay_17_1;
  reg                 io_A_Valid_4_delay_18;
  reg                 io_B_Valid_18_delay_1_3;
  reg                 io_B_Valid_18_delay_2_2;
  reg                 io_B_Valid_18_delay_3_1;
  reg                 io_B_Valid_18_delay_4;
  reg                 io_A_Valid_4_delay_1_18;
  reg                 io_A_Valid_4_delay_2_17;
  reg                 io_A_Valid_4_delay_3_16;
  reg                 io_A_Valid_4_delay_4_15;
  reg                 io_A_Valid_4_delay_5_14;
  reg                 io_A_Valid_4_delay_6_13;
  reg                 io_A_Valid_4_delay_7_12;
  reg                 io_A_Valid_4_delay_8_11;
  reg                 io_A_Valid_4_delay_9_10;
  reg                 io_A_Valid_4_delay_10_9;
  reg                 io_A_Valid_4_delay_11_8;
  reg                 io_A_Valid_4_delay_12_7;
  reg                 io_A_Valid_4_delay_13_6;
  reg                 io_A_Valid_4_delay_14_5;
  reg                 io_A_Valid_4_delay_15_4;
  reg                 io_A_Valid_4_delay_16_3;
  reg                 io_A_Valid_4_delay_17_2;
  reg                 io_A_Valid_4_delay_18_1;
  reg                 io_A_Valid_4_delay_19;
  reg                 io_B_Valid_19_delay_1_3;
  reg                 io_B_Valid_19_delay_2_2;
  reg                 io_B_Valid_19_delay_3_1;
  reg                 io_B_Valid_19_delay_4;
  reg                 io_A_Valid_4_delay_1_19;
  reg                 io_A_Valid_4_delay_2_18;
  reg                 io_A_Valid_4_delay_3_17;
  reg                 io_A_Valid_4_delay_4_16;
  reg                 io_A_Valid_4_delay_5_15;
  reg                 io_A_Valid_4_delay_6_14;
  reg                 io_A_Valid_4_delay_7_13;
  reg                 io_A_Valid_4_delay_8_12;
  reg                 io_A_Valid_4_delay_9_11;
  reg                 io_A_Valid_4_delay_10_10;
  reg                 io_A_Valid_4_delay_11_9;
  reg                 io_A_Valid_4_delay_12_8;
  reg                 io_A_Valid_4_delay_13_7;
  reg                 io_A_Valid_4_delay_14_6;
  reg                 io_A_Valid_4_delay_15_5;
  reg                 io_A_Valid_4_delay_16_4;
  reg                 io_A_Valid_4_delay_17_3;
  reg                 io_A_Valid_4_delay_18_2;
  reg                 io_A_Valid_4_delay_19_1;
  reg                 io_A_Valid_4_delay_20;
  reg                 io_B_Valid_20_delay_1_3;
  reg                 io_B_Valid_20_delay_2_2;
  reg                 io_B_Valid_20_delay_3_1;
  reg                 io_B_Valid_20_delay_4;
  reg                 io_A_Valid_4_delay_1_20;
  reg                 io_A_Valid_4_delay_2_19;
  reg                 io_A_Valid_4_delay_3_18;
  reg                 io_A_Valid_4_delay_4_17;
  reg                 io_A_Valid_4_delay_5_16;
  reg                 io_A_Valid_4_delay_6_15;
  reg                 io_A_Valid_4_delay_7_14;
  reg                 io_A_Valid_4_delay_8_13;
  reg                 io_A_Valid_4_delay_9_12;
  reg                 io_A_Valid_4_delay_10_11;
  reg                 io_A_Valid_4_delay_11_10;
  reg                 io_A_Valid_4_delay_12_9;
  reg                 io_A_Valid_4_delay_13_8;
  reg                 io_A_Valid_4_delay_14_7;
  reg                 io_A_Valid_4_delay_15_6;
  reg                 io_A_Valid_4_delay_16_5;
  reg                 io_A_Valid_4_delay_17_4;
  reg                 io_A_Valid_4_delay_18_3;
  reg                 io_A_Valid_4_delay_19_2;
  reg                 io_A_Valid_4_delay_20_1;
  reg                 io_A_Valid_4_delay_21;
  reg                 io_B_Valid_21_delay_1_3;
  reg                 io_B_Valid_21_delay_2_2;
  reg                 io_B_Valid_21_delay_3_1;
  reg                 io_B_Valid_21_delay_4;
  reg                 io_A_Valid_4_delay_1_21;
  reg                 io_A_Valid_4_delay_2_20;
  reg                 io_A_Valid_4_delay_3_19;
  reg                 io_A_Valid_4_delay_4_18;
  reg                 io_A_Valid_4_delay_5_17;
  reg                 io_A_Valid_4_delay_6_16;
  reg                 io_A_Valid_4_delay_7_15;
  reg                 io_A_Valid_4_delay_8_14;
  reg                 io_A_Valid_4_delay_9_13;
  reg                 io_A_Valid_4_delay_10_12;
  reg                 io_A_Valid_4_delay_11_11;
  reg                 io_A_Valid_4_delay_12_10;
  reg                 io_A_Valid_4_delay_13_9;
  reg                 io_A_Valid_4_delay_14_8;
  reg                 io_A_Valid_4_delay_15_7;
  reg                 io_A_Valid_4_delay_16_6;
  reg                 io_A_Valid_4_delay_17_5;
  reg                 io_A_Valid_4_delay_18_4;
  reg                 io_A_Valid_4_delay_19_3;
  reg                 io_A_Valid_4_delay_20_2;
  reg                 io_A_Valid_4_delay_21_1;
  reg                 io_A_Valid_4_delay_22;
  reg                 io_B_Valid_22_delay_1_3;
  reg                 io_B_Valid_22_delay_2_2;
  reg                 io_B_Valid_22_delay_3_1;
  reg                 io_B_Valid_22_delay_4;
  reg                 io_A_Valid_4_delay_1_22;
  reg                 io_A_Valid_4_delay_2_21;
  reg                 io_A_Valid_4_delay_3_20;
  reg                 io_A_Valid_4_delay_4_19;
  reg                 io_A_Valid_4_delay_5_18;
  reg                 io_A_Valid_4_delay_6_17;
  reg                 io_A_Valid_4_delay_7_16;
  reg                 io_A_Valid_4_delay_8_15;
  reg                 io_A_Valid_4_delay_9_14;
  reg                 io_A_Valid_4_delay_10_13;
  reg                 io_A_Valid_4_delay_11_12;
  reg                 io_A_Valid_4_delay_12_11;
  reg                 io_A_Valid_4_delay_13_10;
  reg                 io_A_Valid_4_delay_14_9;
  reg                 io_A_Valid_4_delay_15_8;
  reg                 io_A_Valid_4_delay_16_7;
  reg                 io_A_Valid_4_delay_17_6;
  reg                 io_A_Valid_4_delay_18_5;
  reg                 io_A_Valid_4_delay_19_4;
  reg                 io_A_Valid_4_delay_20_3;
  reg                 io_A_Valid_4_delay_21_2;
  reg                 io_A_Valid_4_delay_22_1;
  reg                 io_A_Valid_4_delay_23;
  reg                 io_B_Valid_23_delay_1_3;
  reg                 io_B_Valid_23_delay_2_2;
  reg                 io_B_Valid_23_delay_3_1;
  reg                 io_B_Valid_23_delay_4;
  reg                 io_A_Valid_4_delay_1_23;
  reg                 io_A_Valid_4_delay_2_22;
  reg                 io_A_Valid_4_delay_3_21;
  reg                 io_A_Valid_4_delay_4_20;
  reg                 io_A_Valid_4_delay_5_19;
  reg                 io_A_Valid_4_delay_6_18;
  reg                 io_A_Valid_4_delay_7_17;
  reg                 io_A_Valid_4_delay_8_16;
  reg                 io_A_Valid_4_delay_9_15;
  reg                 io_A_Valid_4_delay_10_14;
  reg                 io_A_Valid_4_delay_11_13;
  reg                 io_A_Valid_4_delay_12_12;
  reg                 io_A_Valid_4_delay_13_11;
  reg                 io_A_Valid_4_delay_14_10;
  reg                 io_A_Valid_4_delay_15_9;
  reg                 io_A_Valid_4_delay_16_8;
  reg                 io_A_Valid_4_delay_17_7;
  reg                 io_A_Valid_4_delay_18_6;
  reg                 io_A_Valid_4_delay_19_5;
  reg                 io_A_Valid_4_delay_20_4;
  reg                 io_A_Valid_4_delay_21_3;
  reg                 io_A_Valid_4_delay_22_2;
  reg                 io_A_Valid_4_delay_23_1;
  reg                 io_A_Valid_4_delay_24;
  reg                 io_B_Valid_24_delay_1_3;
  reg                 io_B_Valid_24_delay_2_2;
  reg                 io_B_Valid_24_delay_3_1;
  reg                 io_B_Valid_24_delay_4;
  reg                 io_A_Valid_4_delay_1_24;
  reg                 io_A_Valid_4_delay_2_23;
  reg                 io_A_Valid_4_delay_3_22;
  reg                 io_A_Valid_4_delay_4_21;
  reg                 io_A_Valid_4_delay_5_20;
  reg                 io_A_Valid_4_delay_6_19;
  reg                 io_A_Valid_4_delay_7_18;
  reg                 io_A_Valid_4_delay_8_17;
  reg                 io_A_Valid_4_delay_9_16;
  reg                 io_A_Valid_4_delay_10_15;
  reg                 io_A_Valid_4_delay_11_14;
  reg                 io_A_Valid_4_delay_12_13;
  reg                 io_A_Valid_4_delay_13_12;
  reg                 io_A_Valid_4_delay_14_11;
  reg                 io_A_Valid_4_delay_15_10;
  reg                 io_A_Valid_4_delay_16_9;
  reg                 io_A_Valid_4_delay_17_8;
  reg                 io_A_Valid_4_delay_18_7;
  reg                 io_A_Valid_4_delay_19_6;
  reg                 io_A_Valid_4_delay_20_5;
  reg                 io_A_Valid_4_delay_21_4;
  reg                 io_A_Valid_4_delay_22_3;
  reg                 io_A_Valid_4_delay_23_2;
  reg                 io_A_Valid_4_delay_24_1;
  reg                 io_A_Valid_4_delay_25;
  reg                 io_B_Valid_25_delay_1_3;
  reg                 io_B_Valid_25_delay_2_2;
  reg                 io_B_Valid_25_delay_3_1;
  reg                 io_B_Valid_25_delay_4;
  reg                 io_A_Valid_4_delay_1_25;
  reg                 io_A_Valid_4_delay_2_24;
  reg                 io_A_Valid_4_delay_3_23;
  reg                 io_A_Valid_4_delay_4_22;
  reg                 io_A_Valid_4_delay_5_21;
  reg                 io_A_Valid_4_delay_6_20;
  reg                 io_A_Valid_4_delay_7_19;
  reg                 io_A_Valid_4_delay_8_18;
  reg                 io_A_Valid_4_delay_9_17;
  reg                 io_A_Valid_4_delay_10_16;
  reg                 io_A_Valid_4_delay_11_15;
  reg                 io_A_Valid_4_delay_12_14;
  reg                 io_A_Valid_4_delay_13_13;
  reg                 io_A_Valid_4_delay_14_12;
  reg                 io_A_Valid_4_delay_15_11;
  reg                 io_A_Valid_4_delay_16_10;
  reg                 io_A_Valid_4_delay_17_9;
  reg                 io_A_Valid_4_delay_18_8;
  reg                 io_A_Valid_4_delay_19_7;
  reg                 io_A_Valid_4_delay_20_6;
  reg                 io_A_Valid_4_delay_21_5;
  reg                 io_A_Valid_4_delay_22_4;
  reg                 io_A_Valid_4_delay_23_3;
  reg                 io_A_Valid_4_delay_24_2;
  reg                 io_A_Valid_4_delay_25_1;
  reg                 io_A_Valid_4_delay_26;
  reg                 io_B_Valid_26_delay_1_3;
  reg                 io_B_Valid_26_delay_2_2;
  reg                 io_B_Valid_26_delay_3_1;
  reg                 io_B_Valid_26_delay_4;
  reg                 io_A_Valid_4_delay_1_26;
  reg                 io_A_Valid_4_delay_2_25;
  reg                 io_A_Valid_4_delay_3_24;
  reg                 io_A_Valid_4_delay_4_23;
  reg                 io_A_Valid_4_delay_5_22;
  reg                 io_A_Valid_4_delay_6_21;
  reg                 io_A_Valid_4_delay_7_20;
  reg                 io_A_Valid_4_delay_8_19;
  reg                 io_A_Valid_4_delay_9_18;
  reg                 io_A_Valid_4_delay_10_17;
  reg                 io_A_Valid_4_delay_11_16;
  reg                 io_A_Valid_4_delay_12_15;
  reg                 io_A_Valid_4_delay_13_14;
  reg                 io_A_Valid_4_delay_14_13;
  reg                 io_A_Valid_4_delay_15_12;
  reg                 io_A_Valid_4_delay_16_11;
  reg                 io_A_Valid_4_delay_17_10;
  reg                 io_A_Valid_4_delay_18_9;
  reg                 io_A_Valid_4_delay_19_8;
  reg                 io_A_Valid_4_delay_20_7;
  reg                 io_A_Valid_4_delay_21_6;
  reg                 io_A_Valid_4_delay_22_5;
  reg                 io_A_Valid_4_delay_23_4;
  reg                 io_A_Valid_4_delay_24_3;
  reg                 io_A_Valid_4_delay_25_2;
  reg                 io_A_Valid_4_delay_26_1;
  reg                 io_A_Valid_4_delay_27;
  reg                 io_B_Valid_27_delay_1_3;
  reg                 io_B_Valid_27_delay_2_2;
  reg                 io_B_Valid_27_delay_3_1;
  reg                 io_B_Valid_27_delay_4;
  reg                 io_A_Valid_4_delay_1_27;
  reg                 io_A_Valid_4_delay_2_26;
  reg                 io_A_Valid_4_delay_3_25;
  reg                 io_A_Valid_4_delay_4_24;
  reg                 io_A_Valid_4_delay_5_23;
  reg                 io_A_Valid_4_delay_6_22;
  reg                 io_A_Valid_4_delay_7_21;
  reg                 io_A_Valid_4_delay_8_20;
  reg                 io_A_Valid_4_delay_9_19;
  reg                 io_A_Valid_4_delay_10_18;
  reg                 io_A_Valid_4_delay_11_17;
  reg                 io_A_Valid_4_delay_12_16;
  reg                 io_A_Valid_4_delay_13_15;
  reg                 io_A_Valid_4_delay_14_14;
  reg                 io_A_Valid_4_delay_15_13;
  reg                 io_A_Valid_4_delay_16_12;
  reg                 io_A_Valid_4_delay_17_11;
  reg                 io_A_Valid_4_delay_18_10;
  reg                 io_A_Valid_4_delay_19_9;
  reg                 io_A_Valid_4_delay_20_8;
  reg                 io_A_Valid_4_delay_21_7;
  reg                 io_A_Valid_4_delay_22_6;
  reg                 io_A_Valid_4_delay_23_5;
  reg                 io_A_Valid_4_delay_24_4;
  reg                 io_A_Valid_4_delay_25_3;
  reg                 io_A_Valid_4_delay_26_2;
  reg                 io_A_Valid_4_delay_27_1;
  reg                 io_A_Valid_4_delay_28;
  reg                 io_B_Valid_28_delay_1_3;
  reg                 io_B_Valid_28_delay_2_2;
  reg                 io_B_Valid_28_delay_3_1;
  reg                 io_B_Valid_28_delay_4;
  reg                 io_A_Valid_4_delay_1_28;
  reg                 io_A_Valid_4_delay_2_27;
  reg                 io_A_Valid_4_delay_3_26;
  reg                 io_A_Valid_4_delay_4_25;
  reg                 io_A_Valid_4_delay_5_24;
  reg                 io_A_Valid_4_delay_6_23;
  reg                 io_A_Valid_4_delay_7_22;
  reg                 io_A_Valid_4_delay_8_21;
  reg                 io_A_Valid_4_delay_9_20;
  reg                 io_A_Valid_4_delay_10_19;
  reg                 io_A_Valid_4_delay_11_18;
  reg                 io_A_Valid_4_delay_12_17;
  reg                 io_A_Valid_4_delay_13_16;
  reg                 io_A_Valid_4_delay_14_15;
  reg                 io_A_Valid_4_delay_15_14;
  reg                 io_A_Valid_4_delay_16_13;
  reg                 io_A_Valid_4_delay_17_12;
  reg                 io_A_Valid_4_delay_18_11;
  reg                 io_A_Valid_4_delay_19_10;
  reg                 io_A_Valid_4_delay_20_9;
  reg                 io_A_Valid_4_delay_21_8;
  reg                 io_A_Valid_4_delay_22_7;
  reg                 io_A_Valid_4_delay_23_6;
  reg                 io_A_Valid_4_delay_24_5;
  reg                 io_A_Valid_4_delay_25_4;
  reg                 io_A_Valid_4_delay_26_3;
  reg                 io_A_Valid_4_delay_27_2;
  reg                 io_A_Valid_4_delay_28_1;
  reg                 io_A_Valid_4_delay_29;
  reg                 io_B_Valid_29_delay_1_3;
  reg                 io_B_Valid_29_delay_2_2;
  reg                 io_B_Valid_29_delay_3_1;
  reg                 io_B_Valid_29_delay_4;
  reg                 io_A_Valid_4_delay_1_29;
  reg                 io_A_Valid_4_delay_2_28;
  reg                 io_A_Valid_4_delay_3_27;
  reg                 io_A_Valid_4_delay_4_26;
  reg                 io_A_Valid_4_delay_5_25;
  reg                 io_A_Valid_4_delay_6_24;
  reg                 io_A_Valid_4_delay_7_23;
  reg                 io_A_Valid_4_delay_8_22;
  reg                 io_A_Valid_4_delay_9_21;
  reg                 io_A_Valid_4_delay_10_20;
  reg                 io_A_Valid_4_delay_11_19;
  reg                 io_A_Valid_4_delay_12_18;
  reg                 io_A_Valid_4_delay_13_17;
  reg                 io_A_Valid_4_delay_14_16;
  reg                 io_A_Valid_4_delay_15_15;
  reg                 io_A_Valid_4_delay_16_14;
  reg                 io_A_Valid_4_delay_17_13;
  reg                 io_A_Valid_4_delay_18_12;
  reg                 io_A_Valid_4_delay_19_11;
  reg                 io_A_Valid_4_delay_20_10;
  reg                 io_A_Valid_4_delay_21_9;
  reg                 io_A_Valid_4_delay_22_8;
  reg                 io_A_Valid_4_delay_23_7;
  reg                 io_A_Valid_4_delay_24_6;
  reg                 io_A_Valid_4_delay_25_5;
  reg                 io_A_Valid_4_delay_26_4;
  reg                 io_A_Valid_4_delay_27_3;
  reg                 io_A_Valid_4_delay_28_2;
  reg                 io_A_Valid_4_delay_29_1;
  reg                 io_A_Valid_4_delay_30;
  reg                 io_B_Valid_30_delay_1_3;
  reg                 io_B_Valid_30_delay_2_2;
  reg                 io_B_Valid_30_delay_3_1;
  reg                 io_B_Valid_30_delay_4;
  reg                 io_A_Valid_4_delay_1_30;
  reg                 io_A_Valid_4_delay_2_29;
  reg                 io_A_Valid_4_delay_3_28;
  reg                 io_A_Valid_4_delay_4_27;
  reg                 io_A_Valid_4_delay_5_26;
  reg                 io_A_Valid_4_delay_6_25;
  reg                 io_A_Valid_4_delay_7_24;
  reg                 io_A_Valid_4_delay_8_23;
  reg                 io_A_Valid_4_delay_9_22;
  reg                 io_A_Valid_4_delay_10_21;
  reg                 io_A_Valid_4_delay_11_20;
  reg                 io_A_Valid_4_delay_12_19;
  reg                 io_A_Valid_4_delay_13_18;
  reg                 io_A_Valid_4_delay_14_17;
  reg                 io_A_Valid_4_delay_15_16;
  reg                 io_A_Valid_4_delay_16_15;
  reg                 io_A_Valid_4_delay_17_14;
  reg                 io_A_Valid_4_delay_18_13;
  reg                 io_A_Valid_4_delay_19_12;
  reg                 io_A_Valid_4_delay_20_11;
  reg                 io_A_Valid_4_delay_21_10;
  reg                 io_A_Valid_4_delay_22_9;
  reg                 io_A_Valid_4_delay_23_8;
  reg                 io_A_Valid_4_delay_24_7;
  reg                 io_A_Valid_4_delay_25_6;
  reg                 io_A_Valid_4_delay_26_5;
  reg                 io_A_Valid_4_delay_27_4;
  reg                 io_A_Valid_4_delay_28_3;
  reg                 io_A_Valid_4_delay_29_2;
  reg                 io_A_Valid_4_delay_30_1;
  reg                 io_A_Valid_4_delay_31;
  reg                 io_B_Valid_31_delay_1_3;
  reg                 io_B_Valid_31_delay_2_2;
  reg                 io_B_Valid_31_delay_3_1;
  reg                 io_B_Valid_31_delay_4;
  reg                 io_A_Valid_4_delay_1_31;
  reg                 io_A_Valid_4_delay_2_30;
  reg                 io_A_Valid_4_delay_3_29;
  reg                 io_A_Valid_4_delay_4_28;
  reg                 io_A_Valid_4_delay_5_27;
  reg                 io_A_Valid_4_delay_6_26;
  reg                 io_A_Valid_4_delay_7_25;
  reg                 io_A_Valid_4_delay_8_24;
  reg                 io_A_Valid_4_delay_9_23;
  reg                 io_A_Valid_4_delay_10_22;
  reg                 io_A_Valid_4_delay_11_21;
  reg                 io_A_Valid_4_delay_12_20;
  reg                 io_A_Valid_4_delay_13_19;
  reg                 io_A_Valid_4_delay_14_18;
  reg                 io_A_Valid_4_delay_15_17;
  reg                 io_A_Valid_4_delay_16_16;
  reg                 io_A_Valid_4_delay_17_15;
  reg                 io_A_Valid_4_delay_18_14;
  reg                 io_A_Valid_4_delay_19_13;
  reg                 io_A_Valid_4_delay_20_12;
  reg                 io_A_Valid_4_delay_21_11;
  reg                 io_A_Valid_4_delay_22_10;
  reg                 io_A_Valid_4_delay_23_9;
  reg                 io_A_Valid_4_delay_24_8;
  reg                 io_A_Valid_4_delay_25_7;
  reg                 io_A_Valid_4_delay_26_6;
  reg                 io_A_Valid_4_delay_27_5;
  reg                 io_A_Valid_4_delay_28_4;
  reg                 io_A_Valid_4_delay_29_3;
  reg                 io_A_Valid_4_delay_30_2;
  reg                 io_A_Valid_4_delay_31_1;
  reg                 io_A_Valid_4_delay_32;
  reg                 io_B_Valid_32_delay_1_3;
  reg                 io_B_Valid_32_delay_2_2;
  reg                 io_B_Valid_32_delay_3_1;
  reg                 io_B_Valid_32_delay_4;
  reg                 io_A_Valid_4_delay_1_32;
  reg                 io_A_Valid_4_delay_2_31;
  reg                 io_A_Valid_4_delay_3_30;
  reg                 io_A_Valid_4_delay_4_29;
  reg                 io_A_Valid_4_delay_5_28;
  reg                 io_A_Valid_4_delay_6_27;
  reg                 io_A_Valid_4_delay_7_26;
  reg                 io_A_Valid_4_delay_8_25;
  reg                 io_A_Valid_4_delay_9_24;
  reg                 io_A_Valid_4_delay_10_23;
  reg                 io_A_Valid_4_delay_11_22;
  reg                 io_A_Valid_4_delay_12_21;
  reg                 io_A_Valid_4_delay_13_20;
  reg                 io_A_Valid_4_delay_14_19;
  reg                 io_A_Valid_4_delay_15_18;
  reg                 io_A_Valid_4_delay_16_17;
  reg                 io_A_Valid_4_delay_17_16;
  reg                 io_A_Valid_4_delay_18_15;
  reg                 io_A_Valid_4_delay_19_14;
  reg                 io_A_Valid_4_delay_20_13;
  reg                 io_A_Valid_4_delay_21_12;
  reg                 io_A_Valid_4_delay_22_11;
  reg                 io_A_Valid_4_delay_23_10;
  reg                 io_A_Valid_4_delay_24_9;
  reg                 io_A_Valid_4_delay_25_8;
  reg                 io_A_Valid_4_delay_26_7;
  reg                 io_A_Valid_4_delay_27_6;
  reg                 io_A_Valid_4_delay_28_5;
  reg                 io_A_Valid_4_delay_29_4;
  reg                 io_A_Valid_4_delay_30_3;
  reg                 io_A_Valid_4_delay_31_2;
  reg                 io_A_Valid_4_delay_32_1;
  reg                 io_A_Valid_4_delay_33;
  reg                 io_B_Valid_33_delay_1_3;
  reg                 io_B_Valid_33_delay_2_2;
  reg                 io_B_Valid_33_delay_3_1;
  reg                 io_B_Valid_33_delay_4;
  reg                 io_A_Valid_4_delay_1_33;
  reg                 io_A_Valid_4_delay_2_32;
  reg                 io_A_Valid_4_delay_3_31;
  reg                 io_A_Valid_4_delay_4_30;
  reg                 io_A_Valid_4_delay_5_29;
  reg                 io_A_Valid_4_delay_6_28;
  reg                 io_A_Valid_4_delay_7_27;
  reg                 io_A_Valid_4_delay_8_26;
  reg                 io_A_Valid_4_delay_9_25;
  reg                 io_A_Valid_4_delay_10_24;
  reg                 io_A_Valid_4_delay_11_23;
  reg                 io_A_Valid_4_delay_12_22;
  reg                 io_A_Valid_4_delay_13_21;
  reg                 io_A_Valid_4_delay_14_20;
  reg                 io_A_Valid_4_delay_15_19;
  reg                 io_A_Valid_4_delay_16_18;
  reg                 io_A_Valid_4_delay_17_17;
  reg                 io_A_Valid_4_delay_18_16;
  reg                 io_A_Valid_4_delay_19_15;
  reg                 io_A_Valid_4_delay_20_14;
  reg                 io_A_Valid_4_delay_21_13;
  reg                 io_A_Valid_4_delay_22_12;
  reg                 io_A_Valid_4_delay_23_11;
  reg                 io_A_Valid_4_delay_24_10;
  reg                 io_A_Valid_4_delay_25_9;
  reg                 io_A_Valid_4_delay_26_8;
  reg                 io_A_Valid_4_delay_27_7;
  reg                 io_A_Valid_4_delay_28_6;
  reg                 io_A_Valid_4_delay_29_5;
  reg                 io_A_Valid_4_delay_30_4;
  reg                 io_A_Valid_4_delay_31_3;
  reg                 io_A_Valid_4_delay_32_2;
  reg                 io_A_Valid_4_delay_33_1;
  reg                 io_A_Valid_4_delay_34;
  reg                 io_B_Valid_34_delay_1_3;
  reg                 io_B_Valid_34_delay_2_2;
  reg                 io_B_Valid_34_delay_3_1;
  reg                 io_B_Valid_34_delay_4;
  reg                 io_A_Valid_4_delay_1_34;
  reg                 io_A_Valid_4_delay_2_33;
  reg                 io_A_Valid_4_delay_3_32;
  reg                 io_A_Valid_4_delay_4_31;
  reg                 io_A_Valid_4_delay_5_30;
  reg                 io_A_Valid_4_delay_6_29;
  reg                 io_A_Valid_4_delay_7_28;
  reg                 io_A_Valid_4_delay_8_27;
  reg                 io_A_Valid_4_delay_9_26;
  reg                 io_A_Valid_4_delay_10_25;
  reg                 io_A_Valid_4_delay_11_24;
  reg                 io_A_Valid_4_delay_12_23;
  reg                 io_A_Valid_4_delay_13_22;
  reg                 io_A_Valid_4_delay_14_21;
  reg                 io_A_Valid_4_delay_15_20;
  reg                 io_A_Valid_4_delay_16_19;
  reg                 io_A_Valid_4_delay_17_18;
  reg                 io_A_Valid_4_delay_18_17;
  reg                 io_A_Valid_4_delay_19_16;
  reg                 io_A_Valid_4_delay_20_15;
  reg                 io_A_Valid_4_delay_21_14;
  reg                 io_A_Valid_4_delay_22_13;
  reg                 io_A_Valid_4_delay_23_12;
  reg                 io_A_Valid_4_delay_24_11;
  reg                 io_A_Valid_4_delay_25_10;
  reg                 io_A_Valid_4_delay_26_9;
  reg                 io_A_Valid_4_delay_27_8;
  reg                 io_A_Valid_4_delay_28_7;
  reg                 io_A_Valid_4_delay_29_6;
  reg                 io_A_Valid_4_delay_30_5;
  reg                 io_A_Valid_4_delay_31_4;
  reg                 io_A_Valid_4_delay_32_3;
  reg                 io_A_Valid_4_delay_33_2;
  reg                 io_A_Valid_4_delay_34_1;
  reg                 io_A_Valid_4_delay_35;
  reg                 io_B_Valid_35_delay_1_3;
  reg                 io_B_Valid_35_delay_2_2;
  reg                 io_B_Valid_35_delay_3_1;
  reg                 io_B_Valid_35_delay_4;
  reg                 io_A_Valid_4_delay_1_35;
  reg                 io_A_Valid_4_delay_2_34;
  reg                 io_A_Valid_4_delay_3_33;
  reg                 io_A_Valid_4_delay_4_32;
  reg                 io_A_Valid_4_delay_5_31;
  reg                 io_A_Valid_4_delay_6_30;
  reg                 io_A_Valid_4_delay_7_29;
  reg                 io_A_Valid_4_delay_8_28;
  reg                 io_A_Valid_4_delay_9_27;
  reg                 io_A_Valid_4_delay_10_26;
  reg                 io_A_Valid_4_delay_11_25;
  reg                 io_A_Valid_4_delay_12_24;
  reg                 io_A_Valid_4_delay_13_23;
  reg                 io_A_Valid_4_delay_14_22;
  reg                 io_A_Valid_4_delay_15_21;
  reg                 io_A_Valid_4_delay_16_20;
  reg                 io_A_Valid_4_delay_17_19;
  reg                 io_A_Valid_4_delay_18_18;
  reg                 io_A_Valid_4_delay_19_17;
  reg                 io_A_Valid_4_delay_20_16;
  reg                 io_A_Valid_4_delay_21_15;
  reg                 io_A_Valid_4_delay_22_14;
  reg                 io_A_Valid_4_delay_23_13;
  reg                 io_A_Valid_4_delay_24_12;
  reg                 io_A_Valid_4_delay_25_11;
  reg                 io_A_Valid_4_delay_26_10;
  reg                 io_A_Valid_4_delay_27_9;
  reg                 io_A_Valid_4_delay_28_8;
  reg                 io_A_Valid_4_delay_29_7;
  reg                 io_A_Valid_4_delay_30_6;
  reg                 io_A_Valid_4_delay_31_5;
  reg                 io_A_Valid_4_delay_32_4;
  reg                 io_A_Valid_4_delay_33_3;
  reg                 io_A_Valid_4_delay_34_2;
  reg                 io_A_Valid_4_delay_35_1;
  reg                 io_A_Valid_4_delay_36;
  reg                 io_B_Valid_36_delay_1_3;
  reg                 io_B_Valid_36_delay_2_2;
  reg                 io_B_Valid_36_delay_3_1;
  reg                 io_B_Valid_36_delay_4;
  reg                 io_A_Valid_4_delay_1_36;
  reg                 io_A_Valid_4_delay_2_35;
  reg                 io_A_Valid_4_delay_3_34;
  reg                 io_A_Valid_4_delay_4_33;
  reg                 io_A_Valid_4_delay_5_32;
  reg                 io_A_Valid_4_delay_6_31;
  reg                 io_A_Valid_4_delay_7_30;
  reg                 io_A_Valid_4_delay_8_29;
  reg                 io_A_Valid_4_delay_9_28;
  reg                 io_A_Valid_4_delay_10_27;
  reg                 io_A_Valid_4_delay_11_26;
  reg                 io_A_Valid_4_delay_12_25;
  reg                 io_A_Valid_4_delay_13_24;
  reg                 io_A_Valid_4_delay_14_23;
  reg                 io_A_Valid_4_delay_15_22;
  reg                 io_A_Valid_4_delay_16_21;
  reg                 io_A_Valid_4_delay_17_20;
  reg                 io_A_Valid_4_delay_18_19;
  reg                 io_A_Valid_4_delay_19_18;
  reg                 io_A_Valid_4_delay_20_17;
  reg                 io_A_Valid_4_delay_21_16;
  reg                 io_A_Valid_4_delay_22_15;
  reg                 io_A_Valid_4_delay_23_14;
  reg                 io_A_Valid_4_delay_24_13;
  reg                 io_A_Valid_4_delay_25_12;
  reg                 io_A_Valid_4_delay_26_11;
  reg                 io_A_Valid_4_delay_27_10;
  reg                 io_A_Valid_4_delay_28_9;
  reg                 io_A_Valid_4_delay_29_8;
  reg                 io_A_Valid_4_delay_30_7;
  reg                 io_A_Valid_4_delay_31_6;
  reg                 io_A_Valid_4_delay_32_5;
  reg                 io_A_Valid_4_delay_33_4;
  reg                 io_A_Valid_4_delay_34_3;
  reg                 io_A_Valid_4_delay_35_2;
  reg                 io_A_Valid_4_delay_36_1;
  reg                 io_A_Valid_4_delay_37;
  reg                 io_B_Valid_37_delay_1_3;
  reg                 io_B_Valid_37_delay_2_2;
  reg                 io_B_Valid_37_delay_3_1;
  reg                 io_B_Valid_37_delay_4;
  reg                 io_A_Valid_4_delay_1_37;
  reg                 io_A_Valid_4_delay_2_36;
  reg                 io_A_Valid_4_delay_3_35;
  reg                 io_A_Valid_4_delay_4_34;
  reg                 io_A_Valid_4_delay_5_33;
  reg                 io_A_Valid_4_delay_6_32;
  reg                 io_A_Valid_4_delay_7_31;
  reg                 io_A_Valid_4_delay_8_30;
  reg                 io_A_Valid_4_delay_9_29;
  reg                 io_A_Valid_4_delay_10_28;
  reg                 io_A_Valid_4_delay_11_27;
  reg                 io_A_Valid_4_delay_12_26;
  reg                 io_A_Valid_4_delay_13_25;
  reg                 io_A_Valid_4_delay_14_24;
  reg                 io_A_Valid_4_delay_15_23;
  reg                 io_A_Valid_4_delay_16_22;
  reg                 io_A_Valid_4_delay_17_21;
  reg                 io_A_Valid_4_delay_18_20;
  reg                 io_A_Valid_4_delay_19_19;
  reg                 io_A_Valid_4_delay_20_18;
  reg                 io_A_Valid_4_delay_21_17;
  reg                 io_A_Valid_4_delay_22_16;
  reg                 io_A_Valid_4_delay_23_15;
  reg                 io_A_Valid_4_delay_24_14;
  reg                 io_A_Valid_4_delay_25_13;
  reg                 io_A_Valid_4_delay_26_12;
  reg                 io_A_Valid_4_delay_27_11;
  reg                 io_A_Valid_4_delay_28_10;
  reg                 io_A_Valid_4_delay_29_9;
  reg                 io_A_Valid_4_delay_30_8;
  reg                 io_A_Valid_4_delay_31_7;
  reg                 io_A_Valid_4_delay_32_6;
  reg                 io_A_Valid_4_delay_33_5;
  reg                 io_A_Valid_4_delay_34_4;
  reg                 io_A_Valid_4_delay_35_3;
  reg                 io_A_Valid_4_delay_36_2;
  reg                 io_A_Valid_4_delay_37_1;
  reg                 io_A_Valid_4_delay_38;
  reg                 io_B_Valid_38_delay_1_3;
  reg                 io_B_Valid_38_delay_2_2;
  reg                 io_B_Valid_38_delay_3_1;
  reg                 io_B_Valid_38_delay_4;
  reg                 io_A_Valid_4_delay_1_38;
  reg                 io_A_Valid_4_delay_2_37;
  reg                 io_A_Valid_4_delay_3_36;
  reg                 io_A_Valid_4_delay_4_35;
  reg                 io_A_Valid_4_delay_5_34;
  reg                 io_A_Valid_4_delay_6_33;
  reg                 io_A_Valid_4_delay_7_32;
  reg                 io_A_Valid_4_delay_8_31;
  reg                 io_A_Valid_4_delay_9_30;
  reg                 io_A_Valid_4_delay_10_29;
  reg                 io_A_Valid_4_delay_11_28;
  reg                 io_A_Valid_4_delay_12_27;
  reg                 io_A_Valid_4_delay_13_26;
  reg                 io_A_Valid_4_delay_14_25;
  reg                 io_A_Valid_4_delay_15_24;
  reg                 io_A_Valid_4_delay_16_23;
  reg                 io_A_Valid_4_delay_17_22;
  reg                 io_A_Valid_4_delay_18_21;
  reg                 io_A_Valid_4_delay_19_20;
  reg                 io_A_Valid_4_delay_20_19;
  reg                 io_A_Valid_4_delay_21_18;
  reg                 io_A_Valid_4_delay_22_17;
  reg                 io_A_Valid_4_delay_23_16;
  reg                 io_A_Valid_4_delay_24_15;
  reg                 io_A_Valid_4_delay_25_14;
  reg                 io_A_Valid_4_delay_26_13;
  reg                 io_A_Valid_4_delay_27_12;
  reg                 io_A_Valid_4_delay_28_11;
  reg                 io_A_Valid_4_delay_29_10;
  reg                 io_A_Valid_4_delay_30_9;
  reg                 io_A_Valid_4_delay_31_8;
  reg                 io_A_Valid_4_delay_32_7;
  reg                 io_A_Valid_4_delay_33_6;
  reg                 io_A_Valid_4_delay_34_5;
  reg                 io_A_Valid_4_delay_35_4;
  reg                 io_A_Valid_4_delay_36_3;
  reg                 io_A_Valid_4_delay_37_2;
  reg                 io_A_Valid_4_delay_38_1;
  reg                 io_A_Valid_4_delay_39;
  reg                 io_B_Valid_39_delay_1_3;
  reg                 io_B_Valid_39_delay_2_2;
  reg                 io_B_Valid_39_delay_3_1;
  reg                 io_B_Valid_39_delay_4;
  reg                 io_A_Valid_4_delay_1_39;
  reg                 io_A_Valid_4_delay_2_38;
  reg                 io_A_Valid_4_delay_3_37;
  reg                 io_A_Valid_4_delay_4_36;
  reg                 io_A_Valid_4_delay_5_35;
  reg                 io_A_Valid_4_delay_6_34;
  reg                 io_A_Valid_4_delay_7_33;
  reg                 io_A_Valid_4_delay_8_32;
  reg                 io_A_Valid_4_delay_9_31;
  reg                 io_A_Valid_4_delay_10_30;
  reg                 io_A_Valid_4_delay_11_29;
  reg                 io_A_Valid_4_delay_12_28;
  reg                 io_A_Valid_4_delay_13_27;
  reg                 io_A_Valid_4_delay_14_26;
  reg                 io_A_Valid_4_delay_15_25;
  reg                 io_A_Valid_4_delay_16_24;
  reg                 io_A_Valid_4_delay_17_23;
  reg                 io_A_Valid_4_delay_18_22;
  reg                 io_A_Valid_4_delay_19_21;
  reg                 io_A_Valid_4_delay_20_20;
  reg                 io_A_Valid_4_delay_21_19;
  reg                 io_A_Valid_4_delay_22_18;
  reg                 io_A_Valid_4_delay_23_17;
  reg                 io_A_Valid_4_delay_24_16;
  reg                 io_A_Valid_4_delay_25_15;
  reg                 io_A_Valid_4_delay_26_14;
  reg                 io_A_Valid_4_delay_27_13;
  reg                 io_A_Valid_4_delay_28_12;
  reg                 io_A_Valid_4_delay_29_11;
  reg                 io_A_Valid_4_delay_30_10;
  reg                 io_A_Valid_4_delay_31_9;
  reg                 io_A_Valid_4_delay_32_8;
  reg                 io_A_Valid_4_delay_33_7;
  reg                 io_A_Valid_4_delay_34_6;
  reg                 io_A_Valid_4_delay_35_5;
  reg                 io_A_Valid_4_delay_36_4;
  reg                 io_A_Valid_4_delay_37_3;
  reg                 io_A_Valid_4_delay_38_2;
  reg                 io_A_Valid_4_delay_39_1;
  reg                 io_A_Valid_4_delay_40;
  reg                 io_B_Valid_40_delay_1_3;
  reg                 io_B_Valid_40_delay_2_2;
  reg                 io_B_Valid_40_delay_3_1;
  reg                 io_B_Valid_40_delay_4;
  reg                 io_A_Valid_4_delay_1_40;
  reg                 io_A_Valid_4_delay_2_39;
  reg                 io_A_Valid_4_delay_3_38;
  reg                 io_A_Valid_4_delay_4_37;
  reg                 io_A_Valid_4_delay_5_36;
  reg                 io_A_Valid_4_delay_6_35;
  reg                 io_A_Valid_4_delay_7_34;
  reg                 io_A_Valid_4_delay_8_33;
  reg                 io_A_Valid_4_delay_9_32;
  reg                 io_A_Valid_4_delay_10_31;
  reg                 io_A_Valid_4_delay_11_30;
  reg                 io_A_Valid_4_delay_12_29;
  reg                 io_A_Valid_4_delay_13_28;
  reg                 io_A_Valid_4_delay_14_27;
  reg                 io_A_Valid_4_delay_15_26;
  reg                 io_A_Valid_4_delay_16_25;
  reg                 io_A_Valid_4_delay_17_24;
  reg                 io_A_Valid_4_delay_18_23;
  reg                 io_A_Valid_4_delay_19_22;
  reg                 io_A_Valid_4_delay_20_21;
  reg                 io_A_Valid_4_delay_21_20;
  reg                 io_A_Valid_4_delay_22_19;
  reg                 io_A_Valid_4_delay_23_18;
  reg                 io_A_Valid_4_delay_24_17;
  reg                 io_A_Valid_4_delay_25_16;
  reg                 io_A_Valid_4_delay_26_15;
  reg                 io_A_Valid_4_delay_27_14;
  reg                 io_A_Valid_4_delay_28_13;
  reg                 io_A_Valid_4_delay_29_12;
  reg                 io_A_Valid_4_delay_30_11;
  reg                 io_A_Valid_4_delay_31_10;
  reg                 io_A_Valid_4_delay_32_9;
  reg                 io_A_Valid_4_delay_33_8;
  reg                 io_A_Valid_4_delay_34_7;
  reg                 io_A_Valid_4_delay_35_6;
  reg                 io_A_Valid_4_delay_36_5;
  reg                 io_A_Valid_4_delay_37_4;
  reg                 io_A_Valid_4_delay_38_3;
  reg                 io_A_Valid_4_delay_39_2;
  reg                 io_A_Valid_4_delay_40_1;
  reg                 io_A_Valid_4_delay_41;
  reg                 io_B_Valid_41_delay_1_3;
  reg                 io_B_Valid_41_delay_2_2;
  reg                 io_B_Valid_41_delay_3_1;
  reg                 io_B_Valid_41_delay_4;
  reg                 io_A_Valid_4_delay_1_41;
  reg                 io_A_Valid_4_delay_2_40;
  reg                 io_A_Valid_4_delay_3_39;
  reg                 io_A_Valid_4_delay_4_38;
  reg                 io_A_Valid_4_delay_5_37;
  reg                 io_A_Valid_4_delay_6_36;
  reg                 io_A_Valid_4_delay_7_35;
  reg                 io_A_Valid_4_delay_8_34;
  reg                 io_A_Valid_4_delay_9_33;
  reg                 io_A_Valid_4_delay_10_32;
  reg                 io_A_Valid_4_delay_11_31;
  reg                 io_A_Valid_4_delay_12_30;
  reg                 io_A_Valid_4_delay_13_29;
  reg                 io_A_Valid_4_delay_14_28;
  reg                 io_A_Valid_4_delay_15_27;
  reg                 io_A_Valid_4_delay_16_26;
  reg                 io_A_Valid_4_delay_17_25;
  reg                 io_A_Valid_4_delay_18_24;
  reg                 io_A_Valid_4_delay_19_23;
  reg                 io_A_Valid_4_delay_20_22;
  reg                 io_A_Valid_4_delay_21_21;
  reg                 io_A_Valid_4_delay_22_20;
  reg                 io_A_Valid_4_delay_23_19;
  reg                 io_A_Valid_4_delay_24_18;
  reg                 io_A_Valid_4_delay_25_17;
  reg                 io_A_Valid_4_delay_26_16;
  reg                 io_A_Valid_4_delay_27_15;
  reg                 io_A_Valid_4_delay_28_14;
  reg                 io_A_Valid_4_delay_29_13;
  reg                 io_A_Valid_4_delay_30_12;
  reg                 io_A_Valid_4_delay_31_11;
  reg                 io_A_Valid_4_delay_32_10;
  reg                 io_A_Valid_4_delay_33_9;
  reg                 io_A_Valid_4_delay_34_8;
  reg                 io_A_Valid_4_delay_35_7;
  reg                 io_A_Valid_4_delay_36_6;
  reg                 io_A_Valid_4_delay_37_5;
  reg                 io_A_Valid_4_delay_38_4;
  reg                 io_A_Valid_4_delay_39_3;
  reg                 io_A_Valid_4_delay_40_2;
  reg                 io_A_Valid_4_delay_41_1;
  reg                 io_A_Valid_4_delay_42;
  reg                 io_B_Valid_42_delay_1_3;
  reg                 io_B_Valid_42_delay_2_2;
  reg                 io_B_Valid_42_delay_3_1;
  reg                 io_B_Valid_42_delay_4;
  reg                 io_A_Valid_4_delay_1_42;
  reg                 io_A_Valid_4_delay_2_41;
  reg                 io_A_Valid_4_delay_3_40;
  reg                 io_A_Valid_4_delay_4_39;
  reg                 io_A_Valid_4_delay_5_38;
  reg                 io_A_Valid_4_delay_6_37;
  reg                 io_A_Valid_4_delay_7_36;
  reg                 io_A_Valid_4_delay_8_35;
  reg                 io_A_Valid_4_delay_9_34;
  reg                 io_A_Valid_4_delay_10_33;
  reg                 io_A_Valid_4_delay_11_32;
  reg                 io_A_Valid_4_delay_12_31;
  reg                 io_A_Valid_4_delay_13_30;
  reg                 io_A_Valid_4_delay_14_29;
  reg                 io_A_Valid_4_delay_15_28;
  reg                 io_A_Valid_4_delay_16_27;
  reg                 io_A_Valid_4_delay_17_26;
  reg                 io_A_Valid_4_delay_18_25;
  reg                 io_A_Valid_4_delay_19_24;
  reg                 io_A_Valid_4_delay_20_23;
  reg                 io_A_Valid_4_delay_21_22;
  reg                 io_A_Valid_4_delay_22_21;
  reg                 io_A_Valid_4_delay_23_20;
  reg                 io_A_Valid_4_delay_24_19;
  reg                 io_A_Valid_4_delay_25_18;
  reg                 io_A_Valid_4_delay_26_17;
  reg                 io_A_Valid_4_delay_27_16;
  reg                 io_A_Valid_4_delay_28_15;
  reg                 io_A_Valid_4_delay_29_14;
  reg                 io_A_Valid_4_delay_30_13;
  reg                 io_A_Valid_4_delay_31_12;
  reg                 io_A_Valid_4_delay_32_11;
  reg                 io_A_Valid_4_delay_33_10;
  reg                 io_A_Valid_4_delay_34_9;
  reg                 io_A_Valid_4_delay_35_8;
  reg                 io_A_Valid_4_delay_36_7;
  reg                 io_A_Valid_4_delay_37_6;
  reg                 io_A_Valid_4_delay_38_5;
  reg                 io_A_Valid_4_delay_39_4;
  reg                 io_A_Valid_4_delay_40_3;
  reg                 io_A_Valid_4_delay_41_2;
  reg                 io_A_Valid_4_delay_42_1;
  reg                 io_A_Valid_4_delay_43;
  reg                 io_B_Valid_43_delay_1_3;
  reg                 io_B_Valid_43_delay_2_2;
  reg                 io_B_Valid_43_delay_3_1;
  reg                 io_B_Valid_43_delay_4;
  reg                 io_A_Valid_4_delay_1_43;
  reg                 io_A_Valid_4_delay_2_42;
  reg                 io_A_Valid_4_delay_3_41;
  reg                 io_A_Valid_4_delay_4_40;
  reg                 io_A_Valid_4_delay_5_39;
  reg                 io_A_Valid_4_delay_6_38;
  reg                 io_A_Valid_4_delay_7_37;
  reg                 io_A_Valid_4_delay_8_36;
  reg                 io_A_Valid_4_delay_9_35;
  reg                 io_A_Valid_4_delay_10_34;
  reg                 io_A_Valid_4_delay_11_33;
  reg                 io_A_Valid_4_delay_12_32;
  reg                 io_A_Valid_4_delay_13_31;
  reg                 io_A_Valid_4_delay_14_30;
  reg                 io_A_Valid_4_delay_15_29;
  reg                 io_A_Valid_4_delay_16_28;
  reg                 io_A_Valid_4_delay_17_27;
  reg                 io_A_Valid_4_delay_18_26;
  reg                 io_A_Valid_4_delay_19_25;
  reg                 io_A_Valid_4_delay_20_24;
  reg                 io_A_Valid_4_delay_21_23;
  reg                 io_A_Valid_4_delay_22_22;
  reg                 io_A_Valid_4_delay_23_21;
  reg                 io_A_Valid_4_delay_24_20;
  reg                 io_A_Valid_4_delay_25_19;
  reg                 io_A_Valid_4_delay_26_18;
  reg                 io_A_Valid_4_delay_27_17;
  reg                 io_A_Valid_4_delay_28_16;
  reg                 io_A_Valid_4_delay_29_15;
  reg                 io_A_Valid_4_delay_30_14;
  reg                 io_A_Valid_4_delay_31_13;
  reg                 io_A_Valid_4_delay_32_12;
  reg                 io_A_Valid_4_delay_33_11;
  reg                 io_A_Valid_4_delay_34_10;
  reg                 io_A_Valid_4_delay_35_9;
  reg                 io_A_Valid_4_delay_36_8;
  reg                 io_A_Valid_4_delay_37_7;
  reg                 io_A_Valid_4_delay_38_6;
  reg                 io_A_Valid_4_delay_39_5;
  reg                 io_A_Valid_4_delay_40_4;
  reg                 io_A_Valid_4_delay_41_3;
  reg                 io_A_Valid_4_delay_42_2;
  reg                 io_A_Valid_4_delay_43_1;
  reg                 io_A_Valid_4_delay_44;
  reg                 io_B_Valid_44_delay_1_3;
  reg                 io_B_Valid_44_delay_2_2;
  reg                 io_B_Valid_44_delay_3_1;
  reg                 io_B_Valid_44_delay_4;
  reg                 io_A_Valid_4_delay_1_44;
  reg                 io_A_Valid_4_delay_2_43;
  reg                 io_A_Valid_4_delay_3_42;
  reg                 io_A_Valid_4_delay_4_41;
  reg                 io_A_Valid_4_delay_5_40;
  reg                 io_A_Valid_4_delay_6_39;
  reg                 io_A_Valid_4_delay_7_38;
  reg                 io_A_Valid_4_delay_8_37;
  reg                 io_A_Valid_4_delay_9_36;
  reg                 io_A_Valid_4_delay_10_35;
  reg                 io_A_Valid_4_delay_11_34;
  reg                 io_A_Valid_4_delay_12_33;
  reg                 io_A_Valid_4_delay_13_32;
  reg                 io_A_Valid_4_delay_14_31;
  reg                 io_A_Valid_4_delay_15_30;
  reg                 io_A_Valid_4_delay_16_29;
  reg                 io_A_Valid_4_delay_17_28;
  reg                 io_A_Valid_4_delay_18_27;
  reg                 io_A_Valid_4_delay_19_26;
  reg                 io_A_Valid_4_delay_20_25;
  reg                 io_A_Valid_4_delay_21_24;
  reg                 io_A_Valid_4_delay_22_23;
  reg                 io_A_Valid_4_delay_23_22;
  reg                 io_A_Valid_4_delay_24_21;
  reg                 io_A_Valid_4_delay_25_20;
  reg                 io_A_Valid_4_delay_26_19;
  reg                 io_A_Valid_4_delay_27_18;
  reg                 io_A_Valid_4_delay_28_17;
  reg                 io_A_Valid_4_delay_29_16;
  reg                 io_A_Valid_4_delay_30_15;
  reg                 io_A_Valid_4_delay_31_14;
  reg                 io_A_Valid_4_delay_32_13;
  reg                 io_A_Valid_4_delay_33_12;
  reg                 io_A_Valid_4_delay_34_11;
  reg                 io_A_Valid_4_delay_35_10;
  reg                 io_A_Valid_4_delay_36_9;
  reg                 io_A_Valid_4_delay_37_8;
  reg                 io_A_Valid_4_delay_38_7;
  reg                 io_A_Valid_4_delay_39_6;
  reg                 io_A_Valid_4_delay_40_5;
  reg                 io_A_Valid_4_delay_41_4;
  reg                 io_A_Valid_4_delay_42_3;
  reg                 io_A_Valid_4_delay_43_2;
  reg                 io_A_Valid_4_delay_44_1;
  reg                 io_A_Valid_4_delay_45;
  reg                 io_B_Valid_45_delay_1_3;
  reg                 io_B_Valid_45_delay_2_2;
  reg                 io_B_Valid_45_delay_3_1;
  reg                 io_B_Valid_45_delay_4;
  reg                 io_A_Valid_4_delay_1_45;
  reg                 io_A_Valid_4_delay_2_44;
  reg                 io_A_Valid_4_delay_3_43;
  reg                 io_A_Valid_4_delay_4_42;
  reg                 io_A_Valid_4_delay_5_41;
  reg                 io_A_Valid_4_delay_6_40;
  reg                 io_A_Valid_4_delay_7_39;
  reg                 io_A_Valid_4_delay_8_38;
  reg                 io_A_Valid_4_delay_9_37;
  reg                 io_A_Valid_4_delay_10_36;
  reg                 io_A_Valid_4_delay_11_35;
  reg                 io_A_Valid_4_delay_12_34;
  reg                 io_A_Valid_4_delay_13_33;
  reg                 io_A_Valid_4_delay_14_32;
  reg                 io_A_Valid_4_delay_15_31;
  reg                 io_A_Valid_4_delay_16_30;
  reg                 io_A_Valid_4_delay_17_29;
  reg                 io_A_Valid_4_delay_18_28;
  reg                 io_A_Valid_4_delay_19_27;
  reg                 io_A_Valid_4_delay_20_26;
  reg                 io_A_Valid_4_delay_21_25;
  reg                 io_A_Valid_4_delay_22_24;
  reg                 io_A_Valid_4_delay_23_23;
  reg                 io_A_Valid_4_delay_24_22;
  reg                 io_A_Valid_4_delay_25_21;
  reg                 io_A_Valid_4_delay_26_20;
  reg                 io_A_Valid_4_delay_27_19;
  reg                 io_A_Valid_4_delay_28_18;
  reg                 io_A_Valid_4_delay_29_17;
  reg                 io_A_Valid_4_delay_30_16;
  reg                 io_A_Valid_4_delay_31_15;
  reg                 io_A_Valid_4_delay_32_14;
  reg                 io_A_Valid_4_delay_33_13;
  reg                 io_A_Valid_4_delay_34_12;
  reg                 io_A_Valid_4_delay_35_11;
  reg                 io_A_Valid_4_delay_36_10;
  reg                 io_A_Valid_4_delay_37_9;
  reg                 io_A_Valid_4_delay_38_8;
  reg                 io_A_Valid_4_delay_39_7;
  reg                 io_A_Valid_4_delay_40_6;
  reg                 io_A_Valid_4_delay_41_5;
  reg                 io_A_Valid_4_delay_42_4;
  reg                 io_A_Valid_4_delay_43_3;
  reg                 io_A_Valid_4_delay_44_2;
  reg                 io_A_Valid_4_delay_45_1;
  reg                 io_A_Valid_4_delay_46;
  reg                 io_B_Valid_46_delay_1_3;
  reg                 io_B_Valid_46_delay_2_2;
  reg                 io_B_Valid_46_delay_3_1;
  reg                 io_B_Valid_46_delay_4;
  reg                 io_A_Valid_4_delay_1_46;
  reg                 io_A_Valid_4_delay_2_45;
  reg                 io_A_Valid_4_delay_3_44;
  reg                 io_A_Valid_4_delay_4_43;
  reg                 io_A_Valid_4_delay_5_42;
  reg                 io_A_Valid_4_delay_6_41;
  reg                 io_A_Valid_4_delay_7_40;
  reg                 io_A_Valid_4_delay_8_39;
  reg                 io_A_Valid_4_delay_9_38;
  reg                 io_A_Valid_4_delay_10_37;
  reg                 io_A_Valid_4_delay_11_36;
  reg                 io_A_Valid_4_delay_12_35;
  reg                 io_A_Valid_4_delay_13_34;
  reg                 io_A_Valid_4_delay_14_33;
  reg                 io_A_Valid_4_delay_15_32;
  reg                 io_A_Valid_4_delay_16_31;
  reg                 io_A_Valid_4_delay_17_30;
  reg                 io_A_Valid_4_delay_18_29;
  reg                 io_A_Valid_4_delay_19_28;
  reg                 io_A_Valid_4_delay_20_27;
  reg                 io_A_Valid_4_delay_21_26;
  reg                 io_A_Valid_4_delay_22_25;
  reg                 io_A_Valid_4_delay_23_24;
  reg                 io_A_Valid_4_delay_24_23;
  reg                 io_A_Valid_4_delay_25_22;
  reg                 io_A_Valid_4_delay_26_21;
  reg                 io_A_Valid_4_delay_27_20;
  reg                 io_A_Valid_4_delay_28_19;
  reg                 io_A_Valid_4_delay_29_18;
  reg                 io_A_Valid_4_delay_30_17;
  reg                 io_A_Valid_4_delay_31_16;
  reg                 io_A_Valid_4_delay_32_15;
  reg                 io_A_Valid_4_delay_33_14;
  reg                 io_A_Valid_4_delay_34_13;
  reg                 io_A_Valid_4_delay_35_12;
  reg                 io_A_Valid_4_delay_36_11;
  reg                 io_A_Valid_4_delay_37_10;
  reg                 io_A_Valid_4_delay_38_9;
  reg                 io_A_Valid_4_delay_39_8;
  reg                 io_A_Valid_4_delay_40_7;
  reg                 io_A_Valid_4_delay_41_6;
  reg                 io_A_Valid_4_delay_42_5;
  reg                 io_A_Valid_4_delay_43_4;
  reg                 io_A_Valid_4_delay_44_3;
  reg                 io_A_Valid_4_delay_45_2;
  reg                 io_A_Valid_4_delay_46_1;
  reg                 io_A_Valid_4_delay_47;
  reg                 io_B_Valid_47_delay_1_3;
  reg                 io_B_Valid_47_delay_2_2;
  reg                 io_B_Valid_47_delay_3_1;
  reg                 io_B_Valid_47_delay_4;
  reg                 io_A_Valid_4_delay_1_47;
  reg                 io_A_Valid_4_delay_2_46;
  reg                 io_A_Valid_4_delay_3_45;
  reg                 io_A_Valid_4_delay_4_44;
  reg                 io_A_Valid_4_delay_5_43;
  reg                 io_A_Valid_4_delay_6_42;
  reg                 io_A_Valid_4_delay_7_41;
  reg                 io_A_Valid_4_delay_8_40;
  reg                 io_A_Valid_4_delay_9_39;
  reg                 io_A_Valid_4_delay_10_38;
  reg                 io_A_Valid_4_delay_11_37;
  reg                 io_A_Valid_4_delay_12_36;
  reg                 io_A_Valid_4_delay_13_35;
  reg                 io_A_Valid_4_delay_14_34;
  reg                 io_A_Valid_4_delay_15_33;
  reg                 io_A_Valid_4_delay_16_32;
  reg                 io_A_Valid_4_delay_17_31;
  reg                 io_A_Valid_4_delay_18_30;
  reg                 io_A_Valid_4_delay_19_29;
  reg                 io_A_Valid_4_delay_20_28;
  reg                 io_A_Valid_4_delay_21_27;
  reg                 io_A_Valid_4_delay_22_26;
  reg                 io_A_Valid_4_delay_23_25;
  reg                 io_A_Valid_4_delay_24_24;
  reg                 io_A_Valid_4_delay_25_23;
  reg                 io_A_Valid_4_delay_26_22;
  reg                 io_A_Valid_4_delay_27_21;
  reg                 io_A_Valid_4_delay_28_20;
  reg                 io_A_Valid_4_delay_29_19;
  reg                 io_A_Valid_4_delay_30_18;
  reg                 io_A_Valid_4_delay_31_17;
  reg                 io_A_Valid_4_delay_32_16;
  reg                 io_A_Valid_4_delay_33_15;
  reg                 io_A_Valid_4_delay_34_14;
  reg                 io_A_Valid_4_delay_35_13;
  reg                 io_A_Valid_4_delay_36_12;
  reg                 io_A_Valid_4_delay_37_11;
  reg                 io_A_Valid_4_delay_38_10;
  reg                 io_A_Valid_4_delay_39_9;
  reg                 io_A_Valid_4_delay_40_8;
  reg                 io_A_Valid_4_delay_41_7;
  reg                 io_A_Valid_4_delay_42_6;
  reg                 io_A_Valid_4_delay_43_5;
  reg                 io_A_Valid_4_delay_44_4;
  reg                 io_A_Valid_4_delay_45_3;
  reg                 io_A_Valid_4_delay_46_2;
  reg                 io_A_Valid_4_delay_47_1;
  reg                 io_A_Valid_4_delay_48;
  reg                 io_B_Valid_48_delay_1_3;
  reg                 io_B_Valid_48_delay_2_2;
  reg                 io_B_Valid_48_delay_3_1;
  reg                 io_B_Valid_48_delay_4;
  reg                 io_A_Valid_4_delay_1_48;
  reg                 io_A_Valid_4_delay_2_47;
  reg                 io_A_Valid_4_delay_3_46;
  reg                 io_A_Valid_4_delay_4_45;
  reg                 io_A_Valid_4_delay_5_44;
  reg                 io_A_Valid_4_delay_6_43;
  reg                 io_A_Valid_4_delay_7_42;
  reg                 io_A_Valid_4_delay_8_41;
  reg                 io_A_Valid_4_delay_9_40;
  reg                 io_A_Valid_4_delay_10_39;
  reg                 io_A_Valid_4_delay_11_38;
  reg                 io_A_Valid_4_delay_12_37;
  reg                 io_A_Valid_4_delay_13_36;
  reg                 io_A_Valid_4_delay_14_35;
  reg                 io_A_Valid_4_delay_15_34;
  reg                 io_A_Valid_4_delay_16_33;
  reg                 io_A_Valid_4_delay_17_32;
  reg                 io_A_Valid_4_delay_18_31;
  reg                 io_A_Valid_4_delay_19_30;
  reg                 io_A_Valid_4_delay_20_29;
  reg                 io_A_Valid_4_delay_21_28;
  reg                 io_A_Valid_4_delay_22_27;
  reg                 io_A_Valid_4_delay_23_26;
  reg                 io_A_Valid_4_delay_24_25;
  reg                 io_A_Valid_4_delay_25_24;
  reg                 io_A_Valid_4_delay_26_23;
  reg                 io_A_Valid_4_delay_27_22;
  reg                 io_A_Valid_4_delay_28_21;
  reg                 io_A_Valid_4_delay_29_20;
  reg                 io_A_Valid_4_delay_30_19;
  reg                 io_A_Valid_4_delay_31_18;
  reg                 io_A_Valid_4_delay_32_17;
  reg                 io_A_Valid_4_delay_33_16;
  reg                 io_A_Valid_4_delay_34_15;
  reg                 io_A_Valid_4_delay_35_14;
  reg                 io_A_Valid_4_delay_36_13;
  reg                 io_A_Valid_4_delay_37_12;
  reg                 io_A_Valid_4_delay_38_11;
  reg                 io_A_Valid_4_delay_39_10;
  reg                 io_A_Valid_4_delay_40_9;
  reg                 io_A_Valid_4_delay_41_8;
  reg                 io_A_Valid_4_delay_42_7;
  reg                 io_A_Valid_4_delay_43_6;
  reg                 io_A_Valid_4_delay_44_5;
  reg                 io_A_Valid_4_delay_45_4;
  reg                 io_A_Valid_4_delay_46_3;
  reg                 io_A_Valid_4_delay_47_2;
  reg                 io_A_Valid_4_delay_48_1;
  reg                 io_A_Valid_4_delay_49;
  reg                 io_B_Valid_49_delay_1_3;
  reg                 io_B_Valid_49_delay_2_2;
  reg                 io_B_Valid_49_delay_3_1;
  reg                 io_B_Valid_49_delay_4;
  reg                 io_A_Valid_4_delay_1_49;
  reg                 io_A_Valid_4_delay_2_48;
  reg                 io_A_Valid_4_delay_3_47;
  reg                 io_A_Valid_4_delay_4_46;
  reg                 io_A_Valid_4_delay_5_45;
  reg                 io_A_Valid_4_delay_6_44;
  reg                 io_A_Valid_4_delay_7_43;
  reg                 io_A_Valid_4_delay_8_42;
  reg                 io_A_Valid_4_delay_9_41;
  reg                 io_A_Valid_4_delay_10_40;
  reg                 io_A_Valid_4_delay_11_39;
  reg                 io_A_Valid_4_delay_12_38;
  reg                 io_A_Valid_4_delay_13_37;
  reg                 io_A_Valid_4_delay_14_36;
  reg                 io_A_Valid_4_delay_15_35;
  reg                 io_A_Valid_4_delay_16_34;
  reg                 io_A_Valid_4_delay_17_33;
  reg                 io_A_Valid_4_delay_18_32;
  reg                 io_A_Valid_4_delay_19_31;
  reg                 io_A_Valid_4_delay_20_30;
  reg                 io_A_Valid_4_delay_21_29;
  reg                 io_A_Valid_4_delay_22_28;
  reg                 io_A_Valid_4_delay_23_27;
  reg                 io_A_Valid_4_delay_24_26;
  reg                 io_A_Valid_4_delay_25_25;
  reg                 io_A_Valid_4_delay_26_24;
  reg                 io_A_Valid_4_delay_27_23;
  reg                 io_A_Valid_4_delay_28_22;
  reg                 io_A_Valid_4_delay_29_21;
  reg                 io_A_Valid_4_delay_30_20;
  reg                 io_A_Valid_4_delay_31_19;
  reg                 io_A_Valid_4_delay_32_18;
  reg                 io_A_Valid_4_delay_33_17;
  reg                 io_A_Valid_4_delay_34_16;
  reg                 io_A_Valid_4_delay_35_15;
  reg                 io_A_Valid_4_delay_36_14;
  reg                 io_A_Valid_4_delay_37_13;
  reg                 io_A_Valid_4_delay_38_12;
  reg                 io_A_Valid_4_delay_39_11;
  reg                 io_A_Valid_4_delay_40_10;
  reg                 io_A_Valid_4_delay_41_9;
  reg                 io_A_Valid_4_delay_42_8;
  reg                 io_A_Valid_4_delay_43_7;
  reg                 io_A_Valid_4_delay_44_6;
  reg                 io_A_Valid_4_delay_45_5;
  reg                 io_A_Valid_4_delay_46_4;
  reg                 io_A_Valid_4_delay_47_3;
  reg                 io_A_Valid_4_delay_48_2;
  reg                 io_A_Valid_4_delay_49_1;
  reg                 io_A_Valid_4_delay_50;
  reg                 io_B_Valid_50_delay_1_3;
  reg                 io_B_Valid_50_delay_2_2;
  reg                 io_B_Valid_50_delay_3_1;
  reg                 io_B_Valid_50_delay_4;
  reg                 io_A_Valid_4_delay_1_50;
  reg                 io_A_Valid_4_delay_2_49;
  reg                 io_A_Valid_4_delay_3_48;
  reg                 io_A_Valid_4_delay_4_47;
  reg                 io_A_Valid_4_delay_5_46;
  reg                 io_A_Valid_4_delay_6_45;
  reg                 io_A_Valid_4_delay_7_44;
  reg                 io_A_Valid_4_delay_8_43;
  reg                 io_A_Valid_4_delay_9_42;
  reg                 io_A_Valid_4_delay_10_41;
  reg                 io_A_Valid_4_delay_11_40;
  reg                 io_A_Valid_4_delay_12_39;
  reg                 io_A_Valid_4_delay_13_38;
  reg                 io_A_Valid_4_delay_14_37;
  reg                 io_A_Valid_4_delay_15_36;
  reg                 io_A_Valid_4_delay_16_35;
  reg                 io_A_Valid_4_delay_17_34;
  reg                 io_A_Valid_4_delay_18_33;
  reg                 io_A_Valid_4_delay_19_32;
  reg                 io_A_Valid_4_delay_20_31;
  reg                 io_A_Valid_4_delay_21_30;
  reg                 io_A_Valid_4_delay_22_29;
  reg                 io_A_Valid_4_delay_23_28;
  reg                 io_A_Valid_4_delay_24_27;
  reg                 io_A_Valid_4_delay_25_26;
  reg                 io_A_Valid_4_delay_26_25;
  reg                 io_A_Valid_4_delay_27_24;
  reg                 io_A_Valid_4_delay_28_23;
  reg                 io_A_Valid_4_delay_29_22;
  reg                 io_A_Valid_4_delay_30_21;
  reg                 io_A_Valid_4_delay_31_20;
  reg                 io_A_Valid_4_delay_32_19;
  reg                 io_A_Valid_4_delay_33_18;
  reg                 io_A_Valid_4_delay_34_17;
  reg                 io_A_Valid_4_delay_35_16;
  reg                 io_A_Valid_4_delay_36_15;
  reg                 io_A_Valid_4_delay_37_14;
  reg                 io_A_Valid_4_delay_38_13;
  reg                 io_A_Valid_4_delay_39_12;
  reg                 io_A_Valid_4_delay_40_11;
  reg                 io_A_Valid_4_delay_41_10;
  reg                 io_A_Valid_4_delay_42_9;
  reg                 io_A_Valid_4_delay_43_8;
  reg                 io_A_Valid_4_delay_44_7;
  reg                 io_A_Valid_4_delay_45_6;
  reg                 io_A_Valid_4_delay_46_5;
  reg                 io_A_Valid_4_delay_47_4;
  reg                 io_A_Valid_4_delay_48_3;
  reg                 io_A_Valid_4_delay_49_2;
  reg                 io_A_Valid_4_delay_50_1;
  reg                 io_A_Valid_4_delay_51;
  reg                 io_B_Valid_51_delay_1_3;
  reg                 io_B_Valid_51_delay_2_2;
  reg                 io_B_Valid_51_delay_3_1;
  reg                 io_B_Valid_51_delay_4;
  reg                 io_A_Valid_4_delay_1_51;
  reg                 io_A_Valid_4_delay_2_50;
  reg                 io_A_Valid_4_delay_3_49;
  reg                 io_A_Valid_4_delay_4_48;
  reg                 io_A_Valid_4_delay_5_47;
  reg                 io_A_Valid_4_delay_6_46;
  reg                 io_A_Valid_4_delay_7_45;
  reg                 io_A_Valid_4_delay_8_44;
  reg                 io_A_Valid_4_delay_9_43;
  reg                 io_A_Valid_4_delay_10_42;
  reg                 io_A_Valid_4_delay_11_41;
  reg                 io_A_Valid_4_delay_12_40;
  reg                 io_A_Valid_4_delay_13_39;
  reg                 io_A_Valid_4_delay_14_38;
  reg                 io_A_Valid_4_delay_15_37;
  reg                 io_A_Valid_4_delay_16_36;
  reg                 io_A_Valid_4_delay_17_35;
  reg                 io_A_Valid_4_delay_18_34;
  reg                 io_A_Valid_4_delay_19_33;
  reg                 io_A_Valid_4_delay_20_32;
  reg                 io_A_Valid_4_delay_21_31;
  reg                 io_A_Valid_4_delay_22_30;
  reg                 io_A_Valid_4_delay_23_29;
  reg                 io_A_Valid_4_delay_24_28;
  reg                 io_A_Valid_4_delay_25_27;
  reg                 io_A_Valid_4_delay_26_26;
  reg                 io_A_Valid_4_delay_27_25;
  reg                 io_A_Valid_4_delay_28_24;
  reg                 io_A_Valid_4_delay_29_23;
  reg                 io_A_Valid_4_delay_30_22;
  reg                 io_A_Valid_4_delay_31_21;
  reg                 io_A_Valid_4_delay_32_20;
  reg                 io_A_Valid_4_delay_33_19;
  reg                 io_A_Valid_4_delay_34_18;
  reg                 io_A_Valid_4_delay_35_17;
  reg                 io_A_Valid_4_delay_36_16;
  reg                 io_A_Valid_4_delay_37_15;
  reg                 io_A_Valid_4_delay_38_14;
  reg                 io_A_Valid_4_delay_39_13;
  reg                 io_A_Valid_4_delay_40_12;
  reg                 io_A_Valid_4_delay_41_11;
  reg                 io_A_Valid_4_delay_42_10;
  reg                 io_A_Valid_4_delay_43_9;
  reg                 io_A_Valid_4_delay_44_8;
  reg                 io_A_Valid_4_delay_45_7;
  reg                 io_A_Valid_4_delay_46_6;
  reg                 io_A_Valid_4_delay_47_5;
  reg                 io_A_Valid_4_delay_48_4;
  reg                 io_A_Valid_4_delay_49_3;
  reg                 io_A_Valid_4_delay_50_2;
  reg                 io_A_Valid_4_delay_51_1;
  reg                 io_A_Valid_4_delay_52;
  reg                 io_B_Valid_52_delay_1_3;
  reg                 io_B_Valid_52_delay_2_2;
  reg                 io_B_Valid_52_delay_3_1;
  reg                 io_B_Valid_52_delay_4;
  reg                 io_A_Valid_4_delay_1_52;
  reg                 io_A_Valid_4_delay_2_51;
  reg                 io_A_Valid_4_delay_3_50;
  reg                 io_A_Valid_4_delay_4_49;
  reg                 io_A_Valid_4_delay_5_48;
  reg                 io_A_Valid_4_delay_6_47;
  reg                 io_A_Valid_4_delay_7_46;
  reg                 io_A_Valid_4_delay_8_45;
  reg                 io_A_Valid_4_delay_9_44;
  reg                 io_A_Valid_4_delay_10_43;
  reg                 io_A_Valid_4_delay_11_42;
  reg                 io_A_Valid_4_delay_12_41;
  reg                 io_A_Valid_4_delay_13_40;
  reg                 io_A_Valid_4_delay_14_39;
  reg                 io_A_Valid_4_delay_15_38;
  reg                 io_A_Valid_4_delay_16_37;
  reg                 io_A_Valid_4_delay_17_36;
  reg                 io_A_Valid_4_delay_18_35;
  reg                 io_A_Valid_4_delay_19_34;
  reg                 io_A_Valid_4_delay_20_33;
  reg                 io_A_Valid_4_delay_21_32;
  reg                 io_A_Valid_4_delay_22_31;
  reg                 io_A_Valid_4_delay_23_30;
  reg                 io_A_Valid_4_delay_24_29;
  reg                 io_A_Valid_4_delay_25_28;
  reg                 io_A_Valid_4_delay_26_27;
  reg                 io_A_Valid_4_delay_27_26;
  reg                 io_A_Valid_4_delay_28_25;
  reg                 io_A_Valid_4_delay_29_24;
  reg                 io_A_Valid_4_delay_30_23;
  reg                 io_A_Valid_4_delay_31_22;
  reg                 io_A_Valid_4_delay_32_21;
  reg                 io_A_Valid_4_delay_33_20;
  reg                 io_A_Valid_4_delay_34_19;
  reg                 io_A_Valid_4_delay_35_18;
  reg                 io_A_Valid_4_delay_36_17;
  reg                 io_A_Valid_4_delay_37_16;
  reg                 io_A_Valid_4_delay_38_15;
  reg                 io_A_Valid_4_delay_39_14;
  reg                 io_A_Valid_4_delay_40_13;
  reg                 io_A_Valid_4_delay_41_12;
  reg                 io_A_Valid_4_delay_42_11;
  reg                 io_A_Valid_4_delay_43_10;
  reg                 io_A_Valid_4_delay_44_9;
  reg                 io_A_Valid_4_delay_45_8;
  reg                 io_A_Valid_4_delay_46_7;
  reg                 io_A_Valid_4_delay_47_6;
  reg                 io_A_Valid_4_delay_48_5;
  reg                 io_A_Valid_4_delay_49_4;
  reg                 io_A_Valid_4_delay_50_3;
  reg                 io_A_Valid_4_delay_51_2;
  reg                 io_A_Valid_4_delay_52_1;
  reg                 io_A_Valid_4_delay_53;
  reg                 io_B_Valid_53_delay_1_3;
  reg                 io_B_Valid_53_delay_2_2;
  reg                 io_B_Valid_53_delay_3_1;
  reg                 io_B_Valid_53_delay_4;
  reg                 io_A_Valid_4_delay_1_53;
  reg                 io_A_Valid_4_delay_2_52;
  reg                 io_A_Valid_4_delay_3_51;
  reg                 io_A_Valid_4_delay_4_50;
  reg                 io_A_Valid_4_delay_5_49;
  reg                 io_A_Valid_4_delay_6_48;
  reg                 io_A_Valid_4_delay_7_47;
  reg                 io_A_Valid_4_delay_8_46;
  reg                 io_A_Valid_4_delay_9_45;
  reg                 io_A_Valid_4_delay_10_44;
  reg                 io_A_Valid_4_delay_11_43;
  reg                 io_A_Valid_4_delay_12_42;
  reg                 io_A_Valid_4_delay_13_41;
  reg                 io_A_Valid_4_delay_14_40;
  reg                 io_A_Valid_4_delay_15_39;
  reg                 io_A_Valid_4_delay_16_38;
  reg                 io_A_Valid_4_delay_17_37;
  reg                 io_A_Valid_4_delay_18_36;
  reg                 io_A_Valid_4_delay_19_35;
  reg                 io_A_Valid_4_delay_20_34;
  reg                 io_A_Valid_4_delay_21_33;
  reg                 io_A_Valid_4_delay_22_32;
  reg                 io_A_Valid_4_delay_23_31;
  reg                 io_A_Valid_4_delay_24_30;
  reg                 io_A_Valid_4_delay_25_29;
  reg                 io_A_Valid_4_delay_26_28;
  reg                 io_A_Valid_4_delay_27_27;
  reg                 io_A_Valid_4_delay_28_26;
  reg                 io_A_Valid_4_delay_29_25;
  reg                 io_A_Valid_4_delay_30_24;
  reg                 io_A_Valid_4_delay_31_23;
  reg                 io_A_Valid_4_delay_32_22;
  reg                 io_A_Valid_4_delay_33_21;
  reg                 io_A_Valid_4_delay_34_20;
  reg                 io_A_Valid_4_delay_35_19;
  reg                 io_A_Valid_4_delay_36_18;
  reg                 io_A_Valid_4_delay_37_17;
  reg                 io_A_Valid_4_delay_38_16;
  reg                 io_A_Valid_4_delay_39_15;
  reg                 io_A_Valid_4_delay_40_14;
  reg                 io_A_Valid_4_delay_41_13;
  reg                 io_A_Valid_4_delay_42_12;
  reg                 io_A_Valid_4_delay_43_11;
  reg                 io_A_Valid_4_delay_44_10;
  reg                 io_A_Valid_4_delay_45_9;
  reg                 io_A_Valid_4_delay_46_8;
  reg                 io_A_Valid_4_delay_47_7;
  reg                 io_A_Valid_4_delay_48_6;
  reg                 io_A_Valid_4_delay_49_5;
  reg                 io_A_Valid_4_delay_50_4;
  reg                 io_A_Valid_4_delay_51_3;
  reg                 io_A_Valid_4_delay_52_2;
  reg                 io_A_Valid_4_delay_53_1;
  reg                 io_A_Valid_4_delay_54;
  reg                 io_B_Valid_54_delay_1_3;
  reg                 io_B_Valid_54_delay_2_2;
  reg                 io_B_Valid_54_delay_3_1;
  reg                 io_B_Valid_54_delay_4;
  reg                 io_A_Valid_4_delay_1_54;
  reg                 io_A_Valid_4_delay_2_53;
  reg                 io_A_Valid_4_delay_3_52;
  reg                 io_A_Valid_4_delay_4_51;
  reg                 io_A_Valid_4_delay_5_50;
  reg                 io_A_Valid_4_delay_6_49;
  reg                 io_A_Valid_4_delay_7_48;
  reg                 io_A_Valid_4_delay_8_47;
  reg                 io_A_Valid_4_delay_9_46;
  reg                 io_A_Valid_4_delay_10_45;
  reg                 io_A_Valid_4_delay_11_44;
  reg                 io_A_Valid_4_delay_12_43;
  reg                 io_A_Valid_4_delay_13_42;
  reg                 io_A_Valid_4_delay_14_41;
  reg                 io_A_Valid_4_delay_15_40;
  reg                 io_A_Valid_4_delay_16_39;
  reg                 io_A_Valid_4_delay_17_38;
  reg                 io_A_Valid_4_delay_18_37;
  reg                 io_A_Valid_4_delay_19_36;
  reg                 io_A_Valid_4_delay_20_35;
  reg                 io_A_Valid_4_delay_21_34;
  reg                 io_A_Valid_4_delay_22_33;
  reg                 io_A_Valid_4_delay_23_32;
  reg                 io_A_Valid_4_delay_24_31;
  reg                 io_A_Valid_4_delay_25_30;
  reg                 io_A_Valid_4_delay_26_29;
  reg                 io_A_Valid_4_delay_27_28;
  reg                 io_A_Valid_4_delay_28_27;
  reg                 io_A_Valid_4_delay_29_26;
  reg                 io_A_Valid_4_delay_30_25;
  reg                 io_A_Valid_4_delay_31_24;
  reg                 io_A_Valid_4_delay_32_23;
  reg                 io_A_Valid_4_delay_33_22;
  reg                 io_A_Valid_4_delay_34_21;
  reg                 io_A_Valid_4_delay_35_20;
  reg                 io_A_Valid_4_delay_36_19;
  reg                 io_A_Valid_4_delay_37_18;
  reg                 io_A_Valid_4_delay_38_17;
  reg                 io_A_Valid_4_delay_39_16;
  reg                 io_A_Valid_4_delay_40_15;
  reg                 io_A_Valid_4_delay_41_14;
  reg                 io_A_Valid_4_delay_42_13;
  reg                 io_A_Valid_4_delay_43_12;
  reg                 io_A_Valid_4_delay_44_11;
  reg                 io_A_Valid_4_delay_45_10;
  reg                 io_A_Valid_4_delay_46_9;
  reg                 io_A_Valid_4_delay_47_8;
  reg                 io_A_Valid_4_delay_48_7;
  reg                 io_A_Valid_4_delay_49_6;
  reg                 io_A_Valid_4_delay_50_5;
  reg                 io_A_Valid_4_delay_51_4;
  reg                 io_A_Valid_4_delay_52_3;
  reg                 io_A_Valid_4_delay_53_2;
  reg                 io_A_Valid_4_delay_54_1;
  reg                 io_A_Valid_4_delay_55;
  reg                 io_B_Valid_55_delay_1_3;
  reg                 io_B_Valid_55_delay_2_2;
  reg                 io_B_Valid_55_delay_3_1;
  reg                 io_B_Valid_55_delay_4;
  reg                 io_A_Valid_4_delay_1_55;
  reg                 io_A_Valid_4_delay_2_54;
  reg                 io_A_Valid_4_delay_3_53;
  reg                 io_A_Valid_4_delay_4_52;
  reg                 io_A_Valid_4_delay_5_51;
  reg                 io_A_Valid_4_delay_6_50;
  reg                 io_A_Valid_4_delay_7_49;
  reg                 io_A_Valid_4_delay_8_48;
  reg                 io_A_Valid_4_delay_9_47;
  reg                 io_A_Valid_4_delay_10_46;
  reg                 io_A_Valid_4_delay_11_45;
  reg                 io_A_Valid_4_delay_12_44;
  reg                 io_A_Valid_4_delay_13_43;
  reg                 io_A_Valid_4_delay_14_42;
  reg                 io_A_Valid_4_delay_15_41;
  reg                 io_A_Valid_4_delay_16_40;
  reg                 io_A_Valid_4_delay_17_39;
  reg                 io_A_Valid_4_delay_18_38;
  reg                 io_A_Valid_4_delay_19_37;
  reg                 io_A_Valid_4_delay_20_36;
  reg                 io_A_Valid_4_delay_21_35;
  reg                 io_A_Valid_4_delay_22_34;
  reg                 io_A_Valid_4_delay_23_33;
  reg                 io_A_Valid_4_delay_24_32;
  reg                 io_A_Valid_4_delay_25_31;
  reg                 io_A_Valid_4_delay_26_30;
  reg                 io_A_Valid_4_delay_27_29;
  reg                 io_A_Valid_4_delay_28_28;
  reg                 io_A_Valid_4_delay_29_27;
  reg                 io_A_Valid_4_delay_30_26;
  reg                 io_A_Valid_4_delay_31_25;
  reg                 io_A_Valid_4_delay_32_24;
  reg                 io_A_Valid_4_delay_33_23;
  reg                 io_A_Valid_4_delay_34_22;
  reg                 io_A_Valid_4_delay_35_21;
  reg                 io_A_Valid_4_delay_36_20;
  reg                 io_A_Valid_4_delay_37_19;
  reg                 io_A_Valid_4_delay_38_18;
  reg                 io_A_Valid_4_delay_39_17;
  reg                 io_A_Valid_4_delay_40_16;
  reg                 io_A_Valid_4_delay_41_15;
  reg                 io_A_Valid_4_delay_42_14;
  reg                 io_A_Valid_4_delay_43_13;
  reg                 io_A_Valid_4_delay_44_12;
  reg                 io_A_Valid_4_delay_45_11;
  reg                 io_A_Valid_4_delay_46_10;
  reg                 io_A_Valid_4_delay_47_9;
  reg                 io_A_Valid_4_delay_48_8;
  reg                 io_A_Valid_4_delay_49_7;
  reg                 io_A_Valid_4_delay_50_6;
  reg                 io_A_Valid_4_delay_51_5;
  reg                 io_A_Valid_4_delay_52_4;
  reg                 io_A_Valid_4_delay_53_3;
  reg                 io_A_Valid_4_delay_54_2;
  reg                 io_A_Valid_4_delay_55_1;
  reg                 io_A_Valid_4_delay_56;
  reg                 io_B_Valid_56_delay_1_3;
  reg                 io_B_Valid_56_delay_2_2;
  reg                 io_B_Valid_56_delay_3_1;
  reg                 io_B_Valid_56_delay_4;
  reg                 io_A_Valid_4_delay_1_56;
  reg                 io_A_Valid_4_delay_2_55;
  reg                 io_A_Valid_4_delay_3_54;
  reg                 io_A_Valid_4_delay_4_53;
  reg                 io_A_Valid_4_delay_5_52;
  reg                 io_A_Valid_4_delay_6_51;
  reg                 io_A_Valid_4_delay_7_50;
  reg                 io_A_Valid_4_delay_8_49;
  reg                 io_A_Valid_4_delay_9_48;
  reg                 io_A_Valid_4_delay_10_47;
  reg                 io_A_Valid_4_delay_11_46;
  reg                 io_A_Valid_4_delay_12_45;
  reg                 io_A_Valid_4_delay_13_44;
  reg                 io_A_Valid_4_delay_14_43;
  reg                 io_A_Valid_4_delay_15_42;
  reg                 io_A_Valid_4_delay_16_41;
  reg                 io_A_Valid_4_delay_17_40;
  reg                 io_A_Valid_4_delay_18_39;
  reg                 io_A_Valid_4_delay_19_38;
  reg                 io_A_Valid_4_delay_20_37;
  reg                 io_A_Valid_4_delay_21_36;
  reg                 io_A_Valid_4_delay_22_35;
  reg                 io_A_Valid_4_delay_23_34;
  reg                 io_A_Valid_4_delay_24_33;
  reg                 io_A_Valid_4_delay_25_32;
  reg                 io_A_Valid_4_delay_26_31;
  reg                 io_A_Valid_4_delay_27_30;
  reg                 io_A_Valid_4_delay_28_29;
  reg                 io_A_Valid_4_delay_29_28;
  reg                 io_A_Valid_4_delay_30_27;
  reg                 io_A_Valid_4_delay_31_26;
  reg                 io_A_Valid_4_delay_32_25;
  reg                 io_A_Valid_4_delay_33_24;
  reg                 io_A_Valid_4_delay_34_23;
  reg                 io_A_Valid_4_delay_35_22;
  reg                 io_A_Valid_4_delay_36_21;
  reg                 io_A_Valid_4_delay_37_20;
  reg                 io_A_Valid_4_delay_38_19;
  reg                 io_A_Valid_4_delay_39_18;
  reg                 io_A_Valid_4_delay_40_17;
  reg                 io_A_Valid_4_delay_41_16;
  reg                 io_A_Valid_4_delay_42_15;
  reg                 io_A_Valid_4_delay_43_14;
  reg                 io_A_Valid_4_delay_44_13;
  reg                 io_A_Valid_4_delay_45_12;
  reg                 io_A_Valid_4_delay_46_11;
  reg                 io_A_Valid_4_delay_47_10;
  reg                 io_A_Valid_4_delay_48_9;
  reg                 io_A_Valid_4_delay_49_8;
  reg                 io_A_Valid_4_delay_50_7;
  reg                 io_A_Valid_4_delay_51_6;
  reg                 io_A_Valid_4_delay_52_5;
  reg                 io_A_Valid_4_delay_53_4;
  reg                 io_A_Valid_4_delay_54_3;
  reg                 io_A_Valid_4_delay_55_2;
  reg                 io_A_Valid_4_delay_56_1;
  reg                 io_A_Valid_4_delay_57;
  reg                 io_B_Valid_57_delay_1_3;
  reg                 io_B_Valid_57_delay_2_2;
  reg                 io_B_Valid_57_delay_3_1;
  reg                 io_B_Valid_57_delay_4;
  reg                 io_A_Valid_4_delay_1_57;
  reg                 io_A_Valid_4_delay_2_56;
  reg                 io_A_Valid_4_delay_3_55;
  reg                 io_A_Valid_4_delay_4_54;
  reg                 io_A_Valid_4_delay_5_53;
  reg                 io_A_Valid_4_delay_6_52;
  reg                 io_A_Valid_4_delay_7_51;
  reg                 io_A_Valid_4_delay_8_50;
  reg                 io_A_Valid_4_delay_9_49;
  reg                 io_A_Valid_4_delay_10_48;
  reg                 io_A_Valid_4_delay_11_47;
  reg                 io_A_Valid_4_delay_12_46;
  reg                 io_A_Valid_4_delay_13_45;
  reg                 io_A_Valid_4_delay_14_44;
  reg                 io_A_Valid_4_delay_15_43;
  reg                 io_A_Valid_4_delay_16_42;
  reg                 io_A_Valid_4_delay_17_41;
  reg                 io_A_Valid_4_delay_18_40;
  reg                 io_A_Valid_4_delay_19_39;
  reg                 io_A_Valid_4_delay_20_38;
  reg                 io_A_Valid_4_delay_21_37;
  reg                 io_A_Valid_4_delay_22_36;
  reg                 io_A_Valid_4_delay_23_35;
  reg                 io_A_Valid_4_delay_24_34;
  reg                 io_A_Valid_4_delay_25_33;
  reg                 io_A_Valid_4_delay_26_32;
  reg                 io_A_Valid_4_delay_27_31;
  reg                 io_A_Valid_4_delay_28_30;
  reg                 io_A_Valid_4_delay_29_29;
  reg                 io_A_Valid_4_delay_30_28;
  reg                 io_A_Valid_4_delay_31_27;
  reg                 io_A_Valid_4_delay_32_26;
  reg                 io_A_Valid_4_delay_33_25;
  reg                 io_A_Valid_4_delay_34_24;
  reg                 io_A_Valid_4_delay_35_23;
  reg                 io_A_Valid_4_delay_36_22;
  reg                 io_A_Valid_4_delay_37_21;
  reg                 io_A_Valid_4_delay_38_20;
  reg                 io_A_Valid_4_delay_39_19;
  reg                 io_A_Valid_4_delay_40_18;
  reg                 io_A_Valid_4_delay_41_17;
  reg                 io_A_Valid_4_delay_42_16;
  reg                 io_A_Valid_4_delay_43_15;
  reg                 io_A_Valid_4_delay_44_14;
  reg                 io_A_Valid_4_delay_45_13;
  reg                 io_A_Valid_4_delay_46_12;
  reg                 io_A_Valid_4_delay_47_11;
  reg                 io_A_Valid_4_delay_48_10;
  reg                 io_A_Valid_4_delay_49_9;
  reg                 io_A_Valid_4_delay_50_8;
  reg                 io_A_Valid_4_delay_51_7;
  reg                 io_A_Valid_4_delay_52_6;
  reg                 io_A_Valid_4_delay_53_5;
  reg                 io_A_Valid_4_delay_54_4;
  reg                 io_A_Valid_4_delay_55_3;
  reg                 io_A_Valid_4_delay_56_2;
  reg                 io_A_Valid_4_delay_57_1;
  reg                 io_A_Valid_4_delay_58;
  reg                 io_B_Valid_58_delay_1_3;
  reg                 io_B_Valid_58_delay_2_2;
  reg                 io_B_Valid_58_delay_3_1;
  reg                 io_B_Valid_58_delay_4;
  reg                 io_A_Valid_4_delay_1_58;
  reg                 io_A_Valid_4_delay_2_57;
  reg                 io_A_Valid_4_delay_3_56;
  reg                 io_A_Valid_4_delay_4_55;
  reg                 io_A_Valid_4_delay_5_54;
  reg                 io_A_Valid_4_delay_6_53;
  reg                 io_A_Valid_4_delay_7_52;
  reg                 io_A_Valid_4_delay_8_51;
  reg                 io_A_Valid_4_delay_9_50;
  reg                 io_A_Valid_4_delay_10_49;
  reg                 io_A_Valid_4_delay_11_48;
  reg                 io_A_Valid_4_delay_12_47;
  reg                 io_A_Valid_4_delay_13_46;
  reg                 io_A_Valid_4_delay_14_45;
  reg                 io_A_Valid_4_delay_15_44;
  reg                 io_A_Valid_4_delay_16_43;
  reg                 io_A_Valid_4_delay_17_42;
  reg                 io_A_Valid_4_delay_18_41;
  reg                 io_A_Valid_4_delay_19_40;
  reg                 io_A_Valid_4_delay_20_39;
  reg                 io_A_Valid_4_delay_21_38;
  reg                 io_A_Valid_4_delay_22_37;
  reg                 io_A_Valid_4_delay_23_36;
  reg                 io_A_Valid_4_delay_24_35;
  reg                 io_A_Valid_4_delay_25_34;
  reg                 io_A_Valid_4_delay_26_33;
  reg                 io_A_Valid_4_delay_27_32;
  reg                 io_A_Valid_4_delay_28_31;
  reg                 io_A_Valid_4_delay_29_30;
  reg                 io_A_Valid_4_delay_30_29;
  reg                 io_A_Valid_4_delay_31_28;
  reg                 io_A_Valid_4_delay_32_27;
  reg                 io_A_Valid_4_delay_33_26;
  reg                 io_A_Valid_4_delay_34_25;
  reg                 io_A_Valid_4_delay_35_24;
  reg                 io_A_Valid_4_delay_36_23;
  reg                 io_A_Valid_4_delay_37_22;
  reg                 io_A_Valid_4_delay_38_21;
  reg                 io_A_Valid_4_delay_39_20;
  reg                 io_A_Valid_4_delay_40_19;
  reg                 io_A_Valid_4_delay_41_18;
  reg                 io_A_Valid_4_delay_42_17;
  reg                 io_A_Valid_4_delay_43_16;
  reg                 io_A_Valid_4_delay_44_15;
  reg                 io_A_Valid_4_delay_45_14;
  reg                 io_A_Valid_4_delay_46_13;
  reg                 io_A_Valid_4_delay_47_12;
  reg                 io_A_Valid_4_delay_48_11;
  reg                 io_A_Valid_4_delay_49_10;
  reg                 io_A_Valid_4_delay_50_9;
  reg                 io_A_Valid_4_delay_51_8;
  reg                 io_A_Valid_4_delay_52_7;
  reg                 io_A_Valid_4_delay_53_6;
  reg                 io_A_Valid_4_delay_54_5;
  reg                 io_A_Valid_4_delay_55_4;
  reg                 io_A_Valid_4_delay_56_3;
  reg                 io_A_Valid_4_delay_57_2;
  reg                 io_A_Valid_4_delay_58_1;
  reg                 io_A_Valid_4_delay_59;
  reg                 io_B_Valid_59_delay_1_3;
  reg                 io_B_Valid_59_delay_2_2;
  reg                 io_B_Valid_59_delay_3_1;
  reg                 io_B_Valid_59_delay_4;
  reg                 io_A_Valid_4_delay_1_59;
  reg                 io_A_Valid_4_delay_2_58;
  reg                 io_A_Valid_4_delay_3_57;
  reg                 io_A_Valid_4_delay_4_56;
  reg                 io_A_Valid_4_delay_5_55;
  reg                 io_A_Valid_4_delay_6_54;
  reg                 io_A_Valid_4_delay_7_53;
  reg                 io_A_Valid_4_delay_8_52;
  reg                 io_A_Valid_4_delay_9_51;
  reg                 io_A_Valid_4_delay_10_50;
  reg                 io_A_Valid_4_delay_11_49;
  reg                 io_A_Valid_4_delay_12_48;
  reg                 io_A_Valid_4_delay_13_47;
  reg                 io_A_Valid_4_delay_14_46;
  reg                 io_A_Valid_4_delay_15_45;
  reg                 io_A_Valid_4_delay_16_44;
  reg                 io_A_Valid_4_delay_17_43;
  reg                 io_A_Valid_4_delay_18_42;
  reg                 io_A_Valid_4_delay_19_41;
  reg                 io_A_Valid_4_delay_20_40;
  reg                 io_A_Valid_4_delay_21_39;
  reg                 io_A_Valid_4_delay_22_38;
  reg                 io_A_Valid_4_delay_23_37;
  reg                 io_A_Valid_4_delay_24_36;
  reg                 io_A_Valid_4_delay_25_35;
  reg                 io_A_Valid_4_delay_26_34;
  reg                 io_A_Valid_4_delay_27_33;
  reg                 io_A_Valid_4_delay_28_32;
  reg                 io_A_Valid_4_delay_29_31;
  reg                 io_A_Valid_4_delay_30_30;
  reg                 io_A_Valid_4_delay_31_29;
  reg                 io_A_Valid_4_delay_32_28;
  reg                 io_A_Valid_4_delay_33_27;
  reg                 io_A_Valid_4_delay_34_26;
  reg                 io_A_Valid_4_delay_35_25;
  reg                 io_A_Valid_4_delay_36_24;
  reg                 io_A_Valid_4_delay_37_23;
  reg                 io_A_Valid_4_delay_38_22;
  reg                 io_A_Valid_4_delay_39_21;
  reg                 io_A_Valid_4_delay_40_20;
  reg                 io_A_Valid_4_delay_41_19;
  reg                 io_A_Valid_4_delay_42_18;
  reg                 io_A_Valid_4_delay_43_17;
  reg                 io_A_Valid_4_delay_44_16;
  reg                 io_A_Valid_4_delay_45_15;
  reg                 io_A_Valid_4_delay_46_14;
  reg                 io_A_Valid_4_delay_47_13;
  reg                 io_A_Valid_4_delay_48_12;
  reg                 io_A_Valid_4_delay_49_11;
  reg                 io_A_Valid_4_delay_50_10;
  reg                 io_A_Valid_4_delay_51_9;
  reg                 io_A_Valid_4_delay_52_8;
  reg                 io_A_Valid_4_delay_53_7;
  reg                 io_A_Valid_4_delay_54_6;
  reg                 io_A_Valid_4_delay_55_5;
  reg                 io_A_Valid_4_delay_56_4;
  reg                 io_A_Valid_4_delay_57_3;
  reg                 io_A_Valid_4_delay_58_2;
  reg                 io_A_Valid_4_delay_59_1;
  reg                 io_A_Valid_4_delay_60;
  reg                 io_B_Valid_60_delay_1_3;
  reg                 io_B_Valid_60_delay_2_2;
  reg                 io_B_Valid_60_delay_3_1;
  reg                 io_B_Valid_60_delay_4;
  reg                 io_A_Valid_4_delay_1_60;
  reg                 io_A_Valid_4_delay_2_59;
  reg                 io_A_Valid_4_delay_3_58;
  reg                 io_A_Valid_4_delay_4_57;
  reg                 io_A_Valid_4_delay_5_56;
  reg                 io_A_Valid_4_delay_6_55;
  reg                 io_A_Valid_4_delay_7_54;
  reg                 io_A_Valid_4_delay_8_53;
  reg                 io_A_Valid_4_delay_9_52;
  reg                 io_A_Valid_4_delay_10_51;
  reg                 io_A_Valid_4_delay_11_50;
  reg                 io_A_Valid_4_delay_12_49;
  reg                 io_A_Valid_4_delay_13_48;
  reg                 io_A_Valid_4_delay_14_47;
  reg                 io_A_Valid_4_delay_15_46;
  reg                 io_A_Valid_4_delay_16_45;
  reg                 io_A_Valid_4_delay_17_44;
  reg                 io_A_Valid_4_delay_18_43;
  reg                 io_A_Valid_4_delay_19_42;
  reg                 io_A_Valid_4_delay_20_41;
  reg                 io_A_Valid_4_delay_21_40;
  reg                 io_A_Valid_4_delay_22_39;
  reg                 io_A_Valid_4_delay_23_38;
  reg                 io_A_Valid_4_delay_24_37;
  reg                 io_A_Valid_4_delay_25_36;
  reg                 io_A_Valid_4_delay_26_35;
  reg                 io_A_Valid_4_delay_27_34;
  reg                 io_A_Valid_4_delay_28_33;
  reg                 io_A_Valid_4_delay_29_32;
  reg                 io_A_Valid_4_delay_30_31;
  reg                 io_A_Valid_4_delay_31_30;
  reg                 io_A_Valid_4_delay_32_29;
  reg                 io_A_Valid_4_delay_33_28;
  reg                 io_A_Valid_4_delay_34_27;
  reg                 io_A_Valid_4_delay_35_26;
  reg                 io_A_Valid_4_delay_36_25;
  reg                 io_A_Valid_4_delay_37_24;
  reg                 io_A_Valid_4_delay_38_23;
  reg                 io_A_Valid_4_delay_39_22;
  reg                 io_A_Valid_4_delay_40_21;
  reg                 io_A_Valid_4_delay_41_20;
  reg                 io_A_Valid_4_delay_42_19;
  reg                 io_A_Valid_4_delay_43_18;
  reg                 io_A_Valid_4_delay_44_17;
  reg                 io_A_Valid_4_delay_45_16;
  reg                 io_A_Valid_4_delay_46_15;
  reg                 io_A_Valid_4_delay_47_14;
  reg                 io_A_Valid_4_delay_48_13;
  reg                 io_A_Valid_4_delay_49_12;
  reg                 io_A_Valid_4_delay_50_11;
  reg                 io_A_Valid_4_delay_51_10;
  reg                 io_A_Valid_4_delay_52_9;
  reg                 io_A_Valid_4_delay_53_8;
  reg                 io_A_Valid_4_delay_54_7;
  reg                 io_A_Valid_4_delay_55_6;
  reg                 io_A_Valid_4_delay_56_5;
  reg                 io_A_Valid_4_delay_57_4;
  reg                 io_A_Valid_4_delay_58_3;
  reg                 io_A_Valid_4_delay_59_2;
  reg                 io_A_Valid_4_delay_60_1;
  reg                 io_A_Valid_4_delay_61;
  reg                 io_B_Valid_61_delay_1_3;
  reg                 io_B_Valid_61_delay_2_2;
  reg                 io_B_Valid_61_delay_3_1;
  reg                 io_B_Valid_61_delay_4;
  reg                 io_A_Valid_4_delay_1_61;
  reg                 io_A_Valid_4_delay_2_60;
  reg                 io_A_Valid_4_delay_3_59;
  reg                 io_A_Valid_4_delay_4_58;
  reg                 io_A_Valid_4_delay_5_57;
  reg                 io_A_Valid_4_delay_6_56;
  reg                 io_A_Valid_4_delay_7_55;
  reg                 io_A_Valid_4_delay_8_54;
  reg                 io_A_Valid_4_delay_9_53;
  reg                 io_A_Valid_4_delay_10_52;
  reg                 io_A_Valid_4_delay_11_51;
  reg                 io_A_Valid_4_delay_12_50;
  reg                 io_A_Valid_4_delay_13_49;
  reg                 io_A_Valid_4_delay_14_48;
  reg                 io_A_Valid_4_delay_15_47;
  reg                 io_A_Valid_4_delay_16_46;
  reg                 io_A_Valid_4_delay_17_45;
  reg                 io_A_Valid_4_delay_18_44;
  reg                 io_A_Valid_4_delay_19_43;
  reg                 io_A_Valid_4_delay_20_42;
  reg                 io_A_Valid_4_delay_21_41;
  reg                 io_A_Valid_4_delay_22_40;
  reg                 io_A_Valid_4_delay_23_39;
  reg                 io_A_Valid_4_delay_24_38;
  reg                 io_A_Valid_4_delay_25_37;
  reg                 io_A_Valid_4_delay_26_36;
  reg                 io_A_Valid_4_delay_27_35;
  reg                 io_A_Valid_4_delay_28_34;
  reg                 io_A_Valid_4_delay_29_33;
  reg                 io_A_Valid_4_delay_30_32;
  reg                 io_A_Valid_4_delay_31_31;
  reg                 io_A_Valid_4_delay_32_30;
  reg                 io_A_Valid_4_delay_33_29;
  reg                 io_A_Valid_4_delay_34_28;
  reg                 io_A_Valid_4_delay_35_27;
  reg                 io_A_Valid_4_delay_36_26;
  reg                 io_A_Valid_4_delay_37_25;
  reg                 io_A_Valid_4_delay_38_24;
  reg                 io_A_Valid_4_delay_39_23;
  reg                 io_A_Valid_4_delay_40_22;
  reg                 io_A_Valid_4_delay_41_21;
  reg                 io_A_Valid_4_delay_42_20;
  reg                 io_A_Valid_4_delay_43_19;
  reg                 io_A_Valid_4_delay_44_18;
  reg                 io_A_Valid_4_delay_45_17;
  reg                 io_A_Valid_4_delay_46_16;
  reg                 io_A_Valid_4_delay_47_15;
  reg                 io_A_Valid_4_delay_48_14;
  reg                 io_A_Valid_4_delay_49_13;
  reg                 io_A_Valid_4_delay_50_12;
  reg                 io_A_Valid_4_delay_51_11;
  reg                 io_A_Valid_4_delay_52_10;
  reg                 io_A_Valid_4_delay_53_9;
  reg                 io_A_Valid_4_delay_54_8;
  reg                 io_A_Valid_4_delay_55_7;
  reg                 io_A_Valid_4_delay_56_6;
  reg                 io_A_Valid_4_delay_57_5;
  reg                 io_A_Valid_4_delay_58_4;
  reg                 io_A_Valid_4_delay_59_3;
  reg                 io_A_Valid_4_delay_60_2;
  reg                 io_A_Valid_4_delay_61_1;
  reg                 io_A_Valid_4_delay_62;
  reg                 io_B_Valid_62_delay_1_3;
  reg                 io_B_Valid_62_delay_2_2;
  reg                 io_B_Valid_62_delay_3_1;
  reg                 io_B_Valid_62_delay_4;
  reg                 io_A_Valid_4_delay_1_62;
  reg                 io_A_Valid_4_delay_2_61;
  reg                 io_A_Valid_4_delay_3_60;
  reg                 io_A_Valid_4_delay_4_59;
  reg                 io_A_Valid_4_delay_5_58;
  reg                 io_A_Valid_4_delay_6_57;
  reg                 io_A_Valid_4_delay_7_56;
  reg                 io_A_Valid_4_delay_8_55;
  reg                 io_A_Valid_4_delay_9_54;
  reg                 io_A_Valid_4_delay_10_53;
  reg                 io_A_Valid_4_delay_11_52;
  reg                 io_A_Valid_4_delay_12_51;
  reg                 io_A_Valid_4_delay_13_50;
  reg                 io_A_Valid_4_delay_14_49;
  reg                 io_A_Valid_4_delay_15_48;
  reg                 io_A_Valid_4_delay_16_47;
  reg                 io_A_Valid_4_delay_17_46;
  reg                 io_A_Valid_4_delay_18_45;
  reg                 io_A_Valid_4_delay_19_44;
  reg                 io_A_Valid_4_delay_20_43;
  reg                 io_A_Valid_4_delay_21_42;
  reg                 io_A_Valid_4_delay_22_41;
  reg                 io_A_Valid_4_delay_23_40;
  reg                 io_A_Valid_4_delay_24_39;
  reg                 io_A_Valid_4_delay_25_38;
  reg                 io_A_Valid_4_delay_26_37;
  reg                 io_A_Valid_4_delay_27_36;
  reg                 io_A_Valid_4_delay_28_35;
  reg                 io_A_Valid_4_delay_29_34;
  reg                 io_A_Valid_4_delay_30_33;
  reg                 io_A_Valid_4_delay_31_32;
  reg                 io_A_Valid_4_delay_32_31;
  reg                 io_A_Valid_4_delay_33_30;
  reg                 io_A_Valid_4_delay_34_29;
  reg                 io_A_Valid_4_delay_35_28;
  reg                 io_A_Valid_4_delay_36_27;
  reg                 io_A_Valid_4_delay_37_26;
  reg                 io_A_Valid_4_delay_38_25;
  reg                 io_A_Valid_4_delay_39_24;
  reg                 io_A_Valid_4_delay_40_23;
  reg                 io_A_Valid_4_delay_41_22;
  reg                 io_A_Valid_4_delay_42_21;
  reg                 io_A_Valid_4_delay_43_20;
  reg                 io_A_Valid_4_delay_44_19;
  reg                 io_A_Valid_4_delay_45_18;
  reg                 io_A_Valid_4_delay_46_17;
  reg                 io_A_Valid_4_delay_47_16;
  reg                 io_A_Valid_4_delay_48_15;
  reg                 io_A_Valid_4_delay_49_14;
  reg                 io_A_Valid_4_delay_50_13;
  reg                 io_A_Valid_4_delay_51_12;
  reg                 io_A_Valid_4_delay_52_11;
  reg                 io_A_Valid_4_delay_53_10;
  reg                 io_A_Valid_4_delay_54_9;
  reg                 io_A_Valid_4_delay_55_8;
  reg                 io_A_Valid_4_delay_56_7;
  reg                 io_A_Valid_4_delay_57_6;
  reg                 io_A_Valid_4_delay_58_5;
  reg                 io_A_Valid_4_delay_59_4;
  reg                 io_A_Valid_4_delay_60_3;
  reg                 io_A_Valid_4_delay_61_2;
  reg                 io_A_Valid_4_delay_62_1;
  reg                 io_A_Valid_4_delay_63;
  reg                 io_B_Valid_63_delay_1_3;
  reg                 io_B_Valid_63_delay_2_2;
  reg                 io_B_Valid_63_delay_3_1;
  reg                 io_B_Valid_63_delay_4;
  reg        [15:0]   io_signCount_regNextWhen_5;
  reg                 io_B_Valid_0_delay_1_4;
  reg                 io_B_Valid_0_delay_2_3;
  reg                 io_B_Valid_0_delay_3_2;
  reg                 io_B_Valid_0_delay_4_1;
  reg                 io_B_Valid_0_delay_5;
  reg                 io_A_Valid_5_delay_1;
  reg                 io_B_Valid_1_delay_1_4;
  reg                 io_B_Valid_1_delay_2_3;
  reg                 io_B_Valid_1_delay_3_2;
  reg                 io_B_Valid_1_delay_4_1;
  reg                 io_B_Valid_1_delay_5;
  reg                 io_A_Valid_5_delay_1_1;
  reg                 io_A_Valid_5_delay_2;
  reg                 io_B_Valid_2_delay_1_4;
  reg                 io_B_Valid_2_delay_2_3;
  reg                 io_B_Valid_2_delay_3_2;
  reg                 io_B_Valid_2_delay_4_1;
  reg                 io_B_Valid_2_delay_5;
  reg                 io_A_Valid_5_delay_1_2;
  reg                 io_A_Valid_5_delay_2_1;
  reg                 io_A_Valid_5_delay_3;
  reg                 io_B_Valid_3_delay_1_4;
  reg                 io_B_Valid_3_delay_2_3;
  reg                 io_B_Valid_3_delay_3_2;
  reg                 io_B_Valid_3_delay_4_1;
  reg                 io_B_Valid_3_delay_5;
  reg                 io_A_Valid_5_delay_1_3;
  reg                 io_A_Valid_5_delay_2_2;
  reg                 io_A_Valid_5_delay_3_1;
  reg                 io_A_Valid_5_delay_4;
  reg                 io_B_Valid_4_delay_1_4;
  reg                 io_B_Valid_4_delay_2_3;
  reg                 io_B_Valid_4_delay_3_2;
  reg                 io_B_Valid_4_delay_4_1;
  reg                 io_B_Valid_4_delay_5;
  reg                 io_A_Valid_5_delay_1_4;
  reg                 io_A_Valid_5_delay_2_3;
  reg                 io_A_Valid_5_delay_3_2;
  reg                 io_A_Valid_5_delay_4_1;
  reg                 io_A_Valid_5_delay_5;
  reg                 io_B_Valid_5_delay_1_4;
  reg                 io_B_Valid_5_delay_2_3;
  reg                 io_B_Valid_5_delay_3_2;
  reg                 io_B_Valid_5_delay_4_1;
  reg                 io_B_Valid_5_delay_5;
  reg                 io_A_Valid_5_delay_1_5;
  reg                 io_A_Valid_5_delay_2_4;
  reg                 io_A_Valid_5_delay_3_3;
  reg                 io_A_Valid_5_delay_4_2;
  reg                 io_A_Valid_5_delay_5_1;
  reg                 io_A_Valid_5_delay_6;
  reg                 io_B_Valid_6_delay_1_4;
  reg                 io_B_Valid_6_delay_2_3;
  reg                 io_B_Valid_6_delay_3_2;
  reg                 io_B_Valid_6_delay_4_1;
  reg                 io_B_Valid_6_delay_5;
  reg                 io_A_Valid_5_delay_1_6;
  reg                 io_A_Valid_5_delay_2_5;
  reg                 io_A_Valid_5_delay_3_4;
  reg                 io_A_Valid_5_delay_4_3;
  reg                 io_A_Valid_5_delay_5_2;
  reg                 io_A_Valid_5_delay_6_1;
  reg                 io_A_Valid_5_delay_7;
  reg                 io_B_Valid_7_delay_1_4;
  reg                 io_B_Valid_7_delay_2_3;
  reg                 io_B_Valid_7_delay_3_2;
  reg                 io_B_Valid_7_delay_4_1;
  reg                 io_B_Valid_7_delay_5;
  reg                 io_A_Valid_5_delay_1_7;
  reg                 io_A_Valid_5_delay_2_6;
  reg                 io_A_Valid_5_delay_3_5;
  reg                 io_A_Valid_5_delay_4_4;
  reg                 io_A_Valid_5_delay_5_3;
  reg                 io_A_Valid_5_delay_6_2;
  reg                 io_A_Valid_5_delay_7_1;
  reg                 io_A_Valid_5_delay_8;
  reg                 io_B_Valid_8_delay_1_4;
  reg                 io_B_Valid_8_delay_2_3;
  reg                 io_B_Valid_8_delay_3_2;
  reg                 io_B_Valid_8_delay_4_1;
  reg                 io_B_Valid_8_delay_5;
  reg                 io_A_Valid_5_delay_1_8;
  reg                 io_A_Valid_5_delay_2_7;
  reg                 io_A_Valid_5_delay_3_6;
  reg                 io_A_Valid_5_delay_4_5;
  reg                 io_A_Valid_5_delay_5_4;
  reg                 io_A_Valid_5_delay_6_3;
  reg                 io_A_Valid_5_delay_7_2;
  reg                 io_A_Valid_5_delay_8_1;
  reg                 io_A_Valid_5_delay_9;
  reg                 io_B_Valid_9_delay_1_4;
  reg                 io_B_Valid_9_delay_2_3;
  reg                 io_B_Valid_9_delay_3_2;
  reg                 io_B_Valid_9_delay_4_1;
  reg                 io_B_Valid_9_delay_5;
  reg                 io_A_Valid_5_delay_1_9;
  reg                 io_A_Valid_5_delay_2_8;
  reg                 io_A_Valid_5_delay_3_7;
  reg                 io_A_Valid_5_delay_4_6;
  reg                 io_A_Valid_5_delay_5_5;
  reg                 io_A_Valid_5_delay_6_4;
  reg                 io_A_Valid_5_delay_7_3;
  reg                 io_A_Valid_5_delay_8_2;
  reg                 io_A_Valid_5_delay_9_1;
  reg                 io_A_Valid_5_delay_10;
  reg                 io_B_Valid_10_delay_1_4;
  reg                 io_B_Valid_10_delay_2_3;
  reg                 io_B_Valid_10_delay_3_2;
  reg                 io_B_Valid_10_delay_4_1;
  reg                 io_B_Valid_10_delay_5;
  reg                 io_A_Valid_5_delay_1_10;
  reg                 io_A_Valid_5_delay_2_9;
  reg                 io_A_Valid_5_delay_3_8;
  reg                 io_A_Valid_5_delay_4_7;
  reg                 io_A_Valid_5_delay_5_6;
  reg                 io_A_Valid_5_delay_6_5;
  reg                 io_A_Valid_5_delay_7_4;
  reg                 io_A_Valid_5_delay_8_3;
  reg                 io_A_Valid_5_delay_9_2;
  reg                 io_A_Valid_5_delay_10_1;
  reg                 io_A_Valid_5_delay_11;
  reg                 io_B_Valid_11_delay_1_4;
  reg                 io_B_Valid_11_delay_2_3;
  reg                 io_B_Valid_11_delay_3_2;
  reg                 io_B_Valid_11_delay_4_1;
  reg                 io_B_Valid_11_delay_5;
  reg                 io_A_Valid_5_delay_1_11;
  reg                 io_A_Valid_5_delay_2_10;
  reg                 io_A_Valid_5_delay_3_9;
  reg                 io_A_Valid_5_delay_4_8;
  reg                 io_A_Valid_5_delay_5_7;
  reg                 io_A_Valid_5_delay_6_6;
  reg                 io_A_Valid_5_delay_7_5;
  reg                 io_A_Valid_5_delay_8_4;
  reg                 io_A_Valid_5_delay_9_3;
  reg                 io_A_Valid_5_delay_10_2;
  reg                 io_A_Valid_5_delay_11_1;
  reg                 io_A_Valid_5_delay_12;
  reg                 io_B_Valid_12_delay_1_4;
  reg                 io_B_Valid_12_delay_2_3;
  reg                 io_B_Valid_12_delay_3_2;
  reg                 io_B_Valid_12_delay_4_1;
  reg                 io_B_Valid_12_delay_5;
  reg                 io_A_Valid_5_delay_1_12;
  reg                 io_A_Valid_5_delay_2_11;
  reg                 io_A_Valid_5_delay_3_10;
  reg                 io_A_Valid_5_delay_4_9;
  reg                 io_A_Valid_5_delay_5_8;
  reg                 io_A_Valid_5_delay_6_7;
  reg                 io_A_Valid_5_delay_7_6;
  reg                 io_A_Valid_5_delay_8_5;
  reg                 io_A_Valid_5_delay_9_4;
  reg                 io_A_Valid_5_delay_10_3;
  reg                 io_A_Valid_5_delay_11_2;
  reg                 io_A_Valid_5_delay_12_1;
  reg                 io_A_Valid_5_delay_13;
  reg                 io_B_Valid_13_delay_1_4;
  reg                 io_B_Valid_13_delay_2_3;
  reg                 io_B_Valid_13_delay_3_2;
  reg                 io_B_Valid_13_delay_4_1;
  reg                 io_B_Valid_13_delay_5;
  reg                 io_A_Valid_5_delay_1_13;
  reg                 io_A_Valid_5_delay_2_12;
  reg                 io_A_Valid_5_delay_3_11;
  reg                 io_A_Valid_5_delay_4_10;
  reg                 io_A_Valid_5_delay_5_9;
  reg                 io_A_Valid_5_delay_6_8;
  reg                 io_A_Valid_5_delay_7_7;
  reg                 io_A_Valid_5_delay_8_6;
  reg                 io_A_Valid_5_delay_9_5;
  reg                 io_A_Valid_5_delay_10_4;
  reg                 io_A_Valid_5_delay_11_3;
  reg                 io_A_Valid_5_delay_12_2;
  reg                 io_A_Valid_5_delay_13_1;
  reg                 io_A_Valid_5_delay_14;
  reg                 io_B_Valid_14_delay_1_4;
  reg                 io_B_Valid_14_delay_2_3;
  reg                 io_B_Valid_14_delay_3_2;
  reg                 io_B_Valid_14_delay_4_1;
  reg                 io_B_Valid_14_delay_5;
  reg                 io_A_Valid_5_delay_1_14;
  reg                 io_A_Valid_5_delay_2_13;
  reg                 io_A_Valid_5_delay_3_12;
  reg                 io_A_Valid_5_delay_4_11;
  reg                 io_A_Valid_5_delay_5_10;
  reg                 io_A_Valid_5_delay_6_9;
  reg                 io_A_Valid_5_delay_7_8;
  reg                 io_A_Valid_5_delay_8_7;
  reg                 io_A_Valid_5_delay_9_6;
  reg                 io_A_Valid_5_delay_10_5;
  reg                 io_A_Valid_5_delay_11_4;
  reg                 io_A_Valid_5_delay_12_3;
  reg                 io_A_Valid_5_delay_13_2;
  reg                 io_A_Valid_5_delay_14_1;
  reg                 io_A_Valid_5_delay_15;
  reg                 io_B_Valid_15_delay_1_4;
  reg                 io_B_Valid_15_delay_2_3;
  reg                 io_B_Valid_15_delay_3_2;
  reg                 io_B_Valid_15_delay_4_1;
  reg                 io_B_Valid_15_delay_5;
  reg                 io_A_Valid_5_delay_1_15;
  reg                 io_A_Valid_5_delay_2_14;
  reg                 io_A_Valid_5_delay_3_13;
  reg                 io_A_Valid_5_delay_4_12;
  reg                 io_A_Valid_5_delay_5_11;
  reg                 io_A_Valid_5_delay_6_10;
  reg                 io_A_Valid_5_delay_7_9;
  reg                 io_A_Valid_5_delay_8_8;
  reg                 io_A_Valid_5_delay_9_7;
  reg                 io_A_Valid_5_delay_10_6;
  reg                 io_A_Valid_5_delay_11_5;
  reg                 io_A_Valid_5_delay_12_4;
  reg                 io_A_Valid_5_delay_13_3;
  reg                 io_A_Valid_5_delay_14_2;
  reg                 io_A_Valid_5_delay_15_1;
  reg                 io_A_Valid_5_delay_16;
  reg                 io_B_Valid_16_delay_1_4;
  reg                 io_B_Valid_16_delay_2_3;
  reg                 io_B_Valid_16_delay_3_2;
  reg                 io_B_Valid_16_delay_4_1;
  reg                 io_B_Valid_16_delay_5;
  reg                 io_A_Valid_5_delay_1_16;
  reg                 io_A_Valid_5_delay_2_15;
  reg                 io_A_Valid_5_delay_3_14;
  reg                 io_A_Valid_5_delay_4_13;
  reg                 io_A_Valid_5_delay_5_12;
  reg                 io_A_Valid_5_delay_6_11;
  reg                 io_A_Valid_5_delay_7_10;
  reg                 io_A_Valid_5_delay_8_9;
  reg                 io_A_Valid_5_delay_9_8;
  reg                 io_A_Valid_5_delay_10_7;
  reg                 io_A_Valid_5_delay_11_6;
  reg                 io_A_Valid_5_delay_12_5;
  reg                 io_A_Valid_5_delay_13_4;
  reg                 io_A_Valid_5_delay_14_3;
  reg                 io_A_Valid_5_delay_15_2;
  reg                 io_A_Valid_5_delay_16_1;
  reg                 io_A_Valid_5_delay_17;
  reg                 io_B_Valid_17_delay_1_4;
  reg                 io_B_Valid_17_delay_2_3;
  reg                 io_B_Valid_17_delay_3_2;
  reg                 io_B_Valid_17_delay_4_1;
  reg                 io_B_Valid_17_delay_5;
  reg                 io_A_Valid_5_delay_1_17;
  reg                 io_A_Valid_5_delay_2_16;
  reg                 io_A_Valid_5_delay_3_15;
  reg                 io_A_Valid_5_delay_4_14;
  reg                 io_A_Valid_5_delay_5_13;
  reg                 io_A_Valid_5_delay_6_12;
  reg                 io_A_Valid_5_delay_7_11;
  reg                 io_A_Valid_5_delay_8_10;
  reg                 io_A_Valid_5_delay_9_9;
  reg                 io_A_Valid_5_delay_10_8;
  reg                 io_A_Valid_5_delay_11_7;
  reg                 io_A_Valid_5_delay_12_6;
  reg                 io_A_Valid_5_delay_13_5;
  reg                 io_A_Valid_5_delay_14_4;
  reg                 io_A_Valid_5_delay_15_3;
  reg                 io_A_Valid_5_delay_16_2;
  reg                 io_A_Valid_5_delay_17_1;
  reg                 io_A_Valid_5_delay_18;
  reg                 io_B_Valid_18_delay_1_4;
  reg                 io_B_Valid_18_delay_2_3;
  reg                 io_B_Valid_18_delay_3_2;
  reg                 io_B_Valid_18_delay_4_1;
  reg                 io_B_Valid_18_delay_5;
  reg                 io_A_Valid_5_delay_1_18;
  reg                 io_A_Valid_5_delay_2_17;
  reg                 io_A_Valid_5_delay_3_16;
  reg                 io_A_Valid_5_delay_4_15;
  reg                 io_A_Valid_5_delay_5_14;
  reg                 io_A_Valid_5_delay_6_13;
  reg                 io_A_Valid_5_delay_7_12;
  reg                 io_A_Valid_5_delay_8_11;
  reg                 io_A_Valid_5_delay_9_10;
  reg                 io_A_Valid_5_delay_10_9;
  reg                 io_A_Valid_5_delay_11_8;
  reg                 io_A_Valid_5_delay_12_7;
  reg                 io_A_Valid_5_delay_13_6;
  reg                 io_A_Valid_5_delay_14_5;
  reg                 io_A_Valid_5_delay_15_4;
  reg                 io_A_Valid_5_delay_16_3;
  reg                 io_A_Valid_5_delay_17_2;
  reg                 io_A_Valid_5_delay_18_1;
  reg                 io_A_Valid_5_delay_19;
  reg                 io_B_Valid_19_delay_1_4;
  reg                 io_B_Valid_19_delay_2_3;
  reg                 io_B_Valid_19_delay_3_2;
  reg                 io_B_Valid_19_delay_4_1;
  reg                 io_B_Valid_19_delay_5;
  reg                 io_A_Valid_5_delay_1_19;
  reg                 io_A_Valid_5_delay_2_18;
  reg                 io_A_Valid_5_delay_3_17;
  reg                 io_A_Valid_5_delay_4_16;
  reg                 io_A_Valid_5_delay_5_15;
  reg                 io_A_Valid_5_delay_6_14;
  reg                 io_A_Valid_5_delay_7_13;
  reg                 io_A_Valid_5_delay_8_12;
  reg                 io_A_Valid_5_delay_9_11;
  reg                 io_A_Valid_5_delay_10_10;
  reg                 io_A_Valid_5_delay_11_9;
  reg                 io_A_Valid_5_delay_12_8;
  reg                 io_A_Valid_5_delay_13_7;
  reg                 io_A_Valid_5_delay_14_6;
  reg                 io_A_Valid_5_delay_15_5;
  reg                 io_A_Valid_5_delay_16_4;
  reg                 io_A_Valid_5_delay_17_3;
  reg                 io_A_Valid_5_delay_18_2;
  reg                 io_A_Valid_5_delay_19_1;
  reg                 io_A_Valid_5_delay_20;
  reg                 io_B_Valid_20_delay_1_4;
  reg                 io_B_Valid_20_delay_2_3;
  reg                 io_B_Valid_20_delay_3_2;
  reg                 io_B_Valid_20_delay_4_1;
  reg                 io_B_Valid_20_delay_5;
  reg                 io_A_Valid_5_delay_1_20;
  reg                 io_A_Valid_5_delay_2_19;
  reg                 io_A_Valid_5_delay_3_18;
  reg                 io_A_Valid_5_delay_4_17;
  reg                 io_A_Valid_5_delay_5_16;
  reg                 io_A_Valid_5_delay_6_15;
  reg                 io_A_Valid_5_delay_7_14;
  reg                 io_A_Valid_5_delay_8_13;
  reg                 io_A_Valid_5_delay_9_12;
  reg                 io_A_Valid_5_delay_10_11;
  reg                 io_A_Valid_5_delay_11_10;
  reg                 io_A_Valid_5_delay_12_9;
  reg                 io_A_Valid_5_delay_13_8;
  reg                 io_A_Valid_5_delay_14_7;
  reg                 io_A_Valid_5_delay_15_6;
  reg                 io_A_Valid_5_delay_16_5;
  reg                 io_A_Valid_5_delay_17_4;
  reg                 io_A_Valid_5_delay_18_3;
  reg                 io_A_Valid_5_delay_19_2;
  reg                 io_A_Valid_5_delay_20_1;
  reg                 io_A_Valid_5_delay_21;
  reg                 io_B_Valid_21_delay_1_4;
  reg                 io_B_Valid_21_delay_2_3;
  reg                 io_B_Valid_21_delay_3_2;
  reg                 io_B_Valid_21_delay_4_1;
  reg                 io_B_Valid_21_delay_5;
  reg                 io_A_Valid_5_delay_1_21;
  reg                 io_A_Valid_5_delay_2_20;
  reg                 io_A_Valid_5_delay_3_19;
  reg                 io_A_Valid_5_delay_4_18;
  reg                 io_A_Valid_5_delay_5_17;
  reg                 io_A_Valid_5_delay_6_16;
  reg                 io_A_Valid_5_delay_7_15;
  reg                 io_A_Valid_5_delay_8_14;
  reg                 io_A_Valid_5_delay_9_13;
  reg                 io_A_Valid_5_delay_10_12;
  reg                 io_A_Valid_5_delay_11_11;
  reg                 io_A_Valid_5_delay_12_10;
  reg                 io_A_Valid_5_delay_13_9;
  reg                 io_A_Valid_5_delay_14_8;
  reg                 io_A_Valid_5_delay_15_7;
  reg                 io_A_Valid_5_delay_16_6;
  reg                 io_A_Valid_5_delay_17_5;
  reg                 io_A_Valid_5_delay_18_4;
  reg                 io_A_Valid_5_delay_19_3;
  reg                 io_A_Valid_5_delay_20_2;
  reg                 io_A_Valid_5_delay_21_1;
  reg                 io_A_Valid_5_delay_22;
  reg                 io_B_Valid_22_delay_1_4;
  reg                 io_B_Valid_22_delay_2_3;
  reg                 io_B_Valid_22_delay_3_2;
  reg                 io_B_Valid_22_delay_4_1;
  reg                 io_B_Valid_22_delay_5;
  reg                 io_A_Valid_5_delay_1_22;
  reg                 io_A_Valid_5_delay_2_21;
  reg                 io_A_Valid_5_delay_3_20;
  reg                 io_A_Valid_5_delay_4_19;
  reg                 io_A_Valid_5_delay_5_18;
  reg                 io_A_Valid_5_delay_6_17;
  reg                 io_A_Valid_5_delay_7_16;
  reg                 io_A_Valid_5_delay_8_15;
  reg                 io_A_Valid_5_delay_9_14;
  reg                 io_A_Valid_5_delay_10_13;
  reg                 io_A_Valid_5_delay_11_12;
  reg                 io_A_Valid_5_delay_12_11;
  reg                 io_A_Valid_5_delay_13_10;
  reg                 io_A_Valid_5_delay_14_9;
  reg                 io_A_Valid_5_delay_15_8;
  reg                 io_A_Valid_5_delay_16_7;
  reg                 io_A_Valid_5_delay_17_6;
  reg                 io_A_Valid_5_delay_18_5;
  reg                 io_A_Valid_5_delay_19_4;
  reg                 io_A_Valid_5_delay_20_3;
  reg                 io_A_Valid_5_delay_21_2;
  reg                 io_A_Valid_5_delay_22_1;
  reg                 io_A_Valid_5_delay_23;
  reg                 io_B_Valid_23_delay_1_4;
  reg                 io_B_Valid_23_delay_2_3;
  reg                 io_B_Valid_23_delay_3_2;
  reg                 io_B_Valid_23_delay_4_1;
  reg                 io_B_Valid_23_delay_5;
  reg                 io_A_Valid_5_delay_1_23;
  reg                 io_A_Valid_5_delay_2_22;
  reg                 io_A_Valid_5_delay_3_21;
  reg                 io_A_Valid_5_delay_4_20;
  reg                 io_A_Valid_5_delay_5_19;
  reg                 io_A_Valid_5_delay_6_18;
  reg                 io_A_Valid_5_delay_7_17;
  reg                 io_A_Valid_5_delay_8_16;
  reg                 io_A_Valid_5_delay_9_15;
  reg                 io_A_Valid_5_delay_10_14;
  reg                 io_A_Valid_5_delay_11_13;
  reg                 io_A_Valid_5_delay_12_12;
  reg                 io_A_Valid_5_delay_13_11;
  reg                 io_A_Valid_5_delay_14_10;
  reg                 io_A_Valid_5_delay_15_9;
  reg                 io_A_Valid_5_delay_16_8;
  reg                 io_A_Valid_5_delay_17_7;
  reg                 io_A_Valid_5_delay_18_6;
  reg                 io_A_Valid_5_delay_19_5;
  reg                 io_A_Valid_5_delay_20_4;
  reg                 io_A_Valid_5_delay_21_3;
  reg                 io_A_Valid_5_delay_22_2;
  reg                 io_A_Valid_5_delay_23_1;
  reg                 io_A_Valid_5_delay_24;
  reg                 io_B_Valid_24_delay_1_4;
  reg                 io_B_Valid_24_delay_2_3;
  reg                 io_B_Valid_24_delay_3_2;
  reg                 io_B_Valid_24_delay_4_1;
  reg                 io_B_Valid_24_delay_5;
  reg                 io_A_Valid_5_delay_1_24;
  reg                 io_A_Valid_5_delay_2_23;
  reg                 io_A_Valid_5_delay_3_22;
  reg                 io_A_Valid_5_delay_4_21;
  reg                 io_A_Valid_5_delay_5_20;
  reg                 io_A_Valid_5_delay_6_19;
  reg                 io_A_Valid_5_delay_7_18;
  reg                 io_A_Valid_5_delay_8_17;
  reg                 io_A_Valid_5_delay_9_16;
  reg                 io_A_Valid_5_delay_10_15;
  reg                 io_A_Valid_5_delay_11_14;
  reg                 io_A_Valid_5_delay_12_13;
  reg                 io_A_Valid_5_delay_13_12;
  reg                 io_A_Valid_5_delay_14_11;
  reg                 io_A_Valid_5_delay_15_10;
  reg                 io_A_Valid_5_delay_16_9;
  reg                 io_A_Valid_5_delay_17_8;
  reg                 io_A_Valid_5_delay_18_7;
  reg                 io_A_Valid_5_delay_19_6;
  reg                 io_A_Valid_5_delay_20_5;
  reg                 io_A_Valid_5_delay_21_4;
  reg                 io_A_Valid_5_delay_22_3;
  reg                 io_A_Valid_5_delay_23_2;
  reg                 io_A_Valid_5_delay_24_1;
  reg                 io_A_Valid_5_delay_25;
  reg                 io_B_Valid_25_delay_1_4;
  reg                 io_B_Valid_25_delay_2_3;
  reg                 io_B_Valid_25_delay_3_2;
  reg                 io_B_Valid_25_delay_4_1;
  reg                 io_B_Valid_25_delay_5;
  reg                 io_A_Valid_5_delay_1_25;
  reg                 io_A_Valid_5_delay_2_24;
  reg                 io_A_Valid_5_delay_3_23;
  reg                 io_A_Valid_5_delay_4_22;
  reg                 io_A_Valid_5_delay_5_21;
  reg                 io_A_Valid_5_delay_6_20;
  reg                 io_A_Valid_5_delay_7_19;
  reg                 io_A_Valid_5_delay_8_18;
  reg                 io_A_Valid_5_delay_9_17;
  reg                 io_A_Valid_5_delay_10_16;
  reg                 io_A_Valid_5_delay_11_15;
  reg                 io_A_Valid_5_delay_12_14;
  reg                 io_A_Valid_5_delay_13_13;
  reg                 io_A_Valid_5_delay_14_12;
  reg                 io_A_Valid_5_delay_15_11;
  reg                 io_A_Valid_5_delay_16_10;
  reg                 io_A_Valid_5_delay_17_9;
  reg                 io_A_Valid_5_delay_18_8;
  reg                 io_A_Valid_5_delay_19_7;
  reg                 io_A_Valid_5_delay_20_6;
  reg                 io_A_Valid_5_delay_21_5;
  reg                 io_A_Valid_5_delay_22_4;
  reg                 io_A_Valid_5_delay_23_3;
  reg                 io_A_Valid_5_delay_24_2;
  reg                 io_A_Valid_5_delay_25_1;
  reg                 io_A_Valid_5_delay_26;
  reg                 io_B_Valid_26_delay_1_4;
  reg                 io_B_Valid_26_delay_2_3;
  reg                 io_B_Valid_26_delay_3_2;
  reg                 io_B_Valid_26_delay_4_1;
  reg                 io_B_Valid_26_delay_5;
  reg                 io_A_Valid_5_delay_1_26;
  reg                 io_A_Valid_5_delay_2_25;
  reg                 io_A_Valid_5_delay_3_24;
  reg                 io_A_Valid_5_delay_4_23;
  reg                 io_A_Valid_5_delay_5_22;
  reg                 io_A_Valid_5_delay_6_21;
  reg                 io_A_Valid_5_delay_7_20;
  reg                 io_A_Valid_5_delay_8_19;
  reg                 io_A_Valid_5_delay_9_18;
  reg                 io_A_Valid_5_delay_10_17;
  reg                 io_A_Valid_5_delay_11_16;
  reg                 io_A_Valid_5_delay_12_15;
  reg                 io_A_Valid_5_delay_13_14;
  reg                 io_A_Valid_5_delay_14_13;
  reg                 io_A_Valid_5_delay_15_12;
  reg                 io_A_Valid_5_delay_16_11;
  reg                 io_A_Valid_5_delay_17_10;
  reg                 io_A_Valid_5_delay_18_9;
  reg                 io_A_Valid_5_delay_19_8;
  reg                 io_A_Valid_5_delay_20_7;
  reg                 io_A_Valid_5_delay_21_6;
  reg                 io_A_Valid_5_delay_22_5;
  reg                 io_A_Valid_5_delay_23_4;
  reg                 io_A_Valid_5_delay_24_3;
  reg                 io_A_Valid_5_delay_25_2;
  reg                 io_A_Valid_5_delay_26_1;
  reg                 io_A_Valid_5_delay_27;
  reg                 io_B_Valid_27_delay_1_4;
  reg                 io_B_Valid_27_delay_2_3;
  reg                 io_B_Valid_27_delay_3_2;
  reg                 io_B_Valid_27_delay_4_1;
  reg                 io_B_Valid_27_delay_5;
  reg                 io_A_Valid_5_delay_1_27;
  reg                 io_A_Valid_5_delay_2_26;
  reg                 io_A_Valid_5_delay_3_25;
  reg                 io_A_Valid_5_delay_4_24;
  reg                 io_A_Valid_5_delay_5_23;
  reg                 io_A_Valid_5_delay_6_22;
  reg                 io_A_Valid_5_delay_7_21;
  reg                 io_A_Valid_5_delay_8_20;
  reg                 io_A_Valid_5_delay_9_19;
  reg                 io_A_Valid_5_delay_10_18;
  reg                 io_A_Valid_5_delay_11_17;
  reg                 io_A_Valid_5_delay_12_16;
  reg                 io_A_Valid_5_delay_13_15;
  reg                 io_A_Valid_5_delay_14_14;
  reg                 io_A_Valid_5_delay_15_13;
  reg                 io_A_Valid_5_delay_16_12;
  reg                 io_A_Valid_5_delay_17_11;
  reg                 io_A_Valid_5_delay_18_10;
  reg                 io_A_Valid_5_delay_19_9;
  reg                 io_A_Valid_5_delay_20_8;
  reg                 io_A_Valid_5_delay_21_7;
  reg                 io_A_Valid_5_delay_22_6;
  reg                 io_A_Valid_5_delay_23_5;
  reg                 io_A_Valid_5_delay_24_4;
  reg                 io_A_Valid_5_delay_25_3;
  reg                 io_A_Valid_5_delay_26_2;
  reg                 io_A_Valid_5_delay_27_1;
  reg                 io_A_Valid_5_delay_28;
  reg                 io_B_Valid_28_delay_1_4;
  reg                 io_B_Valid_28_delay_2_3;
  reg                 io_B_Valid_28_delay_3_2;
  reg                 io_B_Valid_28_delay_4_1;
  reg                 io_B_Valid_28_delay_5;
  reg                 io_A_Valid_5_delay_1_28;
  reg                 io_A_Valid_5_delay_2_27;
  reg                 io_A_Valid_5_delay_3_26;
  reg                 io_A_Valid_5_delay_4_25;
  reg                 io_A_Valid_5_delay_5_24;
  reg                 io_A_Valid_5_delay_6_23;
  reg                 io_A_Valid_5_delay_7_22;
  reg                 io_A_Valid_5_delay_8_21;
  reg                 io_A_Valid_5_delay_9_20;
  reg                 io_A_Valid_5_delay_10_19;
  reg                 io_A_Valid_5_delay_11_18;
  reg                 io_A_Valid_5_delay_12_17;
  reg                 io_A_Valid_5_delay_13_16;
  reg                 io_A_Valid_5_delay_14_15;
  reg                 io_A_Valid_5_delay_15_14;
  reg                 io_A_Valid_5_delay_16_13;
  reg                 io_A_Valid_5_delay_17_12;
  reg                 io_A_Valid_5_delay_18_11;
  reg                 io_A_Valid_5_delay_19_10;
  reg                 io_A_Valid_5_delay_20_9;
  reg                 io_A_Valid_5_delay_21_8;
  reg                 io_A_Valid_5_delay_22_7;
  reg                 io_A_Valid_5_delay_23_6;
  reg                 io_A_Valid_5_delay_24_5;
  reg                 io_A_Valid_5_delay_25_4;
  reg                 io_A_Valid_5_delay_26_3;
  reg                 io_A_Valid_5_delay_27_2;
  reg                 io_A_Valid_5_delay_28_1;
  reg                 io_A_Valid_5_delay_29;
  reg                 io_B_Valid_29_delay_1_4;
  reg                 io_B_Valid_29_delay_2_3;
  reg                 io_B_Valid_29_delay_3_2;
  reg                 io_B_Valid_29_delay_4_1;
  reg                 io_B_Valid_29_delay_5;
  reg                 io_A_Valid_5_delay_1_29;
  reg                 io_A_Valid_5_delay_2_28;
  reg                 io_A_Valid_5_delay_3_27;
  reg                 io_A_Valid_5_delay_4_26;
  reg                 io_A_Valid_5_delay_5_25;
  reg                 io_A_Valid_5_delay_6_24;
  reg                 io_A_Valid_5_delay_7_23;
  reg                 io_A_Valid_5_delay_8_22;
  reg                 io_A_Valid_5_delay_9_21;
  reg                 io_A_Valid_5_delay_10_20;
  reg                 io_A_Valid_5_delay_11_19;
  reg                 io_A_Valid_5_delay_12_18;
  reg                 io_A_Valid_5_delay_13_17;
  reg                 io_A_Valid_5_delay_14_16;
  reg                 io_A_Valid_5_delay_15_15;
  reg                 io_A_Valid_5_delay_16_14;
  reg                 io_A_Valid_5_delay_17_13;
  reg                 io_A_Valid_5_delay_18_12;
  reg                 io_A_Valid_5_delay_19_11;
  reg                 io_A_Valid_5_delay_20_10;
  reg                 io_A_Valid_5_delay_21_9;
  reg                 io_A_Valid_5_delay_22_8;
  reg                 io_A_Valid_5_delay_23_7;
  reg                 io_A_Valid_5_delay_24_6;
  reg                 io_A_Valid_5_delay_25_5;
  reg                 io_A_Valid_5_delay_26_4;
  reg                 io_A_Valid_5_delay_27_3;
  reg                 io_A_Valid_5_delay_28_2;
  reg                 io_A_Valid_5_delay_29_1;
  reg                 io_A_Valid_5_delay_30;
  reg                 io_B_Valid_30_delay_1_4;
  reg                 io_B_Valid_30_delay_2_3;
  reg                 io_B_Valid_30_delay_3_2;
  reg                 io_B_Valid_30_delay_4_1;
  reg                 io_B_Valid_30_delay_5;
  reg                 io_A_Valid_5_delay_1_30;
  reg                 io_A_Valid_5_delay_2_29;
  reg                 io_A_Valid_5_delay_3_28;
  reg                 io_A_Valid_5_delay_4_27;
  reg                 io_A_Valid_5_delay_5_26;
  reg                 io_A_Valid_5_delay_6_25;
  reg                 io_A_Valid_5_delay_7_24;
  reg                 io_A_Valid_5_delay_8_23;
  reg                 io_A_Valid_5_delay_9_22;
  reg                 io_A_Valid_5_delay_10_21;
  reg                 io_A_Valid_5_delay_11_20;
  reg                 io_A_Valid_5_delay_12_19;
  reg                 io_A_Valid_5_delay_13_18;
  reg                 io_A_Valid_5_delay_14_17;
  reg                 io_A_Valid_5_delay_15_16;
  reg                 io_A_Valid_5_delay_16_15;
  reg                 io_A_Valid_5_delay_17_14;
  reg                 io_A_Valid_5_delay_18_13;
  reg                 io_A_Valid_5_delay_19_12;
  reg                 io_A_Valid_5_delay_20_11;
  reg                 io_A_Valid_5_delay_21_10;
  reg                 io_A_Valid_5_delay_22_9;
  reg                 io_A_Valid_5_delay_23_8;
  reg                 io_A_Valid_5_delay_24_7;
  reg                 io_A_Valid_5_delay_25_6;
  reg                 io_A_Valid_5_delay_26_5;
  reg                 io_A_Valid_5_delay_27_4;
  reg                 io_A_Valid_5_delay_28_3;
  reg                 io_A_Valid_5_delay_29_2;
  reg                 io_A_Valid_5_delay_30_1;
  reg                 io_A_Valid_5_delay_31;
  reg                 io_B_Valid_31_delay_1_4;
  reg                 io_B_Valid_31_delay_2_3;
  reg                 io_B_Valid_31_delay_3_2;
  reg                 io_B_Valid_31_delay_4_1;
  reg                 io_B_Valid_31_delay_5;
  reg                 io_A_Valid_5_delay_1_31;
  reg                 io_A_Valid_5_delay_2_30;
  reg                 io_A_Valid_5_delay_3_29;
  reg                 io_A_Valid_5_delay_4_28;
  reg                 io_A_Valid_5_delay_5_27;
  reg                 io_A_Valid_5_delay_6_26;
  reg                 io_A_Valid_5_delay_7_25;
  reg                 io_A_Valid_5_delay_8_24;
  reg                 io_A_Valid_5_delay_9_23;
  reg                 io_A_Valid_5_delay_10_22;
  reg                 io_A_Valid_5_delay_11_21;
  reg                 io_A_Valid_5_delay_12_20;
  reg                 io_A_Valid_5_delay_13_19;
  reg                 io_A_Valid_5_delay_14_18;
  reg                 io_A_Valid_5_delay_15_17;
  reg                 io_A_Valid_5_delay_16_16;
  reg                 io_A_Valid_5_delay_17_15;
  reg                 io_A_Valid_5_delay_18_14;
  reg                 io_A_Valid_5_delay_19_13;
  reg                 io_A_Valid_5_delay_20_12;
  reg                 io_A_Valid_5_delay_21_11;
  reg                 io_A_Valid_5_delay_22_10;
  reg                 io_A_Valid_5_delay_23_9;
  reg                 io_A_Valid_5_delay_24_8;
  reg                 io_A_Valid_5_delay_25_7;
  reg                 io_A_Valid_5_delay_26_6;
  reg                 io_A_Valid_5_delay_27_5;
  reg                 io_A_Valid_5_delay_28_4;
  reg                 io_A_Valid_5_delay_29_3;
  reg                 io_A_Valid_5_delay_30_2;
  reg                 io_A_Valid_5_delay_31_1;
  reg                 io_A_Valid_5_delay_32;
  reg                 io_B_Valid_32_delay_1_4;
  reg                 io_B_Valid_32_delay_2_3;
  reg                 io_B_Valid_32_delay_3_2;
  reg                 io_B_Valid_32_delay_4_1;
  reg                 io_B_Valid_32_delay_5;
  reg                 io_A_Valid_5_delay_1_32;
  reg                 io_A_Valid_5_delay_2_31;
  reg                 io_A_Valid_5_delay_3_30;
  reg                 io_A_Valid_5_delay_4_29;
  reg                 io_A_Valid_5_delay_5_28;
  reg                 io_A_Valid_5_delay_6_27;
  reg                 io_A_Valid_5_delay_7_26;
  reg                 io_A_Valid_5_delay_8_25;
  reg                 io_A_Valid_5_delay_9_24;
  reg                 io_A_Valid_5_delay_10_23;
  reg                 io_A_Valid_5_delay_11_22;
  reg                 io_A_Valid_5_delay_12_21;
  reg                 io_A_Valid_5_delay_13_20;
  reg                 io_A_Valid_5_delay_14_19;
  reg                 io_A_Valid_5_delay_15_18;
  reg                 io_A_Valid_5_delay_16_17;
  reg                 io_A_Valid_5_delay_17_16;
  reg                 io_A_Valid_5_delay_18_15;
  reg                 io_A_Valid_5_delay_19_14;
  reg                 io_A_Valid_5_delay_20_13;
  reg                 io_A_Valid_5_delay_21_12;
  reg                 io_A_Valid_5_delay_22_11;
  reg                 io_A_Valid_5_delay_23_10;
  reg                 io_A_Valid_5_delay_24_9;
  reg                 io_A_Valid_5_delay_25_8;
  reg                 io_A_Valid_5_delay_26_7;
  reg                 io_A_Valid_5_delay_27_6;
  reg                 io_A_Valid_5_delay_28_5;
  reg                 io_A_Valid_5_delay_29_4;
  reg                 io_A_Valid_5_delay_30_3;
  reg                 io_A_Valid_5_delay_31_2;
  reg                 io_A_Valid_5_delay_32_1;
  reg                 io_A_Valid_5_delay_33;
  reg                 io_B_Valid_33_delay_1_4;
  reg                 io_B_Valid_33_delay_2_3;
  reg                 io_B_Valid_33_delay_3_2;
  reg                 io_B_Valid_33_delay_4_1;
  reg                 io_B_Valid_33_delay_5;
  reg                 io_A_Valid_5_delay_1_33;
  reg                 io_A_Valid_5_delay_2_32;
  reg                 io_A_Valid_5_delay_3_31;
  reg                 io_A_Valid_5_delay_4_30;
  reg                 io_A_Valid_5_delay_5_29;
  reg                 io_A_Valid_5_delay_6_28;
  reg                 io_A_Valid_5_delay_7_27;
  reg                 io_A_Valid_5_delay_8_26;
  reg                 io_A_Valid_5_delay_9_25;
  reg                 io_A_Valid_5_delay_10_24;
  reg                 io_A_Valid_5_delay_11_23;
  reg                 io_A_Valid_5_delay_12_22;
  reg                 io_A_Valid_5_delay_13_21;
  reg                 io_A_Valid_5_delay_14_20;
  reg                 io_A_Valid_5_delay_15_19;
  reg                 io_A_Valid_5_delay_16_18;
  reg                 io_A_Valid_5_delay_17_17;
  reg                 io_A_Valid_5_delay_18_16;
  reg                 io_A_Valid_5_delay_19_15;
  reg                 io_A_Valid_5_delay_20_14;
  reg                 io_A_Valid_5_delay_21_13;
  reg                 io_A_Valid_5_delay_22_12;
  reg                 io_A_Valid_5_delay_23_11;
  reg                 io_A_Valid_5_delay_24_10;
  reg                 io_A_Valid_5_delay_25_9;
  reg                 io_A_Valid_5_delay_26_8;
  reg                 io_A_Valid_5_delay_27_7;
  reg                 io_A_Valid_5_delay_28_6;
  reg                 io_A_Valid_5_delay_29_5;
  reg                 io_A_Valid_5_delay_30_4;
  reg                 io_A_Valid_5_delay_31_3;
  reg                 io_A_Valid_5_delay_32_2;
  reg                 io_A_Valid_5_delay_33_1;
  reg                 io_A_Valid_5_delay_34;
  reg                 io_B_Valid_34_delay_1_4;
  reg                 io_B_Valid_34_delay_2_3;
  reg                 io_B_Valid_34_delay_3_2;
  reg                 io_B_Valid_34_delay_4_1;
  reg                 io_B_Valid_34_delay_5;
  reg                 io_A_Valid_5_delay_1_34;
  reg                 io_A_Valid_5_delay_2_33;
  reg                 io_A_Valid_5_delay_3_32;
  reg                 io_A_Valid_5_delay_4_31;
  reg                 io_A_Valid_5_delay_5_30;
  reg                 io_A_Valid_5_delay_6_29;
  reg                 io_A_Valid_5_delay_7_28;
  reg                 io_A_Valid_5_delay_8_27;
  reg                 io_A_Valid_5_delay_9_26;
  reg                 io_A_Valid_5_delay_10_25;
  reg                 io_A_Valid_5_delay_11_24;
  reg                 io_A_Valid_5_delay_12_23;
  reg                 io_A_Valid_5_delay_13_22;
  reg                 io_A_Valid_5_delay_14_21;
  reg                 io_A_Valid_5_delay_15_20;
  reg                 io_A_Valid_5_delay_16_19;
  reg                 io_A_Valid_5_delay_17_18;
  reg                 io_A_Valid_5_delay_18_17;
  reg                 io_A_Valid_5_delay_19_16;
  reg                 io_A_Valid_5_delay_20_15;
  reg                 io_A_Valid_5_delay_21_14;
  reg                 io_A_Valid_5_delay_22_13;
  reg                 io_A_Valid_5_delay_23_12;
  reg                 io_A_Valid_5_delay_24_11;
  reg                 io_A_Valid_5_delay_25_10;
  reg                 io_A_Valid_5_delay_26_9;
  reg                 io_A_Valid_5_delay_27_8;
  reg                 io_A_Valid_5_delay_28_7;
  reg                 io_A_Valid_5_delay_29_6;
  reg                 io_A_Valid_5_delay_30_5;
  reg                 io_A_Valid_5_delay_31_4;
  reg                 io_A_Valid_5_delay_32_3;
  reg                 io_A_Valid_5_delay_33_2;
  reg                 io_A_Valid_5_delay_34_1;
  reg                 io_A_Valid_5_delay_35;
  reg                 io_B_Valid_35_delay_1_4;
  reg                 io_B_Valid_35_delay_2_3;
  reg                 io_B_Valid_35_delay_3_2;
  reg                 io_B_Valid_35_delay_4_1;
  reg                 io_B_Valid_35_delay_5;
  reg                 io_A_Valid_5_delay_1_35;
  reg                 io_A_Valid_5_delay_2_34;
  reg                 io_A_Valid_5_delay_3_33;
  reg                 io_A_Valid_5_delay_4_32;
  reg                 io_A_Valid_5_delay_5_31;
  reg                 io_A_Valid_5_delay_6_30;
  reg                 io_A_Valid_5_delay_7_29;
  reg                 io_A_Valid_5_delay_8_28;
  reg                 io_A_Valid_5_delay_9_27;
  reg                 io_A_Valid_5_delay_10_26;
  reg                 io_A_Valid_5_delay_11_25;
  reg                 io_A_Valid_5_delay_12_24;
  reg                 io_A_Valid_5_delay_13_23;
  reg                 io_A_Valid_5_delay_14_22;
  reg                 io_A_Valid_5_delay_15_21;
  reg                 io_A_Valid_5_delay_16_20;
  reg                 io_A_Valid_5_delay_17_19;
  reg                 io_A_Valid_5_delay_18_18;
  reg                 io_A_Valid_5_delay_19_17;
  reg                 io_A_Valid_5_delay_20_16;
  reg                 io_A_Valid_5_delay_21_15;
  reg                 io_A_Valid_5_delay_22_14;
  reg                 io_A_Valid_5_delay_23_13;
  reg                 io_A_Valid_5_delay_24_12;
  reg                 io_A_Valid_5_delay_25_11;
  reg                 io_A_Valid_5_delay_26_10;
  reg                 io_A_Valid_5_delay_27_9;
  reg                 io_A_Valid_5_delay_28_8;
  reg                 io_A_Valid_5_delay_29_7;
  reg                 io_A_Valid_5_delay_30_6;
  reg                 io_A_Valid_5_delay_31_5;
  reg                 io_A_Valid_5_delay_32_4;
  reg                 io_A_Valid_5_delay_33_3;
  reg                 io_A_Valid_5_delay_34_2;
  reg                 io_A_Valid_5_delay_35_1;
  reg                 io_A_Valid_5_delay_36;
  reg                 io_B_Valid_36_delay_1_4;
  reg                 io_B_Valid_36_delay_2_3;
  reg                 io_B_Valid_36_delay_3_2;
  reg                 io_B_Valid_36_delay_4_1;
  reg                 io_B_Valid_36_delay_5;
  reg                 io_A_Valid_5_delay_1_36;
  reg                 io_A_Valid_5_delay_2_35;
  reg                 io_A_Valid_5_delay_3_34;
  reg                 io_A_Valid_5_delay_4_33;
  reg                 io_A_Valid_5_delay_5_32;
  reg                 io_A_Valid_5_delay_6_31;
  reg                 io_A_Valid_5_delay_7_30;
  reg                 io_A_Valid_5_delay_8_29;
  reg                 io_A_Valid_5_delay_9_28;
  reg                 io_A_Valid_5_delay_10_27;
  reg                 io_A_Valid_5_delay_11_26;
  reg                 io_A_Valid_5_delay_12_25;
  reg                 io_A_Valid_5_delay_13_24;
  reg                 io_A_Valid_5_delay_14_23;
  reg                 io_A_Valid_5_delay_15_22;
  reg                 io_A_Valid_5_delay_16_21;
  reg                 io_A_Valid_5_delay_17_20;
  reg                 io_A_Valid_5_delay_18_19;
  reg                 io_A_Valid_5_delay_19_18;
  reg                 io_A_Valid_5_delay_20_17;
  reg                 io_A_Valid_5_delay_21_16;
  reg                 io_A_Valid_5_delay_22_15;
  reg                 io_A_Valid_5_delay_23_14;
  reg                 io_A_Valid_5_delay_24_13;
  reg                 io_A_Valid_5_delay_25_12;
  reg                 io_A_Valid_5_delay_26_11;
  reg                 io_A_Valid_5_delay_27_10;
  reg                 io_A_Valid_5_delay_28_9;
  reg                 io_A_Valid_5_delay_29_8;
  reg                 io_A_Valid_5_delay_30_7;
  reg                 io_A_Valid_5_delay_31_6;
  reg                 io_A_Valid_5_delay_32_5;
  reg                 io_A_Valid_5_delay_33_4;
  reg                 io_A_Valid_5_delay_34_3;
  reg                 io_A_Valid_5_delay_35_2;
  reg                 io_A_Valid_5_delay_36_1;
  reg                 io_A_Valid_5_delay_37;
  reg                 io_B_Valid_37_delay_1_4;
  reg                 io_B_Valid_37_delay_2_3;
  reg                 io_B_Valid_37_delay_3_2;
  reg                 io_B_Valid_37_delay_4_1;
  reg                 io_B_Valid_37_delay_5;
  reg                 io_A_Valid_5_delay_1_37;
  reg                 io_A_Valid_5_delay_2_36;
  reg                 io_A_Valid_5_delay_3_35;
  reg                 io_A_Valid_5_delay_4_34;
  reg                 io_A_Valid_5_delay_5_33;
  reg                 io_A_Valid_5_delay_6_32;
  reg                 io_A_Valid_5_delay_7_31;
  reg                 io_A_Valid_5_delay_8_30;
  reg                 io_A_Valid_5_delay_9_29;
  reg                 io_A_Valid_5_delay_10_28;
  reg                 io_A_Valid_5_delay_11_27;
  reg                 io_A_Valid_5_delay_12_26;
  reg                 io_A_Valid_5_delay_13_25;
  reg                 io_A_Valid_5_delay_14_24;
  reg                 io_A_Valid_5_delay_15_23;
  reg                 io_A_Valid_5_delay_16_22;
  reg                 io_A_Valid_5_delay_17_21;
  reg                 io_A_Valid_5_delay_18_20;
  reg                 io_A_Valid_5_delay_19_19;
  reg                 io_A_Valid_5_delay_20_18;
  reg                 io_A_Valid_5_delay_21_17;
  reg                 io_A_Valid_5_delay_22_16;
  reg                 io_A_Valid_5_delay_23_15;
  reg                 io_A_Valid_5_delay_24_14;
  reg                 io_A_Valid_5_delay_25_13;
  reg                 io_A_Valid_5_delay_26_12;
  reg                 io_A_Valid_5_delay_27_11;
  reg                 io_A_Valid_5_delay_28_10;
  reg                 io_A_Valid_5_delay_29_9;
  reg                 io_A_Valid_5_delay_30_8;
  reg                 io_A_Valid_5_delay_31_7;
  reg                 io_A_Valid_5_delay_32_6;
  reg                 io_A_Valid_5_delay_33_5;
  reg                 io_A_Valid_5_delay_34_4;
  reg                 io_A_Valid_5_delay_35_3;
  reg                 io_A_Valid_5_delay_36_2;
  reg                 io_A_Valid_5_delay_37_1;
  reg                 io_A_Valid_5_delay_38;
  reg                 io_B_Valid_38_delay_1_4;
  reg                 io_B_Valid_38_delay_2_3;
  reg                 io_B_Valid_38_delay_3_2;
  reg                 io_B_Valid_38_delay_4_1;
  reg                 io_B_Valid_38_delay_5;
  reg                 io_A_Valid_5_delay_1_38;
  reg                 io_A_Valid_5_delay_2_37;
  reg                 io_A_Valid_5_delay_3_36;
  reg                 io_A_Valid_5_delay_4_35;
  reg                 io_A_Valid_5_delay_5_34;
  reg                 io_A_Valid_5_delay_6_33;
  reg                 io_A_Valid_5_delay_7_32;
  reg                 io_A_Valid_5_delay_8_31;
  reg                 io_A_Valid_5_delay_9_30;
  reg                 io_A_Valid_5_delay_10_29;
  reg                 io_A_Valid_5_delay_11_28;
  reg                 io_A_Valid_5_delay_12_27;
  reg                 io_A_Valid_5_delay_13_26;
  reg                 io_A_Valid_5_delay_14_25;
  reg                 io_A_Valid_5_delay_15_24;
  reg                 io_A_Valid_5_delay_16_23;
  reg                 io_A_Valid_5_delay_17_22;
  reg                 io_A_Valid_5_delay_18_21;
  reg                 io_A_Valid_5_delay_19_20;
  reg                 io_A_Valid_5_delay_20_19;
  reg                 io_A_Valid_5_delay_21_18;
  reg                 io_A_Valid_5_delay_22_17;
  reg                 io_A_Valid_5_delay_23_16;
  reg                 io_A_Valid_5_delay_24_15;
  reg                 io_A_Valid_5_delay_25_14;
  reg                 io_A_Valid_5_delay_26_13;
  reg                 io_A_Valid_5_delay_27_12;
  reg                 io_A_Valid_5_delay_28_11;
  reg                 io_A_Valid_5_delay_29_10;
  reg                 io_A_Valid_5_delay_30_9;
  reg                 io_A_Valid_5_delay_31_8;
  reg                 io_A_Valid_5_delay_32_7;
  reg                 io_A_Valid_5_delay_33_6;
  reg                 io_A_Valid_5_delay_34_5;
  reg                 io_A_Valid_5_delay_35_4;
  reg                 io_A_Valid_5_delay_36_3;
  reg                 io_A_Valid_5_delay_37_2;
  reg                 io_A_Valid_5_delay_38_1;
  reg                 io_A_Valid_5_delay_39;
  reg                 io_B_Valid_39_delay_1_4;
  reg                 io_B_Valid_39_delay_2_3;
  reg                 io_B_Valid_39_delay_3_2;
  reg                 io_B_Valid_39_delay_4_1;
  reg                 io_B_Valid_39_delay_5;
  reg                 io_A_Valid_5_delay_1_39;
  reg                 io_A_Valid_5_delay_2_38;
  reg                 io_A_Valid_5_delay_3_37;
  reg                 io_A_Valid_5_delay_4_36;
  reg                 io_A_Valid_5_delay_5_35;
  reg                 io_A_Valid_5_delay_6_34;
  reg                 io_A_Valid_5_delay_7_33;
  reg                 io_A_Valid_5_delay_8_32;
  reg                 io_A_Valid_5_delay_9_31;
  reg                 io_A_Valid_5_delay_10_30;
  reg                 io_A_Valid_5_delay_11_29;
  reg                 io_A_Valid_5_delay_12_28;
  reg                 io_A_Valid_5_delay_13_27;
  reg                 io_A_Valid_5_delay_14_26;
  reg                 io_A_Valid_5_delay_15_25;
  reg                 io_A_Valid_5_delay_16_24;
  reg                 io_A_Valid_5_delay_17_23;
  reg                 io_A_Valid_5_delay_18_22;
  reg                 io_A_Valid_5_delay_19_21;
  reg                 io_A_Valid_5_delay_20_20;
  reg                 io_A_Valid_5_delay_21_19;
  reg                 io_A_Valid_5_delay_22_18;
  reg                 io_A_Valid_5_delay_23_17;
  reg                 io_A_Valid_5_delay_24_16;
  reg                 io_A_Valid_5_delay_25_15;
  reg                 io_A_Valid_5_delay_26_14;
  reg                 io_A_Valid_5_delay_27_13;
  reg                 io_A_Valid_5_delay_28_12;
  reg                 io_A_Valid_5_delay_29_11;
  reg                 io_A_Valid_5_delay_30_10;
  reg                 io_A_Valid_5_delay_31_9;
  reg                 io_A_Valid_5_delay_32_8;
  reg                 io_A_Valid_5_delay_33_7;
  reg                 io_A_Valid_5_delay_34_6;
  reg                 io_A_Valid_5_delay_35_5;
  reg                 io_A_Valid_5_delay_36_4;
  reg                 io_A_Valid_5_delay_37_3;
  reg                 io_A_Valid_5_delay_38_2;
  reg                 io_A_Valid_5_delay_39_1;
  reg                 io_A_Valid_5_delay_40;
  reg                 io_B_Valid_40_delay_1_4;
  reg                 io_B_Valid_40_delay_2_3;
  reg                 io_B_Valid_40_delay_3_2;
  reg                 io_B_Valid_40_delay_4_1;
  reg                 io_B_Valid_40_delay_5;
  reg                 io_A_Valid_5_delay_1_40;
  reg                 io_A_Valid_5_delay_2_39;
  reg                 io_A_Valid_5_delay_3_38;
  reg                 io_A_Valid_5_delay_4_37;
  reg                 io_A_Valid_5_delay_5_36;
  reg                 io_A_Valid_5_delay_6_35;
  reg                 io_A_Valid_5_delay_7_34;
  reg                 io_A_Valid_5_delay_8_33;
  reg                 io_A_Valid_5_delay_9_32;
  reg                 io_A_Valid_5_delay_10_31;
  reg                 io_A_Valid_5_delay_11_30;
  reg                 io_A_Valid_5_delay_12_29;
  reg                 io_A_Valid_5_delay_13_28;
  reg                 io_A_Valid_5_delay_14_27;
  reg                 io_A_Valid_5_delay_15_26;
  reg                 io_A_Valid_5_delay_16_25;
  reg                 io_A_Valid_5_delay_17_24;
  reg                 io_A_Valid_5_delay_18_23;
  reg                 io_A_Valid_5_delay_19_22;
  reg                 io_A_Valid_5_delay_20_21;
  reg                 io_A_Valid_5_delay_21_20;
  reg                 io_A_Valid_5_delay_22_19;
  reg                 io_A_Valid_5_delay_23_18;
  reg                 io_A_Valid_5_delay_24_17;
  reg                 io_A_Valid_5_delay_25_16;
  reg                 io_A_Valid_5_delay_26_15;
  reg                 io_A_Valid_5_delay_27_14;
  reg                 io_A_Valid_5_delay_28_13;
  reg                 io_A_Valid_5_delay_29_12;
  reg                 io_A_Valid_5_delay_30_11;
  reg                 io_A_Valid_5_delay_31_10;
  reg                 io_A_Valid_5_delay_32_9;
  reg                 io_A_Valid_5_delay_33_8;
  reg                 io_A_Valid_5_delay_34_7;
  reg                 io_A_Valid_5_delay_35_6;
  reg                 io_A_Valid_5_delay_36_5;
  reg                 io_A_Valid_5_delay_37_4;
  reg                 io_A_Valid_5_delay_38_3;
  reg                 io_A_Valid_5_delay_39_2;
  reg                 io_A_Valid_5_delay_40_1;
  reg                 io_A_Valid_5_delay_41;
  reg                 io_B_Valid_41_delay_1_4;
  reg                 io_B_Valid_41_delay_2_3;
  reg                 io_B_Valid_41_delay_3_2;
  reg                 io_B_Valid_41_delay_4_1;
  reg                 io_B_Valid_41_delay_5;
  reg                 io_A_Valid_5_delay_1_41;
  reg                 io_A_Valid_5_delay_2_40;
  reg                 io_A_Valid_5_delay_3_39;
  reg                 io_A_Valid_5_delay_4_38;
  reg                 io_A_Valid_5_delay_5_37;
  reg                 io_A_Valid_5_delay_6_36;
  reg                 io_A_Valid_5_delay_7_35;
  reg                 io_A_Valid_5_delay_8_34;
  reg                 io_A_Valid_5_delay_9_33;
  reg                 io_A_Valid_5_delay_10_32;
  reg                 io_A_Valid_5_delay_11_31;
  reg                 io_A_Valid_5_delay_12_30;
  reg                 io_A_Valid_5_delay_13_29;
  reg                 io_A_Valid_5_delay_14_28;
  reg                 io_A_Valid_5_delay_15_27;
  reg                 io_A_Valid_5_delay_16_26;
  reg                 io_A_Valid_5_delay_17_25;
  reg                 io_A_Valid_5_delay_18_24;
  reg                 io_A_Valid_5_delay_19_23;
  reg                 io_A_Valid_5_delay_20_22;
  reg                 io_A_Valid_5_delay_21_21;
  reg                 io_A_Valid_5_delay_22_20;
  reg                 io_A_Valid_5_delay_23_19;
  reg                 io_A_Valid_5_delay_24_18;
  reg                 io_A_Valid_5_delay_25_17;
  reg                 io_A_Valid_5_delay_26_16;
  reg                 io_A_Valid_5_delay_27_15;
  reg                 io_A_Valid_5_delay_28_14;
  reg                 io_A_Valid_5_delay_29_13;
  reg                 io_A_Valid_5_delay_30_12;
  reg                 io_A_Valid_5_delay_31_11;
  reg                 io_A_Valid_5_delay_32_10;
  reg                 io_A_Valid_5_delay_33_9;
  reg                 io_A_Valid_5_delay_34_8;
  reg                 io_A_Valid_5_delay_35_7;
  reg                 io_A_Valid_5_delay_36_6;
  reg                 io_A_Valid_5_delay_37_5;
  reg                 io_A_Valid_5_delay_38_4;
  reg                 io_A_Valid_5_delay_39_3;
  reg                 io_A_Valid_5_delay_40_2;
  reg                 io_A_Valid_5_delay_41_1;
  reg                 io_A_Valid_5_delay_42;
  reg                 io_B_Valid_42_delay_1_4;
  reg                 io_B_Valid_42_delay_2_3;
  reg                 io_B_Valid_42_delay_3_2;
  reg                 io_B_Valid_42_delay_4_1;
  reg                 io_B_Valid_42_delay_5;
  reg                 io_A_Valid_5_delay_1_42;
  reg                 io_A_Valid_5_delay_2_41;
  reg                 io_A_Valid_5_delay_3_40;
  reg                 io_A_Valid_5_delay_4_39;
  reg                 io_A_Valid_5_delay_5_38;
  reg                 io_A_Valid_5_delay_6_37;
  reg                 io_A_Valid_5_delay_7_36;
  reg                 io_A_Valid_5_delay_8_35;
  reg                 io_A_Valid_5_delay_9_34;
  reg                 io_A_Valid_5_delay_10_33;
  reg                 io_A_Valid_5_delay_11_32;
  reg                 io_A_Valid_5_delay_12_31;
  reg                 io_A_Valid_5_delay_13_30;
  reg                 io_A_Valid_5_delay_14_29;
  reg                 io_A_Valid_5_delay_15_28;
  reg                 io_A_Valid_5_delay_16_27;
  reg                 io_A_Valid_5_delay_17_26;
  reg                 io_A_Valid_5_delay_18_25;
  reg                 io_A_Valid_5_delay_19_24;
  reg                 io_A_Valid_5_delay_20_23;
  reg                 io_A_Valid_5_delay_21_22;
  reg                 io_A_Valid_5_delay_22_21;
  reg                 io_A_Valid_5_delay_23_20;
  reg                 io_A_Valid_5_delay_24_19;
  reg                 io_A_Valid_5_delay_25_18;
  reg                 io_A_Valid_5_delay_26_17;
  reg                 io_A_Valid_5_delay_27_16;
  reg                 io_A_Valid_5_delay_28_15;
  reg                 io_A_Valid_5_delay_29_14;
  reg                 io_A_Valid_5_delay_30_13;
  reg                 io_A_Valid_5_delay_31_12;
  reg                 io_A_Valid_5_delay_32_11;
  reg                 io_A_Valid_5_delay_33_10;
  reg                 io_A_Valid_5_delay_34_9;
  reg                 io_A_Valid_5_delay_35_8;
  reg                 io_A_Valid_5_delay_36_7;
  reg                 io_A_Valid_5_delay_37_6;
  reg                 io_A_Valid_5_delay_38_5;
  reg                 io_A_Valid_5_delay_39_4;
  reg                 io_A_Valid_5_delay_40_3;
  reg                 io_A_Valid_5_delay_41_2;
  reg                 io_A_Valid_5_delay_42_1;
  reg                 io_A_Valid_5_delay_43;
  reg                 io_B_Valid_43_delay_1_4;
  reg                 io_B_Valid_43_delay_2_3;
  reg                 io_B_Valid_43_delay_3_2;
  reg                 io_B_Valid_43_delay_4_1;
  reg                 io_B_Valid_43_delay_5;
  reg                 io_A_Valid_5_delay_1_43;
  reg                 io_A_Valid_5_delay_2_42;
  reg                 io_A_Valid_5_delay_3_41;
  reg                 io_A_Valid_5_delay_4_40;
  reg                 io_A_Valid_5_delay_5_39;
  reg                 io_A_Valid_5_delay_6_38;
  reg                 io_A_Valid_5_delay_7_37;
  reg                 io_A_Valid_5_delay_8_36;
  reg                 io_A_Valid_5_delay_9_35;
  reg                 io_A_Valid_5_delay_10_34;
  reg                 io_A_Valid_5_delay_11_33;
  reg                 io_A_Valid_5_delay_12_32;
  reg                 io_A_Valid_5_delay_13_31;
  reg                 io_A_Valid_5_delay_14_30;
  reg                 io_A_Valid_5_delay_15_29;
  reg                 io_A_Valid_5_delay_16_28;
  reg                 io_A_Valid_5_delay_17_27;
  reg                 io_A_Valid_5_delay_18_26;
  reg                 io_A_Valid_5_delay_19_25;
  reg                 io_A_Valid_5_delay_20_24;
  reg                 io_A_Valid_5_delay_21_23;
  reg                 io_A_Valid_5_delay_22_22;
  reg                 io_A_Valid_5_delay_23_21;
  reg                 io_A_Valid_5_delay_24_20;
  reg                 io_A_Valid_5_delay_25_19;
  reg                 io_A_Valid_5_delay_26_18;
  reg                 io_A_Valid_5_delay_27_17;
  reg                 io_A_Valid_5_delay_28_16;
  reg                 io_A_Valid_5_delay_29_15;
  reg                 io_A_Valid_5_delay_30_14;
  reg                 io_A_Valid_5_delay_31_13;
  reg                 io_A_Valid_5_delay_32_12;
  reg                 io_A_Valid_5_delay_33_11;
  reg                 io_A_Valid_5_delay_34_10;
  reg                 io_A_Valid_5_delay_35_9;
  reg                 io_A_Valid_5_delay_36_8;
  reg                 io_A_Valid_5_delay_37_7;
  reg                 io_A_Valid_5_delay_38_6;
  reg                 io_A_Valid_5_delay_39_5;
  reg                 io_A_Valid_5_delay_40_4;
  reg                 io_A_Valid_5_delay_41_3;
  reg                 io_A_Valid_5_delay_42_2;
  reg                 io_A_Valid_5_delay_43_1;
  reg                 io_A_Valid_5_delay_44;
  reg                 io_B_Valid_44_delay_1_4;
  reg                 io_B_Valid_44_delay_2_3;
  reg                 io_B_Valid_44_delay_3_2;
  reg                 io_B_Valid_44_delay_4_1;
  reg                 io_B_Valid_44_delay_5;
  reg                 io_A_Valid_5_delay_1_44;
  reg                 io_A_Valid_5_delay_2_43;
  reg                 io_A_Valid_5_delay_3_42;
  reg                 io_A_Valid_5_delay_4_41;
  reg                 io_A_Valid_5_delay_5_40;
  reg                 io_A_Valid_5_delay_6_39;
  reg                 io_A_Valid_5_delay_7_38;
  reg                 io_A_Valid_5_delay_8_37;
  reg                 io_A_Valid_5_delay_9_36;
  reg                 io_A_Valid_5_delay_10_35;
  reg                 io_A_Valid_5_delay_11_34;
  reg                 io_A_Valid_5_delay_12_33;
  reg                 io_A_Valid_5_delay_13_32;
  reg                 io_A_Valid_5_delay_14_31;
  reg                 io_A_Valid_5_delay_15_30;
  reg                 io_A_Valid_5_delay_16_29;
  reg                 io_A_Valid_5_delay_17_28;
  reg                 io_A_Valid_5_delay_18_27;
  reg                 io_A_Valid_5_delay_19_26;
  reg                 io_A_Valid_5_delay_20_25;
  reg                 io_A_Valid_5_delay_21_24;
  reg                 io_A_Valid_5_delay_22_23;
  reg                 io_A_Valid_5_delay_23_22;
  reg                 io_A_Valid_5_delay_24_21;
  reg                 io_A_Valid_5_delay_25_20;
  reg                 io_A_Valid_5_delay_26_19;
  reg                 io_A_Valid_5_delay_27_18;
  reg                 io_A_Valid_5_delay_28_17;
  reg                 io_A_Valid_5_delay_29_16;
  reg                 io_A_Valid_5_delay_30_15;
  reg                 io_A_Valid_5_delay_31_14;
  reg                 io_A_Valid_5_delay_32_13;
  reg                 io_A_Valid_5_delay_33_12;
  reg                 io_A_Valid_5_delay_34_11;
  reg                 io_A_Valid_5_delay_35_10;
  reg                 io_A_Valid_5_delay_36_9;
  reg                 io_A_Valid_5_delay_37_8;
  reg                 io_A_Valid_5_delay_38_7;
  reg                 io_A_Valid_5_delay_39_6;
  reg                 io_A_Valid_5_delay_40_5;
  reg                 io_A_Valid_5_delay_41_4;
  reg                 io_A_Valid_5_delay_42_3;
  reg                 io_A_Valid_5_delay_43_2;
  reg                 io_A_Valid_5_delay_44_1;
  reg                 io_A_Valid_5_delay_45;
  reg                 io_B_Valid_45_delay_1_4;
  reg                 io_B_Valid_45_delay_2_3;
  reg                 io_B_Valid_45_delay_3_2;
  reg                 io_B_Valid_45_delay_4_1;
  reg                 io_B_Valid_45_delay_5;
  reg                 io_A_Valid_5_delay_1_45;
  reg                 io_A_Valid_5_delay_2_44;
  reg                 io_A_Valid_5_delay_3_43;
  reg                 io_A_Valid_5_delay_4_42;
  reg                 io_A_Valid_5_delay_5_41;
  reg                 io_A_Valid_5_delay_6_40;
  reg                 io_A_Valid_5_delay_7_39;
  reg                 io_A_Valid_5_delay_8_38;
  reg                 io_A_Valid_5_delay_9_37;
  reg                 io_A_Valid_5_delay_10_36;
  reg                 io_A_Valid_5_delay_11_35;
  reg                 io_A_Valid_5_delay_12_34;
  reg                 io_A_Valid_5_delay_13_33;
  reg                 io_A_Valid_5_delay_14_32;
  reg                 io_A_Valid_5_delay_15_31;
  reg                 io_A_Valid_5_delay_16_30;
  reg                 io_A_Valid_5_delay_17_29;
  reg                 io_A_Valid_5_delay_18_28;
  reg                 io_A_Valid_5_delay_19_27;
  reg                 io_A_Valid_5_delay_20_26;
  reg                 io_A_Valid_5_delay_21_25;
  reg                 io_A_Valid_5_delay_22_24;
  reg                 io_A_Valid_5_delay_23_23;
  reg                 io_A_Valid_5_delay_24_22;
  reg                 io_A_Valid_5_delay_25_21;
  reg                 io_A_Valid_5_delay_26_20;
  reg                 io_A_Valid_5_delay_27_19;
  reg                 io_A_Valid_5_delay_28_18;
  reg                 io_A_Valid_5_delay_29_17;
  reg                 io_A_Valid_5_delay_30_16;
  reg                 io_A_Valid_5_delay_31_15;
  reg                 io_A_Valid_5_delay_32_14;
  reg                 io_A_Valid_5_delay_33_13;
  reg                 io_A_Valid_5_delay_34_12;
  reg                 io_A_Valid_5_delay_35_11;
  reg                 io_A_Valid_5_delay_36_10;
  reg                 io_A_Valid_5_delay_37_9;
  reg                 io_A_Valid_5_delay_38_8;
  reg                 io_A_Valid_5_delay_39_7;
  reg                 io_A_Valid_5_delay_40_6;
  reg                 io_A_Valid_5_delay_41_5;
  reg                 io_A_Valid_5_delay_42_4;
  reg                 io_A_Valid_5_delay_43_3;
  reg                 io_A_Valid_5_delay_44_2;
  reg                 io_A_Valid_5_delay_45_1;
  reg                 io_A_Valid_5_delay_46;
  reg                 io_B_Valid_46_delay_1_4;
  reg                 io_B_Valid_46_delay_2_3;
  reg                 io_B_Valid_46_delay_3_2;
  reg                 io_B_Valid_46_delay_4_1;
  reg                 io_B_Valid_46_delay_5;
  reg                 io_A_Valid_5_delay_1_46;
  reg                 io_A_Valid_5_delay_2_45;
  reg                 io_A_Valid_5_delay_3_44;
  reg                 io_A_Valid_5_delay_4_43;
  reg                 io_A_Valid_5_delay_5_42;
  reg                 io_A_Valid_5_delay_6_41;
  reg                 io_A_Valid_5_delay_7_40;
  reg                 io_A_Valid_5_delay_8_39;
  reg                 io_A_Valid_5_delay_9_38;
  reg                 io_A_Valid_5_delay_10_37;
  reg                 io_A_Valid_5_delay_11_36;
  reg                 io_A_Valid_5_delay_12_35;
  reg                 io_A_Valid_5_delay_13_34;
  reg                 io_A_Valid_5_delay_14_33;
  reg                 io_A_Valid_5_delay_15_32;
  reg                 io_A_Valid_5_delay_16_31;
  reg                 io_A_Valid_5_delay_17_30;
  reg                 io_A_Valid_5_delay_18_29;
  reg                 io_A_Valid_5_delay_19_28;
  reg                 io_A_Valid_5_delay_20_27;
  reg                 io_A_Valid_5_delay_21_26;
  reg                 io_A_Valid_5_delay_22_25;
  reg                 io_A_Valid_5_delay_23_24;
  reg                 io_A_Valid_5_delay_24_23;
  reg                 io_A_Valid_5_delay_25_22;
  reg                 io_A_Valid_5_delay_26_21;
  reg                 io_A_Valid_5_delay_27_20;
  reg                 io_A_Valid_5_delay_28_19;
  reg                 io_A_Valid_5_delay_29_18;
  reg                 io_A_Valid_5_delay_30_17;
  reg                 io_A_Valid_5_delay_31_16;
  reg                 io_A_Valid_5_delay_32_15;
  reg                 io_A_Valid_5_delay_33_14;
  reg                 io_A_Valid_5_delay_34_13;
  reg                 io_A_Valid_5_delay_35_12;
  reg                 io_A_Valid_5_delay_36_11;
  reg                 io_A_Valid_5_delay_37_10;
  reg                 io_A_Valid_5_delay_38_9;
  reg                 io_A_Valid_5_delay_39_8;
  reg                 io_A_Valid_5_delay_40_7;
  reg                 io_A_Valid_5_delay_41_6;
  reg                 io_A_Valid_5_delay_42_5;
  reg                 io_A_Valid_5_delay_43_4;
  reg                 io_A_Valid_5_delay_44_3;
  reg                 io_A_Valid_5_delay_45_2;
  reg                 io_A_Valid_5_delay_46_1;
  reg                 io_A_Valid_5_delay_47;
  reg                 io_B_Valid_47_delay_1_4;
  reg                 io_B_Valid_47_delay_2_3;
  reg                 io_B_Valid_47_delay_3_2;
  reg                 io_B_Valid_47_delay_4_1;
  reg                 io_B_Valid_47_delay_5;
  reg                 io_A_Valid_5_delay_1_47;
  reg                 io_A_Valid_5_delay_2_46;
  reg                 io_A_Valid_5_delay_3_45;
  reg                 io_A_Valid_5_delay_4_44;
  reg                 io_A_Valid_5_delay_5_43;
  reg                 io_A_Valid_5_delay_6_42;
  reg                 io_A_Valid_5_delay_7_41;
  reg                 io_A_Valid_5_delay_8_40;
  reg                 io_A_Valid_5_delay_9_39;
  reg                 io_A_Valid_5_delay_10_38;
  reg                 io_A_Valid_5_delay_11_37;
  reg                 io_A_Valid_5_delay_12_36;
  reg                 io_A_Valid_5_delay_13_35;
  reg                 io_A_Valid_5_delay_14_34;
  reg                 io_A_Valid_5_delay_15_33;
  reg                 io_A_Valid_5_delay_16_32;
  reg                 io_A_Valid_5_delay_17_31;
  reg                 io_A_Valid_5_delay_18_30;
  reg                 io_A_Valid_5_delay_19_29;
  reg                 io_A_Valid_5_delay_20_28;
  reg                 io_A_Valid_5_delay_21_27;
  reg                 io_A_Valid_5_delay_22_26;
  reg                 io_A_Valid_5_delay_23_25;
  reg                 io_A_Valid_5_delay_24_24;
  reg                 io_A_Valid_5_delay_25_23;
  reg                 io_A_Valid_5_delay_26_22;
  reg                 io_A_Valid_5_delay_27_21;
  reg                 io_A_Valid_5_delay_28_20;
  reg                 io_A_Valid_5_delay_29_19;
  reg                 io_A_Valid_5_delay_30_18;
  reg                 io_A_Valid_5_delay_31_17;
  reg                 io_A_Valid_5_delay_32_16;
  reg                 io_A_Valid_5_delay_33_15;
  reg                 io_A_Valid_5_delay_34_14;
  reg                 io_A_Valid_5_delay_35_13;
  reg                 io_A_Valid_5_delay_36_12;
  reg                 io_A_Valid_5_delay_37_11;
  reg                 io_A_Valid_5_delay_38_10;
  reg                 io_A_Valid_5_delay_39_9;
  reg                 io_A_Valid_5_delay_40_8;
  reg                 io_A_Valid_5_delay_41_7;
  reg                 io_A_Valid_5_delay_42_6;
  reg                 io_A_Valid_5_delay_43_5;
  reg                 io_A_Valid_5_delay_44_4;
  reg                 io_A_Valid_5_delay_45_3;
  reg                 io_A_Valid_5_delay_46_2;
  reg                 io_A_Valid_5_delay_47_1;
  reg                 io_A_Valid_5_delay_48;
  reg                 io_B_Valid_48_delay_1_4;
  reg                 io_B_Valid_48_delay_2_3;
  reg                 io_B_Valid_48_delay_3_2;
  reg                 io_B_Valid_48_delay_4_1;
  reg                 io_B_Valid_48_delay_5;
  reg                 io_A_Valid_5_delay_1_48;
  reg                 io_A_Valid_5_delay_2_47;
  reg                 io_A_Valid_5_delay_3_46;
  reg                 io_A_Valid_5_delay_4_45;
  reg                 io_A_Valid_5_delay_5_44;
  reg                 io_A_Valid_5_delay_6_43;
  reg                 io_A_Valid_5_delay_7_42;
  reg                 io_A_Valid_5_delay_8_41;
  reg                 io_A_Valid_5_delay_9_40;
  reg                 io_A_Valid_5_delay_10_39;
  reg                 io_A_Valid_5_delay_11_38;
  reg                 io_A_Valid_5_delay_12_37;
  reg                 io_A_Valid_5_delay_13_36;
  reg                 io_A_Valid_5_delay_14_35;
  reg                 io_A_Valid_5_delay_15_34;
  reg                 io_A_Valid_5_delay_16_33;
  reg                 io_A_Valid_5_delay_17_32;
  reg                 io_A_Valid_5_delay_18_31;
  reg                 io_A_Valid_5_delay_19_30;
  reg                 io_A_Valid_5_delay_20_29;
  reg                 io_A_Valid_5_delay_21_28;
  reg                 io_A_Valid_5_delay_22_27;
  reg                 io_A_Valid_5_delay_23_26;
  reg                 io_A_Valid_5_delay_24_25;
  reg                 io_A_Valid_5_delay_25_24;
  reg                 io_A_Valid_5_delay_26_23;
  reg                 io_A_Valid_5_delay_27_22;
  reg                 io_A_Valid_5_delay_28_21;
  reg                 io_A_Valid_5_delay_29_20;
  reg                 io_A_Valid_5_delay_30_19;
  reg                 io_A_Valid_5_delay_31_18;
  reg                 io_A_Valid_5_delay_32_17;
  reg                 io_A_Valid_5_delay_33_16;
  reg                 io_A_Valid_5_delay_34_15;
  reg                 io_A_Valid_5_delay_35_14;
  reg                 io_A_Valid_5_delay_36_13;
  reg                 io_A_Valid_5_delay_37_12;
  reg                 io_A_Valid_5_delay_38_11;
  reg                 io_A_Valid_5_delay_39_10;
  reg                 io_A_Valid_5_delay_40_9;
  reg                 io_A_Valid_5_delay_41_8;
  reg                 io_A_Valid_5_delay_42_7;
  reg                 io_A_Valid_5_delay_43_6;
  reg                 io_A_Valid_5_delay_44_5;
  reg                 io_A_Valid_5_delay_45_4;
  reg                 io_A_Valid_5_delay_46_3;
  reg                 io_A_Valid_5_delay_47_2;
  reg                 io_A_Valid_5_delay_48_1;
  reg                 io_A_Valid_5_delay_49;
  reg                 io_B_Valid_49_delay_1_4;
  reg                 io_B_Valid_49_delay_2_3;
  reg                 io_B_Valid_49_delay_3_2;
  reg                 io_B_Valid_49_delay_4_1;
  reg                 io_B_Valid_49_delay_5;
  reg                 io_A_Valid_5_delay_1_49;
  reg                 io_A_Valid_5_delay_2_48;
  reg                 io_A_Valid_5_delay_3_47;
  reg                 io_A_Valid_5_delay_4_46;
  reg                 io_A_Valid_5_delay_5_45;
  reg                 io_A_Valid_5_delay_6_44;
  reg                 io_A_Valid_5_delay_7_43;
  reg                 io_A_Valid_5_delay_8_42;
  reg                 io_A_Valid_5_delay_9_41;
  reg                 io_A_Valid_5_delay_10_40;
  reg                 io_A_Valid_5_delay_11_39;
  reg                 io_A_Valid_5_delay_12_38;
  reg                 io_A_Valid_5_delay_13_37;
  reg                 io_A_Valid_5_delay_14_36;
  reg                 io_A_Valid_5_delay_15_35;
  reg                 io_A_Valid_5_delay_16_34;
  reg                 io_A_Valid_5_delay_17_33;
  reg                 io_A_Valid_5_delay_18_32;
  reg                 io_A_Valid_5_delay_19_31;
  reg                 io_A_Valid_5_delay_20_30;
  reg                 io_A_Valid_5_delay_21_29;
  reg                 io_A_Valid_5_delay_22_28;
  reg                 io_A_Valid_5_delay_23_27;
  reg                 io_A_Valid_5_delay_24_26;
  reg                 io_A_Valid_5_delay_25_25;
  reg                 io_A_Valid_5_delay_26_24;
  reg                 io_A_Valid_5_delay_27_23;
  reg                 io_A_Valid_5_delay_28_22;
  reg                 io_A_Valid_5_delay_29_21;
  reg                 io_A_Valid_5_delay_30_20;
  reg                 io_A_Valid_5_delay_31_19;
  reg                 io_A_Valid_5_delay_32_18;
  reg                 io_A_Valid_5_delay_33_17;
  reg                 io_A_Valid_5_delay_34_16;
  reg                 io_A_Valid_5_delay_35_15;
  reg                 io_A_Valid_5_delay_36_14;
  reg                 io_A_Valid_5_delay_37_13;
  reg                 io_A_Valid_5_delay_38_12;
  reg                 io_A_Valid_5_delay_39_11;
  reg                 io_A_Valid_5_delay_40_10;
  reg                 io_A_Valid_5_delay_41_9;
  reg                 io_A_Valid_5_delay_42_8;
  reg                 io_A_Valid_5_delay_43_7;
  reg                 io_A_Valid_5_delay_44_6;
  reg                 io_A_Valid_5_delay_45_5;
  reg                 io_A_Valid_5_delay_46_4;
  reg                 io_A_Valid_5_delay_47_3;
  reg                 io_A_Valid_5_delay_48_2;
  reg                 io_A_Valid_5_delay_49_1;
  reg                 io_A_Valid_5_delay_50;
  reg                 io_B_Valid_50_delay_1_4;
  reg                 io_B_Valid_50_delay_2_3;
  reg                 io_B_Valid_50_delay_3_2;
  reg                 io_B_Valid_50_delay_4_1;
  reg                 io_B_Valid_50_delay_5;
  reg                 io_A_Valid_5_delay_1_50;
  reg                 io_A_Valid_5_delay_2_49;
  reg                 io_A_Valid_5_delay_3_48;
  reg                 io_A_Valid_5_delay_4_47;
  reg                 io_A_Valid_5_delay_5_46;
  reg                 io_A_Valid_5_delay_6_45;
  reg                 io_A_Valid_5_delay_7_44;
  reg                 io_A_Valid_5_delay_8_43;
  reg                 io_A_Valid_5_delay_9_42;
  reg                 io_A_Valid_5_delay_10_41;
  reg                 io_A_Valid_5_delay_11_40;
  reg                 io_A_Valid_5_delay_12_39;
  reg                 io_A_Valid_5_delay_13_38;
  reg                 io_A_Valid_5_delay_14_37;
  reg                 io_A_Valid_5_delay_15_36;
  reg                 io_A_Valid_5_delay_16_35;
  reg                 io_A_Valid_5_delay_17_34;
  reg                 io_A_Valid_5_delay_18_33;
  reg                 io_A_Valid_5_delay_19_32;
  reg                 io_A_Valid_5_delay_20_31;
  reg                 io_A_Valid_5_delay_21_30;
  reg                 io_A_Valid_5_delay_22_29;
  reg                 io_A_Valid_5_delay_23_28;
  reg                 io_A_Valid_5_delay_24_27;
  reg                 io_A_Valid_5_delay_25_26;
  reg                 io_A_Valid_5_delay_26_25;
  reg                 io_A_Valid_5_delay_27_24;
  reg                 io_A_Valid_5_delay_28_23;
  reg                 io_A_Valid_5_delay_29_22;
  reg                 io_A_Valid_5_delay_30_21;
  reg                 io_A_Valid_5_delay_31_20;
  reg                 io_A_Valid_5_delay_32_19;
  reg                 io_A_Valid_5_delay_33_18;
  reg                 io_A_Valid_5_delay_34_17;
  reg                 io_A_Valid_5_delay_35_16;
  reg                 io_A_Valid_5_delay_36_15;
  reg                 io_A_Valid_5_delay_37_14;
  reg                 io_A_Valid_5_delay_38_13;
  reg                 io_A_Valid_5_delay_39_12;
  reg                 io_A_Valid_5_delay_40_11;
  reg                 io_A_Valid_5_delay_41_10;
  reg                 io_A_Valid_5_delay_42_9;
  reg                 io_A_Valid_5_delay_43_8;
  reg                 io_A_Valid_5_delay_44_7;
  reg                 io_A_Valid_5_delay_45_6;
  reg                 io_A_Valid_5_delay_46_5;
  reg                 io_A_Valid_5_delay_47_4;
  reg                 io_A_Valid_5_delay_48_3;
  reg                 io_A_Valid_5_delay_49_2;
  reg                 io_A_Valid_5_delay_50_1;
  reg                 io_A_Valid_5_delay_51;
  reg                 io_B_Valid_51_delay_1_4;
  reg                 io_B_Valid_51_delay_2_3;
  reg                 io_B_Valid_51_delay_3_2;
  reg                 io_B_Valid_51_delay_4_1;
  reg                 io_B_Valid_51_delay_5;
  reg                 io_A_Valid_5_delay_1_51;
  reg                 io_A_Valid_5_delay_2_50;
  reg                 io_A_Valid_5_delay_3_49;
  reg                 io_A_Valid_5_delay_4_48;
  reg                 io_A_Valid_5_delay_5_47;
  reg                 io_A_Valid_5_delay_6_46;
  reg                 io_A_Valid_5_delay_7_45;
  reg                 io_A_Valid_5_delay_8_44;
  reg                 io_A_Valid_5_delay_9_43;
  reg                 io_A_Valid_5_delay_10_42;
  reg                 io_A_Valid_5_delay_11_41;
  reg                 io_A_Valid_5_delay_12_40;
  reg                 io_A_Valid_5_delay_13_39;
  reg                 io_A_Valid_5_delay_14_38;
  reg                 io_A_Valid_5_delay_15_37;
  reg                 io_A_Valid_5_delay_16_36;
  reg                 io_A_Valid_5_delay_17_35;
  reg                 io_A_Valid_5_delay_18_34;
  reg                 io_A_Valid_5_delay_19_33;
  reg                 io_A_Valid_5_delay_20_32;
  reg                 io_A_Valid_5_delay_21_31;
  reg                 io_A_Valid_5_delay_22_30;
  reg                 io_A_Valid_5_delay_23_29;
  reg                 io_A_Valid_5_delay_24_28;
  reg                 io_A_Valid_5_delay_25_27;
  reg                 io_A_Valid_5_delay_26_26;
  reg                 io_A_Valid_5_delay_27_25;
  reg                 io_A_Valid_5_delay_28_24;
  reg                 io_A_Valid_5_delay_29_23;
  reg                 io_A_Valid_5_delay_30_22;
  reg                 io_A_Valid_5_delay_31_21;
  reg                 io_A_Valid_5_delay_32_20;
  reg                 io_A_Valid_5_delay_33_19;
  reg                 io_A_Valid_5_delay_34_18;
  reg                 io_A_Valid_5_delay_35_17;
  reg                 io_A_Valid_5_delay_36_16;
  reg                 io_A_Valid_5_delay_37_15;
  reg                 io_A_Valid_5_delay_38_14;
  reg                 io_A_Valid_5_delay_39_13;
  reg                 io_A_Valid_5_delay_40_12;
  reg                 io_A_Valid_5_delay_41_11;
  reg                 io_A_Valid_5_delay_42_10;
  reg                 io_A_Valid_5_delay_43_9;
  reg                 io_A_Valid_5_delay_44_8;
  reg                 io_A_Valid_5_delay_45_7;
  reg                 io_A_Valid_5_delay_46_6;
  reg                 io_A_Valid_5_delay_47_5;
  reg                 io_A_Valid_5_delay_48_4;
  reg                 io_A_Valid_5_delay_49_3;
  reg                 io_A_Valid_5_delay_50_2;
  reg                 io_A_Valid_5_delay_51_1;
  reg                 io_A_Valid_5_delay_52;
  reg                 io_B_Valid_52_delay_1_4;
  reg                 io_B_Valid_52_delay_2_3;
  reg                 io_B_Valid_52_delay_3_2;
  reg                 io_B_Valid_52_delay_4_1;
  reg                 io_B_Valid_52_delay_5;
  reg                 io_A_Valid_5_delay_1_52;
  reg                 io_A_Valid_5_delay_2_51;
  reg                 io_A_Valid_5_delay_3_50;
  reg                 io_A_Valid_5_delay_4_49;
  reg                 io_A_Valid_5_delay_5_48;
  reg                 io_A_Valid_5_delay_6_47;
  reg                 io_A_Valid_5_delay_7_46;
  reg                 io_A_Valid_5_delay_8_45;
  reg                 io_A_Valid_5_delay_9_44;
  reg                 io_A_Valid_5_delay_10_43;
  reg                 io_A_Valid_5_delay_11_42;
  reg                 io_A_Valid_5_delay_12_41;
  reg                 io_A_Valid_5_delay_13_40;
  reg                 io_A_Valid_5_delay_14_39;
  reg                 io_A_Valid_5_delay_15_38;
  reg                 io_A_Valid_5_delay_16_37;
  reg                 io_A_Valid_5_delay_17_36;
  reg                 io_A_Valid_5_delay_18_35;
  reg                 io_A_Valid_5_delay_19_34;
  reg                 io_A_Valid_5_delay_20_33;
  reg                 io_A_Valid_5_delay_21_32;
  reg                 io_A_Valid_5_delay_22_31;
  reg                 io_A_Valid_5_delay_23_30;
  reg                 io_A_Valid_5_delay_24_29;
  reg                 io_A_Valid_5_delay_25_28;
  reg                 io_A_Valid_5_delay_26_27;
  reg                 io_A_Valid_5_delay_27_26;
  reg                 io_A_Valid_5_delay_28_25;
  reg                 io_A_Valid_5_delay_29_24;
  reg                 io_A_Valid_5_delay_30_23;
  reg                 io_A_Valid_5_delay_31_22;
  reg                 io_A_Valid_5_delay_32_21;
  reg                 io_A_Valid_5_delay_33_20;
  reg                 io_A_Valid_5_delay_34_19;
  reg                 io_A_Valid_5_delay_35_18;
  reg                 io_A_Valid_5_delay_36_17;
  reg                 io_A_Valid_5_delay_37_16;
  reg                 io_A_Valid_5_delay_38_15;
  reg                 io_A_Valid_5_delay_39_14;
  reg                 io_A_Valid_5_delay_40_13;
  reg                 io_A_Valid_5_delay_41_12;
  reg                 io_A_Valid_5_delay_42_11;
  reg                 io_A_Valid_5_delay_43_10;
  reg                 io_A_Valid_5_delay_44_9;
  reg                 io_A_Valid_5_delay_45_8;
  reg                 io_A_Valid_5_delay_46_7;
  reg                 io_A_Valid_5_delay_47_6;
  reg                 io_A_Valid_5_delay_48_5;
  reg                 io_A_Valid_5_delay_49_4;
  reg                 io_A_Valid_5_delay_50_3;
  reg                 io_A_Valid_5_delay_51_2;
  reg                 io_A_Valid_5_delay_52_1;
  reg                 io_A_Valid_5_delay_53;
  reg                 io_B_Valid_53_delay_1_4;
  reg                 io_B_Valid_53_delay_2_3;
  reg                 io_B_Valid_53_delay_3_2;
  reg                 io_B_Valid_53_delay_4_1;
  reg                 io_B_Valid_53_delay_5;
  reg                 io_A_Valid_5_delay_1_53;
  reg                 io_A_Valid_5_delay_2_52;
  reg                 io_A_Valid_5_delay_3_51;
  reg                 io_A_Valid_5_delay_4_50;
  reg                 io_A_Valid_5_delay_5_49;
  reg                 io_A_Valid_5_delay_6_48;
  reg                 io_A_Valid_5_delay_7_47;
  reg                 io_A_Valid_5_delay_8_46;
  reg                 io_A_Valid_5_delay_9_45;
  reg                 io_A_Valid_5_delay_10_44;
  reg                 io_A_Valid_5_delay_11_43;
  reg                 io_A_Valid_5_delay_12_42;
  reg                 io_A_Valid_5_delay_13_41;
  reg                 io_A_Valid_5_delay_14_40;
  reg                 io_A_Valid_5_delay_15_39;
  reg                 io_A_Valid_5_delay_16_38;
  reg                 io_A_Valid_5_delay_17_37;
  reg                 io_A_Valid_5_delay_18_36;
  reg                 io_A_Valid_5_delay_19_35;
  reg                 io_A_Valid_5_delay_20_34;
  reg                 io_A_Valid_5_delay_21_33;
  reg                 io_A_Valid_5_delay_22_32;
  reg                 io_A_Valid_5_delay_23_31;
  reg                 io_A_Valid_5_delay_24_30;
  reg                 io_A_Valid_5_delay_25_29;
  reg                 io_A_Valid_5_delay_26_28;
  reg                 io_A_Valid_5_delay_27_27;
  reg                 io_A_Valid_5_delay_28_26;
  reg                 io_A_Valid_5_delay_29_25;
  reg                 io_A_Valid_5_delay_30_24;
  reg                 io_A_Valid_5_delay_31_23;
  reg                 io_A_Valid_5_delay_32_22;
  reg                 io_A_Valid_5_delay_33_21;
  reg                 io_A_Valid_5_delay_34_20;
  reg                 io_A_Valid_5_delay_35_19;
  reg                 io_A_Valid_5_delay_36_18;
  reg                 io_A_Valid_5_delay_37_17;
  reg                 io_A_Valid_5_delay_38_16;
  reg                 io_A_Valid_5_delay_39_15;
  reg                 io_A_Valid_5_delay_40_14;
  reg                 io_A_Valid_5_delay_41_13;
  reg                 io_A_Valid_5_delay_42_12;
  reg                 io_A_Valid_5_delay_43_11;
  reg                 io_A_Valid_5_delay_44_10;
  reg                 io_A_Valid_5_delay_45_9;
  reg                 io_A_Valid_5_delay_46_8;
  reg                 io_A_Valid_5_delay_47_7;
  reg                 io_A_Valid_5_delay_48_6;
  reg                 io_A_Valid_5_delay_49_5;
  reg                 io_A_Valid_5_delay_50_4;
  reg                 io_A_Valid_5_delay_51_3;
  reg                 io_A_Valid_5_delay_52_2;
  reg                 io_A_Valid_5_delay_53_1;
  reg                 io_A_Valid_5_delay_54;
  reg                 io_B_Valid_54_delay_1_4;
  reg                 io_B_Valid_54_delay_2_3;
  reg                 io_B_Valid_54_delay_3_2;
  reg                 io_B_Valid_54_delay_4_1;
  reg                 io_B_Valid_54_delay_5;
  reg                 io_A_Valid_5_delay_1_54;
  reg                 io_A_Valid_5_delay_2_53;
  reg                 io_A_Valid_5_delay_3_52;
  reg                 io_A_Valid_5_delay_4_51;
  reg                 io_A_Valid_5_delay_5_50;
  reg                 io_A_Valid_5_delay_6_49;
  reg                 io_A_Valid_5_delay_7_48;
  reg                 io_A_Valid_5_delay_8_47;
  reg                 io_A_Valid_5_delay_9_46;
  reg                 io_A_Valid_5_delay_10_45;
  reg                 io_A_Valid_5_delay_11_44;
  reg                 io_A_Valid_5_delay_12_43;
  reg                 io_A_Valid_5_delay_13_42;
  reg                 io_A_Valid_5_delay_14_41;
  reg                 io_A_Valid_5_delay_15_40;
  reg                 io_A_Valid_5_delay_16_39;
  reg                 io_A_Valid_5_delay_17_38;
  reg                 io_A_Valid_5_delay_18_37;
  reg                 io_A_Valid_5_delay_19_36;
  reg                 io_A_Valid_5_delay_20_35;
  reg                 io_A_Valid_5_delay_21_34;
  reg                 io_A_Valid_5_delay_22_33;
  reg                 io_A_Valid_5_delay_23_32;
  reg                 io_A_Valid_5_delay_24_31;
  reg                 io_A_Valid_5_delay_25_30;
  reg                 io_A_Valid_5_delay_26_29;
  reg                 io_A_Valid_5_delay_27_28;
  reg                 io_A_Valid_5_delay_28_27;
  reg                 io_A_Valid_5_delay_29_26;
  reg                 io_A_Valid_5_delay_30_25;
  reg                 io_A_Valid_5_delay_31_24;
  reg                 io_A_Valid_5_delay_32_23;
  reg                 io_A_Valid_5_delay_33_22;
  reg                 io_A_Valid_5_delay_34_21;
  reg                 io_A_Valid_5_delay_35_20;
  reg                 io_A_Valid_5_delay_36_19;
  reg                 io_A_Valid_5_delay_37_18;
  reg                 io_A_Valid_5_delay_38_17;
  reg                 io_A_Valid_5_delay_39_16;
  reg                 io_A_Valid_5_delay_40_15;
  reg                 io_A_Valid_5_delay_41_14;
  reg                 io_A_Valid_5_delay_42_13;
  reg                 io_A_Valid_5_delay_43_12;
  reg                 io_A_Valid_5_delay_44_11;
  reg                 io_A_Valid_5_delay_45_10;
  reg                 io_A_Valid_5_delay_46_9;
  reg                 io_A_Valid_5_delay_47_8;
  reg                 io_A_Valid_5_delay_48_7;
  reg                 io_A_Valid_5_delay_49_6;
  reg                 io_A_Valid_5_delay_50_5;
  reg                 io_A_Valid_5_delay_51_4;
  reg                 io_A_Valid_5_delay_52_3;
  reg                 io_A_Valid_5_delay_53_2;
  reg                 io_A_Valid_5_delay_54_1;
  reg                 io_A_Valid_5_delay_55;
  reg                 io_B_Valid_55_delay_1_4;
  reg                 io_B_Valid_55_delay_2_3;
  reg                 io_B_Valid_55_delay_3_2;
  reg                 io_B_Valid_55_delay_4_1;
  reg                 io_B_Valid_55_delay_5;
  reg                 io_A_Valid_5_delay_1_55;
  reg                 io_A_Valid_5_delay_2_54;
  reg                 io_A_Valid_5_delay_3_53;
  reg                 io_A_Valid_5_delay_4_52;
  reg                 io_A_Valid_5_delay_5_51;
  reg                 io_A_Valid_5_delay_6_50;
  reg                 io_A_Valid_5_delay_7_49;
  reg                 io_A_Valid_5_delay_8_48;
  reg                 io_A_Valid_5_delay_9_47;
  reg                 io_A_Valid_5_delay_10_46;
  reg                 io_A_Valid_5_delay_11_45;
  reg                 io_A_Valid_5_delay_12_44;
  reg                 io_A_Valid_5_delay_13_43;
  reg                 io_A_Valid_5_delay_14_42;
  reg                 io_A_Valid_5_delay_15_41;
  reg                 io_A_Valid_5_delay_16_40;
  reg                 io_A_Valid_5_delay_17_39;
  reg                 io_A_Valid_5_delay_18_38;
  reg                 io_A_Valid_5_delay_19_37;
  reg                 io_A_Valid_5_delay_20_36;
  reg                 io_A_Valid_5_delay_21_35;
  reg                 io_A_Valid_5_delay_22_34;
  reg                 io_A_Valid_5_delay_23_33;
  reg                 io_A_Valid_5_delay_24_32;
  reg                 io_A_Valid_5_delay_25_31;
  reg                 io_A_Valid_5_delay_26_30;
  reg                 io_A_Valid_5_delay_27_29;
  reg                 io_A_Valid_5_delay_28_28;
  reg                 io_A_Valid_5_delay_29_27;
  reg                 io_A_Valid_5_delay_30_26;
  reg                 io_A_Valid_5_delay_31_25;
  reg                 io_A_Valid_5_delay_32_24;
  reg                 io_A_Valid_5_delay_33_23;
  reg                 io_A_Valid_5_delay_34_22;
  reg                 io_A_Valid_5_delay_35_21;
  reg                 io_A_Valid_5_delay_36_20;
  reg                 io_A_Valid_5_delay_37_19;
  reg                 io_A_Valid_5_delay_38_18;
  reg                 io_A_Valid_5_delay_39_17;
  reg                 io_A_Valid_5_delay_40_16;
  reg                 io_A_Valid_5_delay_41_15;
  reg                 io_A_Valid_5_delay_42_14;
  reg                 io_A_Valid_5_delay_43_13;
  reg                 io_A_Valid_5_delay_44_12;
  reg                 io_A_Valid_5_delay_45_11;
  reg                 io_A_Valid_5_delay_46_10;
  reg                 io_A_Valid_5_delay_47_9;
  reg                 io_A_Valid_5_delay_48_8;
  reg                 io_A_Valid_5_delay_49_7;
  reg                 io_A_Valid_5_delay_50_6;
  reg                 io_A_Valid_5_delay_51_5;
  reg                 io_A_Valid_5_delay_52_4;
  reg                 io_A_Valid_5_delay_53_3;
  reg                 io_A_Valid_5_delay_54_2;
  reg                 io_A_Valid_5_delay_55_1;
  reg                 io_A_Valid_5_delay_56;
  reg                 io_B_Valid_56_delay_1_4;
  reg                 io_B_Valid_56_delay_2_3;
  reg                 io_B_Valid_56_delay_3_2;
  reg                 io_B_Valid_56_delay_4_1;
  reg                 io_B_Valid_56_delay_5;
  reg                 io_A_Valid_5_delay_1_56;
  reg                 io_A_Valid_5_delay_2_55;
  reg                 io_A_Valid_5_delay_3_54;
  reg                 io_A_Valid_5_delay_4_53;
  reg                 io_A_Valid_5_delay_5_52;
  reg                 io_A_Valid_5_delay_6_51;
  reg                 io_A_Valid_5_delay_7_50;
  reg                 io_A_Valid_5_delay_8_49;
  reg                 io_A_Valid_5_delay_9_48;
  reg                 io_A_Valid_5_delay_10_47;
  reg                 io_A_Valid_5_delay_11_46;
  reg                 io_A_Valid_5_delay_12_45;
  reg                 io_A_Valid_5_delay_13_44;
  reg                 io_A_Valid_5_delay_14_43;
  reg                 io_A_Valid_5_delay_15_42;
  reg                 io_A_Valid_5_delay_16_41;
  reg                 io_A_Valid_5_delay_17_40;
  reg                 io_A_Valid_5_delay_18_39;
  reg                 io_A_Valid_5_delay_19_38;
  reg                 io_A_Valid_5_delay_20_37;
  reg                 io_A_Valid_5_delay_21_36;
  reg                 io_A_Valid_5_delay_22_35;
  reg                 io_A_Valid_5_delay_23_34;
  reg                 io_A_Valid_5_delay_24_33;
  reg                 io_A_Valid_5_delay_25_32;
  reg                 io_A_Valid_5_delay_26_31;
  reg                 io_A_Valid_5_delay_27_30;
  reg                 io_A_Valid_5_delay_28_29;
  reg                 io_A_Valid_5_delay_29_28;
  reg                 io_A_Valid_5_delay_30_27;
  reg                 io_A_Valid_5_delay_31_26;
  reg                 io_A_Valid_5_delay_32_25;
  reg                 io_A_Valid_5_delay_33_24;
  reg                 io_A_Valid_5_delay_34_23;
  reg                 io_A_Valid_5_delay_35_22;
  reg                 io_A_Valid_5_delay_36_21;
  reg                 io_A_Valid_5_delay_37_20;
  reg                 io_A_Valid_5_delay_38_19;
  reg                 io_A_Valid_5_delay_39_18;
  reg                 io_A_Valid_5_delay_40_17;
  reg                 io_A_Valid_5_delay_41_16;
  reg                 io_A_Valid_5_delay_42_15;
  reg                 io_A_Valid_5_delay_43_14;
  reg                 io_A_Valid_5_delay_44_13;
  reg                 io_A_Valid_5_delay_45_12;
  reg                 io_A_Valid_5_delay_46_11;
  reg                 io_A_Valid_5_delay_47_10;
  reg                 io_A_Valid_5_delay_48_9;
  reg                 io_A_Valid_5_delay_49_8;
  reg                 io_A_Valid_5_delay_50_7;
  reg                 io_A_Valid_5_delay_51_6;
  reg                 io_A_Valid_5_delay_52_5;
  reg                 io_A_Valid_5_delay_53_4;
  reg                 io_A_Valid_5_delay_54_3;
  reg                 io_A_Valid_5_delay_55_2;
  reg                 io_A_Valid_5_delay_56_1;
  reg                 io_A_Valid_5_delay_57;
  reg                 io_B_Valid_57_delay_1_4;
  reg                 io_B_Valid_57_delay_2_3;
  reg                 io_B_Valid_57_delay_3_2;
  reg                 io_B_Valid_57_delay_4_1;
  reg                 io_B_Valid_57_delay_5;
  reg                 io_A_Valid_5_delay_1_57;
  reg                 io_A_Valid_5_delay_2_56;
  reg                 io_A_Valid_5_delay_3_55;
  reg                 io_A_Valid_5_delay_4_54;
  reg                 io_A_Valid_5_delay_5_53;
  reg                 io_A_Valid_5_delay_6_52;
  reg                 io_A_Valid_5_delay_7_51;
  reg                 io_A_Valid_5_delay_8_50;
  reg                 io_A_Valid_5_delay_9_49;
  reg                 io_A_Valid_5_delay_10_48;
  reg                 io_A_Valid_5_delay_11_47;
  reg                 io_A_Valid_5_delay_12_46;
  reg                 io_A_Valid_5_delay_13_45;
  reg                 io_A_Valid_5_delay_14_44;
  reg                 io_A_Valid_5_delay_15_43;
  reg                 io_A_Valid_5_delay_16_42;
  reg                 io_A_Valid_5_delay_17_41;
  reg                 io_A_Valid_5_delay_18_40;
  reg                 io_A_Valid_5_delay_19_39;
  reg                 io_A_Valid_5_delay_20_38;
  reg                 io_A_Valid_5_delay_21_37;
  reg                 io_A_Valid_5_delay_22_36;
  reg                 io_A_Valid_5_delay_23_35;
  reg                 io_A_Valid_5_delay_24_34;
  reg                 io_A_Valid_5_delay_25_33;
  reg                 io_A_Valid_5_delay_26_32;
  reg                 io_A_Valid_5_delay_27_31;
  reg                 io_A_Valid_5_delay_28_30;
  reg                 io_A_Valid_5_delay_29_29;
  reg                 io_A_Valid_5_delay_30_28;
  reg                 io_A_Valid_5_delay_31_27;
  reg                 io_A_Valid_5_delay_32_26;
  reg                 io_A_Valid_5_delay_33_25;
  reg                 io_A_Valid_5_delay_34_24;
  reg                 io_A_Valid_5_delay_35_23;
  reg                 io_A_Valid_5_delay_36_22;
  reg                 io_A_Valid_5_delay_37_21;
  reg                 io_A_Valid_5_delay_38_20;
  reg                 io_A_Valid_5_delay_39_19;
  reg                 io_A_Valid_5_delay_40_18;
  reg                 io_A_Valid_5_delay_41_17;
  reg                 io_A_Valid_5_delay_42_16;
  reg                 io_A_Valid_5_delay_43_15;
  reg                 io_A_Valid_5_delay_44_14;
  reg                 io_A_Valid_5_delay_45_13;
  reg                 io_A_Valid_5_delay_46_12;
  reg                 io_A_Valid_5_delay_47_11;
  reg                 io_A_Valid_5_delay_48_10;
  reg                 io_A_Valid_5_delay_49_9;
  reg                 io_A_Valid_5_delay_50_8;
  reg                 io_A_Valid_5_delay_51_7;
  reg                 io_A_Valid_5_delay_52_6;
  reg                 io_A_Valid_5_delay_53_5;
  reg                 io_A_Valid_5_delay_54_4;
  reg                 io_A_Valid_5_delay_55_3;
  reg                 io_A_Valid_5_delay_56_2;
  reg                 io_A_Valid_5_delay_57_1;
  reg                 io_A_Valid_5_delay_58;
  reg                 io_B_Valid_58_delay_1_4;
  reg                 io_B_Valid_58_delay_2_3;
  reg                 io_B_Valid_58_delay_3_2;
  reg                 io_B_Valid_58_delay_4_1;
  reg                 io_B_Valid_58_delay_5;
  reg                 io_A_Valid_5_delay_1_58;
  reg                 io_A_Valid_5_delay_2_57;
  reg                 io_A_Valid_5_delay_3_56;
  reg                 io_A_Valid_5_delay_4_55;
  reg                 io_A_Valid_5_delay_5_54;
  reg                 io_A_Valid_5_delay_6_53;
  reg                 io_A_Valid_5_delay_7_52;
  reg                 io_A_Valid_5_delay_8_51;
  reg                 io_A_Valid_5_delay_9_50;
  reg                 io_A_Valid_5_delay_10_49;
  reg                 io_A_Valid_5_delay_11_48;
  reg                 io_A_Valid_5_delay_12_47;
  reg                 io_A_Valid_5_delay_13_46;
  reg                 io_A_Valid_5_delay_14_45;
  reg                 io_A_Valid_5_delay_15_44;
  reg                 io_A_Valid_5_delay_16_43;
  reg                 io_A_Valid_5_delay_17_42;
  reg                 io_A_Valid_5_delay_18_41;
  reg                 io_A_Valid_5_delay_19_40;
  reg                 io_A_Valid_5_delay_20_39;
  reg                 io_A_Valid_5_delay_21_38;
  reg                 io_A_Valid_5_delay_22_37;
  reg                 io_A_Valid_5_delay_23_36;
  reg                 io_A_Valid_5_delay_24_35;
  reg                 io_A_Valid_5_delay_25_34;
  reg                 io_A_Valid_5_delay_26_33;
  reg                 io_A_Valid_5_delay_27_32;
  reg                 io_A_Valid_5_delay_28_31;
  reg                 io_A_Valid_5_delay_29_30;
  reg                 io_A_Valid_5_delay_30_29;
  reg                 io_A_Valid_5_delay_31_28;
  reg                 io_A_Valid_5_delay_32_27;
  reg                 io_A_Valid_5_delay_33_26;
  reg                 io_A_Valid_5_delay_34_25;
  reg                 io_A_Valid_5_delay_35_24;
  reg                 io_A_Valid_5_delay_36_23;
  reg                 io_A_Valid_5_delay_37_22;
  reg                 io_A_Valid_5_delay_38_21;
  reg                 io_A_Valid_5_delay_39_20;
  reg                 io_A_Valid_5_delay_40_19;
  reg                 io_A_Valid_5_delay_41_18;
  reg                 io_A_Valid_5_delay_42_17;
  reg                 io_A_Valid_5_delay_43_16;
  reg                 io_A_Valid_5_delay_44_15;
  reg                 io_A_Valid_5_delay_45_14;
  reg                 io_A_Valid_5_delay_46_13;
  reg                 io_A_Valid_5_delay_47_12;
  reg                 io_A_Valid_5_delay_48_11;
  reg                 io_A_Valid_5_delay_49_10;
  reg                 io_A_Valid_5_delay_50_9;
  reg                 io_A_Valid_5_delay_51_8;
  reg                 io_A_Valid_5_delay_52_7;
  reg                 io_A_Valid_5_delay_53_6;
  reg                 io_A_Valid_5_delay_54_5;
  reg                 io_A_Valid_5_delay_55_4;
  reg                 io_A_Valid_5_delay_56_3;
  reg                 io_A_Valid_5_delay_57_2;
  reg                 io_A_Valid_5_delay_58_1;
  reg                 io_A_Valid_5_delay_59;
  reg                 io_B_Valid_59_delay_1_4;
  reg                 io_B_Valid_59_delay_2_3;
  reg                 io_B_Valid_59_delay_3_2;
  reg                 io_B_Valid_59_delay_4_1;
  reg                 io_B_Valid_59_delay_5;
  reg                 io_A_Valid_5_delay_1_59;
  reg                 io_A_Valid_5_delay_2_58;
  reg                 io_A_Valid_5_delay_3_57;
  reg                 io_A_Valid_5_delay_4_56;
  reg                 io_A_Valid_5_delay_5_55;
  reg                 io_A_Valid_5_delay_6_54;
  reg                 io_A_Valid_5_delay_7_53;
  reg                 io_A_Valid_5_delay_8_52;
  reg                 io_A_Valid_5_delay_9_51;
  reg                 io_A_Valid_5_delay_10_50;
  reg                 io_A_Valid_5_delay_11_49;
  reg                 io_A_Valid_5_delay_12_48;
  reg                 io_A_Valid_5_delay_13_47;
  reg                 io_A_Valid_5_delay_14_46;
  reg                 io_A_Valid_5_delay_15_45;
  reg                 io_A_Valid_5_delay_16_44;
  reg                 io_A_Valid_5_delay_17_43;
  reg                 io_A_Valid_5_delay_18_42;
  reg                 io_A_Valid_5_delay_19_41;
  reg                 io_A_Valid_5_delay_20_40;
  reg                 io_A_Valid_5_delay_21_39;
  reg                 io_A_Valid_5_delay_22_38;
  reg                 io_A_Valid_5_delay_23_37;
  reg                 io_A_Valid_5_delay_24_36;
  reg                 io_A_Valid_5_delay_25_35;
  reg                 io_A_Valid_5_delay_26_34;
  reg                 io_A_Valid_5_delay_27_33;
  reg                 io_A_Valid_5_delay_28_32;
  reg                 io_A_Valid_5_delay_29_31;
  reg                 io_A_Valid_5_delay_30_30;
  reg                 io_A_Valid_5_delay_31_29;
  reg                 io_A_Valid_5_delay_32_28;
  reg                 io_A_Valid_5_delay_33_27;
  reg                 io_A_Valid_5_delay_34_26;
  reg                 io_A_Valid_5_delay_35_25;
  reg                 io_A_Valid_5_delay_36_24;
  reg                 io_A_Valid_5_delay_37_23;
  reg                 io_A_Valid_5_delay_38_22;
  reg                 io_A_Valid_5_delay_39_21;
  reg                 io_A_Valid_5_delay_40_20;
  reg                 io_A_Valid_5_delay_41_19;
  reg                 io_A_Valid_5_delay_42_18;
  reg                 io_A_Valid_5_delay_43_17;
  reg                 io_A_Valid_5_delay_44_16;
  reg                 io_A_Valid_5_delay_45_15;
  reg                 io_A_Valid_5_delay_46_14;
  reg                 io_A_Valid_5_delay_47_13;
  reg                 io_A_Valid_5_delay_48_12;
  reg                 io_A_Valid_5_delay_49_11;
  reg                 io_A_Valid_5_delay_50_10;
  reg                 io_A_Valid_5_delay_51_9;
  reg                 io_A_Valid_5_delay_52_8;
  reg                 io_A_Valid_5_delay_53_7;
  reg                 io_A_Valid_5_delay_54_6;
  reg                 io_A_Valid_5_delay_55_5;
  reg                 io_A_Valid_5_delay_56_4;
  reg                 io_A_Valid_5_delay_57_3;
  reg                 io_A_Valid_5_delay_58_2;
  reg                 io_A_Valid_5_delay_59_1;
  reg                 io_A_Valid_5_delay_60;
  reg                 io_B_Valid_60_delay_1_4;
  reg                 io_B_Valid_60_delay_2_3;
  reg                 io_B_Valid_60_delay_3_2;
  reg                 io_B_Valid_60_delay_4_1;
  reg                 io_B_Valid_60_delay_5;
  reg                 io_A_Valid_5_delay_1_60;
  reg                 io_A_Valid_5_delay_2_59;
  reg                 io_A_Valid_5_delay_3_58;
  reg                 io_A_Valid_5_delay_4_57;
  reg                 io_A_Valid_5_delay_5_56;
  reg                 io_A_Valid_5_delay_6_55;
  reg                 io_A_Valid_5_delay_7_54;
  reg                 io_A_Valid_5_delay_8_53;
  reg                 io_A_Valid_5_delay_9_52;
  reg                 io_A_Valid_5_delay_10_51;
  reg                 io_A_Valid_5_delay_11_50;
  reg                 io_A_Valid_5_delay_12_49;
  reg                 io_A_Valid_5_delay_13_48;
  reg                 io_A_Valid_5_delay_14_47;
  reg                 io_A_Valid_5_delay_15_46;
  reg                 io_A_Valid_5_delay_16_45;
  reg                 io_A_Valid_5_delay_17_44;
  reg                 io_A_Valid_5_delay_18_43;
  reg                 io_A_Valid_5_delay_19_42;
  reg                 io_A_Valid_5_delay_20_41;
  reg                 io_A_Valid_5_delay_21_40;
  reg                 io_A_Valid_5_delay_22_39;
  reg                 io_A_Valid_5_delay_23_38;
  reg                 io_A_Valid_5_delay_24_37;
  reg                 io_A_Valid_5_delay_25_36;
  reg                 io_A_Valid_5_delay_26_35;
  reg                 io_A_Valid_5_delay_27_34;
  reg                 io_A_Valid_5_delay_28_33;
  reg                 io_A_Valid_5_delay_29_32;
  reg                 io_A_Valid_5_delay_30_31;
  reg                 io_A_Valid_5_delay_31_30;
  reg                 io_A_Valid_5_delay_32_29;
  reg                 io_A_Valid_5_delay_33_28;
  reg                 io_A_Valid_5_delay_34_27;
  reg                 io_A_Valid_5_delay_35_26;
  reg                 io_A_Valid_5_delay_36_25;
  reg                 io_A_Valid_5_delay_37_24;
  reg                 io_A_Valid_5_delay_38_23;
  reg                 io_A_Valid_5_delay_39_22;
  reg                 io_A_Valid_5_delay_40_21;
  reg                 io_A_Valid_5_delay_41_20;
  reg                 io_A_Valid_5_delay_42_19;
  reg                 io_A_Valid_5_delay_43_18;
  reg                 io_A_Valid_5_delay_44_17;
  reg                 io_A_Valid_5_delay_45_16;
  reg                 io_A_Valid_5_delay_46_15;
  reg                 io_A_Valid_5_delay_47_14;
  reg                 io_A_Valid_5_delay_48_13;
  reg                 io_A_Valid_5_delay_49_12;
  reg                 io_A_Valid_5_delay_50_11;
  reg                 io_A_Valid_5_delay_51_10;
  reg                 io_A_Valid_5_delay_52_9;
  reg                 io_A_Valid_5_delay_53_8;
  reg                 io_A_Valid_5_delay_54_7;
  reg                 io_A_Valid_5_delay_55_6;
  reg                 io_A_Valid_5_delay_56_5;
  reg                 io_A_Valid_5_delay_57_4;
  reg                 io_A_Valid_5_delay_58_3;
  reg                 io_A_Valid_5_delay_59_2;
  reg                 io_A_Valid_5_delay_60_1;
  reg                 io_A_Valid_5_delay_61;
  reg                 io_B_Valid_61_delay_1_4;
  reg                 io_B_Valid_61_delay_2_3;
  reg                 io_B_Valid_61_delay_3_2;
  reg                 io_B_Valid_61_delay_4_1;
  reg                 io_B_Valid_61_delay_5;
  reg                 io_A_Valid_5_delay_1_61;
  reg                 io_A_Valid_5_delay_2_60;
  reg                 io_A_Valid_5_delay_3_59;
  reg                 io_A_Valid_5_delay_4_58;
  reg                 io_A_Valid_5_delay_5_57;
  reg                 io_A_Valid_5_delay_6_56;
  reg                 io_A_Valid_5_delay_7_55;
  reg                 io_A_Valid_5_delay_8_54;
  reg                 io_A_Valid_5_delay_9_53;
  reg                 io_A_Valid_5_delay_10_52;
  reg                 io_A_Valid_5_delay_11_51;
  reg                 io_A_Valid_5_delay_12_50;
  reg                 io_A_Valid_5_delay_13_49;
  reg                 io_A_Valid_5_delay_14_48;
  reg                 io_A_Valid_5_delay_15_47;
  reg                 io_A_Valid_5_delay_16_46;
  reg                 io_A_Valid_5_delay_17_45;
  reg                 io_A_Valid_5_delay_18_44;
  reg                 io_A_Valid_5_delay_19_43;
  reg                 io_A_Valid_5_delay_20_42;
  reg                 io_A_Valid_5_delay_21_41;
  reg                 io_A_Valid_5_delay_22_40;
  reg                 io_A_Valid_5_delay_23_39;
  reg                 io_A_Valid_5_delay_24_38;
  reg                 io_A_Valid_5_delay_25_37;
  reg                 io_A_Valid_5_delay_26_36;
  reg                 io_A_Valid_5_delay_27_35;
  reg                 io_A_Valid_5_delay_28_34;
  reg                 io_A_Valid_5_delay_29_33;
  reg                 io_A_Valid_5_delay_30_32;
  reg                 io_A_Valid_5_delay_31_31;
  reg                 io_A_Valid_5_delay_32_30;
  reg                 io_A_Valid_5_delay_33_29;
  reg                 io_A_Valid_5_delay_34_28;
  reg                 io_A_Valid_5_delay_35_27;
  reg                 io_A_Valid_5_delay_36_26;
  reg                 io_A_Valid_5_delay_37_25;
  reg                 io_A_Valid_5_delay_38_24;
  reg                 io_A_Valid_5_delay_39_23;
  reg                 io_A_Valid_5_delay_40_22;
  reg                 io_A_Valid_5_delay_41_21;
  reg                 io_A_Valid_5_delay_42_20;
  reg                 io_A_Valid_5_delay_43_19;
  reg                 io_A_Valid_5_delay_44_18;
  reg                 io_A_Valid_5_delay_45_17;
  reg                 io_A_Valid_5_delay_46_16;
  reg                 io_A_Valid_5_delay_47_15;
  reg                 io_A_Valid_5_delay_48_14;
  reg                 io_A_Valid_5_delay_49_13;
  reg                 io_A_Valid_5_delay_50_12;
  reg                 io_A_Valid_5_delay_51_11;
  reg                 io_A_Valid_5_delay_52_10;
  reg                 io_A_Valid_5_delay_53_9;
  reg                 io_A_Valid_5_delay_54_8;
  reg                 io_A_Valid_5_delay_55_7;
  reg                 io_A_Valid_5_delay_56_6;
  reg                 io_A_Valid_5_delay_57_5;
  reg                 io_A_Valid_5_delay_58_4;
  reg                 io_A_Valid_5_delay_59_3;
  reg                 io_A_Valid_5_delay_60_2;
  reg                 io_A_Valid_5_delay_61_1;
  reg                 io_A_Valid_5_delay_62;
  reg                 io_B_Valid_62_delay_1_4;
  reg                 io_B_Valid_62_delay_2_3;
  reg                 io_B_Valid_62_delay_3_2;
  reg                 io_B_Valid_62_delay_4_1;
  reg                 io_B_Valid_62_delay_5;
  reg                 io_A_Valid_5_delay_1_62;
  reg                 io_A_Valid_5_delay_2_61;
  reg                 io_A_Valid_5_delay_3_60;
  reg                 io_A_Valid_5_delay_4_59;
  reg                 io_A_Valid_5_delay_5_58;
  reg                 io_A_Valid_5_delay_6_57;
  reg                 io_A_Valid_5_delay_7_56;
  reg                 io_A_Valid_5_delay_8_55;
  reg                 io_A_Valid_5_delay_9_54;
  reg                 io_A_Valid_5_delay_10_53;
  reg                 io_A_Valid_5_delay_11_52;
  reg                 io_A_Valid_5_delay_12_51;
  reg                 io_A_Valid_5_delay_13_50;
  reg                 io_A_Valid_5_delay_14_49;
  reg                 io_A_Valid_5_delay_15_48;
  reg                 io_A_Valid_5_delay_16_47;
  reg                 io_A_Valid_5_delay_17_46;
  reg                 io_A_Valid_5_delay_18_45;
  reg                 io_A_Valid_5_delay_19_44;
  reg                 io_A_Valid_5_delay_20_43;
  reg                 io_A_Valid_5_delay_21_42;
  reg                 io_A_Valid_5_delay_22_41;
  reg                 io_A_Valid_5_delay_23_40;
  reg                 io_A_Valid_5_delay_24_39;
  reg                 io_A_Valid_5_delay_25_38;
  reg                 io_A_Valid_5_delay_26_37;
  reg                 io_A_Valid_5_delay_27_36;
  reg                 io_A_Valid_5_delay_28_35;
  reg                 io_A_Valid_5_delay_29_34;
  reg                 io_A_Valid_5_delay_30_33;
  reg                 io_A_Valid_5_delay_31_32;
  reg                 io_A_Valid_5_delay_32_31;
  reg                 io_A_Valid_5_delay_33_30;
  reg                 io_A_Valid_5_delay_34_29;
  reg                 io_A_Valid_5_delay_35_28;
  reg                 io_A_Valid_5_delay_36_27;
  reg                 io_A_Valid_5_delay_37_26;
  reg                 io_A_Valid_5_delay_38_25;
  reg                 io_A_Valid_5_delay_39_24;
  reg                 io_A_Valid_5_delay_40_23;
  reg                 io_A_Valid_5_delay_41_22;
  reg                 io_A_Valid_5_delay_42_21;
  reg                 io_A_Valid_5_delay_43_20;
  reg                 io_A_Valid_5_delay_44_19;
  reg                 io_A_Valid_5_delay_45_18;
  reg                 io_A_Valid_5_delay_46_17;
  reg                 io_A_Valid_5_delay_47_16;
  reg                 io_A_Valid_5_delay_48_15;
  reg                 io_A_Valid_5_delay_49_14;
  reg                 io_A_Valid_5_delay_50_13;
  reg                 io_A_Valid_5_delay_51_12;
  reg                 io_A_Valid_5_delay_52_11;
  reg                 io_A_Valid_5_delay_53_10;
  reg                 io_A_Valid_5_delay_54_9;
  reg                 io_A_Valid_5_delay_55_8;
  reg                 io_A_Valid_5_delay_56_7;
  reg                 io_A_Valid_5_delay_57_6;
  reg                 io_A_Valid_5_delay_58_5;
  reg                 io_A_Valid_5_delay_59_4;
  reg                 io_A_Valid_5_delay_60_3;
  reg                 io_A_Valid_5_delay_61_2;
  reg                 io_A_Valid_5_delay_62_1;
  reg                 io_A_Valid_5_delay_63;
  reg                 io_B_Valid_63_delay_1_4;
  reg                 io_B_Valid_63_delay_2_3;
  reg                 io_B_Valid_63_delay_3_2;
  reg                 io_B_Valid_63_delay_4_1;
  reg                 io_B_Valid_63_delay_5;
  reg        [15:0]   io_signCount_regNextWhen_6;
  reg                 io_B_Valid_0_delay_1_5;
  reg                 io_B_Valid_0_delay_2_4;
  reg                 io_B_Valid_0_delay_3_3;
  reg                 io_B_Valid_0_delay_4_2;
  reg                 io_B_Valid_0_delay_5_1;
  reg                 io_B_Valid_0_delay_6;
  reg                 io_A_Valid_6_delay_1;
  reg                 io_B_Valid_1_delay_1_5;
  reg                 io_B_Valid_1_delay_2_4;
  reg                 io_B_Valid_1_delay_3_3;
  reg                 io_B_Valid_1_delay_4_2;
  reg                 io_B_Valid_1_delay_5_1;
  reg                 io_B_Valid_1_delay_6;
  reg                 io_A_Valid_6_delay_1_1;
  reg                 io_A_Valid_6_delay_2;
  reg                 io_B_Valid_2_delay_1_5;
  reg                 io_B_Valid_2_delay_2_4;
  reg                 io_B_Valid_2_delay_3_3;
  reg                 io_B_Valid_2_delay_4_2;
  reg                 io_B_Valid_2_delay_5_1;
  reg                 io_B_Valid_2_delay_6;
  reg                 io_A_Valid_6_delay_1_2;
  reg                 io_A_Valid_6_delay_2_1;
  reg                 io_A_Valid_6_delay_3;
  reg                 io_B_Valid_3_delay_1_5;
  reg                 io_B_Valid_3_delay_2_4;
  reg                 io_B_Valid_3_delay_3_3;
  reg                 io_B_Valid_3_delay_4_2;
  reg                 io_B_Valid_3_delay_5_1;
  reg                 io_B_Valid_3_delay_6;
  reg                 io_A_Valid_6_delay_1_3;
  reg                 io_A_Valid_6_delay_2_2;
  reg                 io_A_Valid_6_delay_3_1;
  reg                 io_A_Valid_6_delay_4;
  reg                 io_B_Valid_4_delay_1_5;
  reg                 io_B_Valid_4_delay_2_4;
  reg                 io_B_Valid_4_delay_3_3;
  reg                 io_B_Valid_4_delay_4_2;
  reg                 io_B_Valid_4_delay_5_1;
  reg                 io_B_Valid_4_delay_6;
  reg                 io_A_Valid_6_delay_1_4;
  reg                 io_A_Valid_6_delay_2_3;
  reg                 io_A_Valid_6_delay_3_2;
  reg                 io_A_Valid_6_delay_4_1;
  reg                 io_A_Valid_6_delay_5;
  reg                 io_B_Valid_5_delay_1_5;
  reg                 io_B_Valid_5_delay_2_4;
  reg                 io_B_Valid_5_delay_3_3;
  reg                 io_B_Valid_5_delay_4_2;
  reg                 io_B_Valid_5_delay_5_1;
  reg                 io_B_Valid_5_delay_6;
  reg                 io_A_Valid_6_delay_1_5;
  reg                 io_A_Valid_6_delay_2_4;
  reg                 io_A_Valid_6_delay_3_3;
  reg                 io_A_Valid_6_delay_4_2;
  reg                 io_A_Valid_6_delay_5_1;
  reg                 io_A_Valid_6_delay_6;
  reg                 io_B_Valid_6_delay_1_5;
  reg                 io_B_Valid_6_delay_2_4;
  reg                 io_B_Valid_6_delay_3_3;
  reg                 io_B_Valid_6_delay_4_2;
  reg                 io_B_Valid_6_delay_5_1;
  reg                 io_B_Valid_6_delay_6;
  reg                 io_A_Valid_6_delay_1_6;
  reg                 io_A_Valid_6_delay_2_5;
  reg                 io_A_Valid_6_delay_3_4;
  reg                 io_A_Valid_6_delay_4_3;
  reg                 io_A_Valid_6_delay_5_2;
  reg                 io_A_Valid_6_delay_6_1;
  reg                 io_A_Valid_6_delay_7;
  reg                 io_B_Valid_7_delay_1_5;
  reg                 io_B_Valid_7_delay_2_4;
  reg                 io_B_Valid_7_delay_3_3;
  reg                 io_B_Valid_7_delay_4_2;
  reg                 io_B_Valid_7_delay_5_1;
  reg                 io_B_Valid_7_delay_6;
  reg                 io_A_Valid_6_delay_1_7;
  reg                 io_A_Valid_6_delay_2_6;
  reg                 io_A_Valid_6_delay_3_5;
  reg                 io_A_Valid_6_delay_4_4;
  reg                 io_A_Valid_6_delay_5_3;
  reg                 io_A_Valid_6_delay_6_2;
  reg                 io_A_Valid_6_delay_7_1;
  reg                 io_A_Valid_6_delay_8;
  reg                 io_B_Valid_8_delay_1_5;
  reg                 io_B_Valid_8_delay_2_4;
  reg                 io_B_Valid_8_delay_3_3;
  reg                 io_B_Valid_8_delay_4_2;
  reg                 io_B_Valid_8_delay_5_1;
  reg                 io_B_Valid_8_delay_6;
  reg                 io_A_Valid_6_delay_1_8;
  reg                 io_A_Valid_6_delay_2_7;
  reg                 io_A_Valid_6_delay_3_6;
  reg                 io_A_Valid_6_delay_4_5;
  reg                 io_A_Valid_6_delay_5_4;
  reg                 io_A_Valid_6_delay_6_3;
  reg                 io_A_Valid_6_delay_7_2;
  reg                 io_A_Valid_6_delay_8_1;
  reg                 io_A_Valid_6_delay_9;
  reg                 io_B_Valid_9_delay_1_5;
  reg                 io_B_Valid_9_delay_2_4;
  reg                 io_B_Valid_9_delay_3_3;
  reg                 io_B_Valid_9_delay_4_2;
  reg                 io_B_Valid_9_delay_5_1;
  reg                 io_B_Valid_9_delay_6;
  reg                 io_A_Valid_6_delay_1_9;
  reg                 io_A_Valid_6_delay_2_8;
  reg                 io_A_Valid_6_delay_3_7;
  reg                 io_A_Valid_6_delay_4_6;
  reg                 io_A_Valid_6_delay_5_5;
  reg                 io_A_Valid_6_delay_6_4;
  reg                 io_A_Valid_6_delay_7_3;
  reg                 io_A_Valid_6_delay_8_2;
  reg                 io_A_Valid_6_delay_9_1;
  reg                 io_A_Valid_6_delay_10;
  reg                 io_B_Valid_10_delay_1_5;
  reg                 io_B_Valid_10_delay_2_4;
  reg                 io_B_Valid_10_delay_3_3;
  reg                 io_B_Valid_10_delay_4_2;
  reg                 io_B_Valid_10_delay_5_1;
  reg                 io_B_Valid_10_delay_6;
  reg                 io_A_Valid_6_delay_1_10;
  reg                 io_A_Valid_6_delay_2_9;
  reg                 io_A_Valid_6_delay_3_8;
  reg                 io_A_Valid_6_delay_4_7;
  reg                 io_A_Valid_6_delay_5_6;
  reg                 io_A_Valid_6_delay_6_5;
  reg                 io_A_Valid_6_delay_7_4;
  reg                 io_A_Valid_6_delay_8_3;
  reg                 io_A_Valid_6_delay_9_2;
  reg                 io_A_Valid_6_delay_10_1;
  reg                 io_A_Valid_6_delay_11;
  reg                 io_B_Valid_11_delay_1_5;
  reg                 io_B_Valid_11_delay_2_4;
  reg                 io_B_Valid_11_delay_3_3;
  reg                 io_B_Valid_11_delay_4_2;
  reg                 io_B_Valid_11_delay_5_1;
  reg                 io_B_Valid_11_delay_6;
  reg                 io_A_Valid_6_delay_1_11;
  reg                 io_A_Valid_6_delay_2_10;
  reg                 io_A_Valid_6_delay_3_9;
  reg                 io_A_Valid_6_delay_4_8;
  reg                 io_A_Valid_6_delay_5_7;
  reg                 io_A_Valid_6_delay_6_6;
  reg                 io_A_Valid_6_delay_7_5;
  reg                 io_A_Valid_6_delay_8_4;
  reg                 io_A_Valid_6_delay_9_3;
  reg                 io_A_Valid_6_delay_10_2;
  reg                 io_A_Valid_6_delay_11_1;
  reg                 io_A_Valid_6_delay_12;
  reg                 io_B_Valid_12_delay_1_5;
  reg                 io_B_Valid_12_delay_2_4;
  reg                 io_B_Valid_12_delay_3_3;
  reg                 io_B_Valid_12_delay_4_2;
  reg                 io_B_Valid_12_delay_5_1;
  reg                 io_B_Valid_12_delay_6;
  reg                 io_A_Valid_6_delay_1_12;
  reg                 io_A_Valid_6_delay_2_11;
  reg                 io_A_Valid_6_delay_3_10;
  reg                 io_A_Valid_6_delay_4_9;
  reg                 io_A_Valid_6_delay_5_8;
  reg                 io_A_Valid_6_delay_6_7;
  reg                 io_A_Valid_6_delay_7_6;
  reg                 io_A_Valid_6_delay_8_5;
  reg                 io_A_Valid_6_delay_9_4;
  reg                 io_A_Valid_6_delay_10_3;
  reg                 io_A_Valid_6_delay_11_2;
  reg                 io_A_Valid_6_delay_12_1;
  reg                 io_A_Valid_6_delay_13;
  reg                 io_B_Valid_13_delay_1_5;
  reg                 io_B_Valid_13_delay_2_4;
  reg                 io_B_Valid_13_delay_3_3;
  reg                 io_B_Valid_13_delay_4_2;
  reg                 io_B_Valid_13_delay_5_1;
  reg                 io_B_Valid_13_delay_6;
  reg                 io_A_Valid_6_delay_1_13;
  reg                 io_A_Valid_6_delay_2_12;
  reg                 io_A_Valid_6_delay_3_11;
  reg                 io_A_Valid_6_delay_4_10;
  reg                 io_A_Valid_6_delay_5_9;
  reg                 io_A_Valid_6_delay_6_8;
  reg                 io_A_Valid_6_delay_7_7;
  reg                 io_A_Valid_6_delay_8_6;
  reg                 io_A_Valid_6_delay_9_5;
  reg                 io_A_Valid_6_delay_10_4;
  reg                 io_A_Valid_6_delay_11_3;
  reg                 io_A_Valid_6_delay_12_2;
  reg                 io_A_Valid_6_delay_13_1;
  reg                 io_A_Valid_6_delay_14;
  reg                 io_B_Valid_14_delay_1_5;
  reg                 io_B_Valid_14_delay_2_4;
  reg                 io_B_Valid_14_delay_3_3;
  reg                 io_B_Valid_14_delay_4_2;
  reg                 io_B_Valid_14_delay_5_1;
  reg                 io_B_Valid_14_delay_6;
  reg                 io_A_Valid_6_delay_1_14;
  reg                 io_A_Valid_6_delay_2_13;
  reg                 io_A_Valid_6_delay_3_12;
  reg                 io_A_Valid_6_delay_4_11;
  reg                 io_A_Valid_6_delay_5_10;
  reg                 io_A_Valid_6_delay_6_9;
  reg                 io_A_Valid_6_delay_7_8;
  reg                 io_A_Valid_6_delay_8_7;
  reg                 io_A_Valid_6_delay_9_6;
  reg                 io_A_Valid_6_delay_10_5;
  reg                 io_A_Valid_6_delay_11_4;
  reg                 io_A_Valid_6_delay_12_3;
  reg                 io_A_Valid_6_delay_13_2;
  reg                 io_A_Valid_6_delay_14_1;
  reg                 io_A_Valid_6_delay_15;
  reg                 io_B_Valid_15_delay_1_5;
  reg                 io_B_Valid_15_delay_2_4;
  reg                 io_B_Valid_15_delay_3_3;
  reg                 io_B_Valid_15_delay_4_2;
  reg                 io_B_Valid_15_delay_5_1;
  reg                 io_B_Valid_15_delay_6;
  reg                 io_A_Valid_6_delay_1_15;
  reg                 io_A_Valid_6_delay_2_14;
  reg                 io_A_Valid_6_delay_3_13;
  reg                 io_A_Valid_6_delay_4_12;
  reg                 io_A_Valid_6_delay_5_11;
  reg                 io_A_Valid_6_delay_6_10;
  reg                 io_A_Valid_6_delay_7_9;
  reg                 io_A_Valid_6_delay_8_8;
  reg                 io_A_Valid_6_delay_9_7;
  reg                 io_A_Valid_6_delay_10_6;
  reg                 io_A_Valid_6_delay_11_5;
  reg                 io_A_Valid_6_delay_12_4;
  reg                 io_A_Valid_6_delay_13_3;
  reg                 io_A_Valid_6_delay_14_2;
  reg                 io_A_Valid_6_delay_15_1;
  reg                 io_A_Valid_6_delay_16;
  reg                 io_B_Valid_16_delay_1_5;
  reg                 io_B_Valid_16_delay_2_4;
  reg                 io_B_Valid_16_delay_3_3;
  reg                 io_B_Valid_16_delay_4_2;
  reg                 io_B_Valid_16_delay_5_1;
  reg                 io_B_Valid_16_delay_6;
  reg                 io_A_Valid_6_delay_1_16;
  reg                 io_A_Valid_6_delay_2_15;
  reg                 io_A_Valid_6_delay_3_14;
  reg                 io_A_Valid_6_delay_4_13;
  reg                 io_A_Valid_6_delay_5_12;
  reg                 io_A_Valid_6_delay_6_11;
  reg                 io_A_Valid_6_delay_7_10;
  reg                 io_A_Valid_6_delay_8_9;
  reg                 io_A_Valid_6_delay_9_8;
  reg                 io_A_Valid_6_delay_10_7;
  reg                 io_A_Valid_6_delay_11_6;
  reg                 io_A_Valid_6_delay_12_5;
  reg                 io_A_Valid_6_delay_13_4;
  reg                 io_A_Valid_6_delay_14_3;
  reg                 io_A_Valid_6_delay_15_2;
  reg                 io_A_Valid_6_delay_16_1;
  reg                 io_A_Valid_6_delay_17;
  reg                 io_B_Valid_17_delay_1_5;
  reg                 io_B_Valid_17_delay_2_4;
  reg                 io_B_Valid_17_delay_3_3;
  reg                 io_B_Valid_17_delay_4_2;
  reg                 io_B_Valid_17_delay_5_1;
  reg                 io_B_Valid_17_delay_6;
  reg                 io_A_Valid_6_delay_1_17;
  reg                 io_A_Valid_6_delay_2_16;
  reg                 io_A_Valid_6_delay_3_15;
  reg                 io_A_Valid_6_delay_4_14;
  reg                 io_A_Valid_6_delay_5_13;
  reg                 io_A_Valid_6_delay_6_12;
  reg                 io_A_Valid_6_delay_7_11;
  reg                 io_A_Valid_6_delay_8_10;
  reg                 io_A_Valid_6_delay_9_9;
  reg                 io_A_Valid_6_delay_10_8;
  reg                 io_A_Valid_6_delay_11_7;
  reg                 io_A_Valid_6_delay_12_6;
  reg                 io_A_Valid_6_delay_13_5;
  reg                 io_A_Valid_6_delay_14_4;
  reg                 io_A_Valid_6_delay_15_3;
  reg                 io_A_Valid_6_delay_16_2;
  reg                 io_A_Valid_6_delay_17_1;
  reg                 io_A_Valid_6_delay_18;
  reg                 io_B_Valid_18_delay_1_5;
  reg                 io_B_Valid_18_delay_2_4;
  reg                 io_B_Valid_18_delay_3_3;
  reg                 io_B_Valid_18_delay_4_2;
  reg                 io_B_Valid_18_delay_5_1;
  reg                 io_B_Valid_18_delay_6;
  reg                 io_A_Valid_6_delay_1_18;
  reg                 io_A_Valid_6_delay_2_17;
  reg                 io_A_Valid_6_delay_3_16;
  reg                 io_A_Valid_6_delay_4_15;
  reg                 io_A_Valid_6_delay_5_14;
  reg                 io_A_Valid_6_delay_6_13;
  reg                 io_A_Valid_6_delay_7_12;
  reg                 io_A_Valid_6_delay_8_11;
  reg                 io_A_Valid_6_delay_9_10;
  reg                 io_A_Valid_6_delay_10_9;
  reg                 io_A_Valid_6_delay_11_8;
  reg                 io_A_Valid_6_delay_12_7;
  reg                 io_A_Valid_6_delay_13_6;
  reg                 io_A_Valid_6_delay_14_5;
  reg                 io_A_Valid_6_delay_15_4;
  reg                 io_A_Valid_6_delay_16_3;
  reg                 io_A_Valid_6_delay_17_2;
  reg                 io_A_Valid_6_delay_18_1;
  reg                 io_A_Valid_6_delay_19;
  reg                 io_B_Valid_19_delay_1_5;
  reg                 io_B_Valid_19_delay_2_4;
  reg                 io_B_Valid_19_delay_3_3;
  reg                 io_B_Valid_19_delay_4_2;
  reg                 io_B_Valid_19_delay_5_1;
  reg                 io_B_Valid_19_delay_6;
  reg                 io_A_Valid_6_delay_1_19;
  reg                 io_A_Valid_6_delay_2_18;
  reg                 io_A_Valid_6_delay_3_17;
  reg                 io_A_Valid_6_delay_4_16;
  reg                 io_A_Valid_6_delay_5_15;
  reg                 io_A_Valid_6_delay_6_14;
  reg                 io_A_Valid_6_delay_7_13;
  reg                 io_A_Valid_6_delay_8_12;
  reg                 io_A_Valid_6_delay_9_11;
  reg                 io_A_Valid_6_delay_10_10;
  reg                 io_A_Valid_6_delay_11_9;
  reg                 io_A_Valid_6_delay_12_8;
  reg                 io_A_Valid_6_delay_13_7;
  reg                 io_A_Valid_6_delay_14_6;
  reg                 io_A_Valid_6_delay_15_5;
  reg                 io_A_Valid_6_delay_16_4;
  reg                 io_A_Valid_6_delay_17_3;
  reg                 io_A_Valid_6_delay_18_2;
  reg                 io_A_Valid_6_delay_19_1;
  reg                 io_A_Valid_6_delay_20;
  reg                 io_B_Valid_20_delay_1_5;
  reg                 io_B_Valid_20_delay_2_4;
  reg                 io_B_Valid_20_delay_3_3;
  reg                 io_B_Valid_20_delay_4_2;
  reg                 io_B_Valid_20_delay_5_1;
  reg                 io_B_Valid_20_delay_6;
  reg                 io_A_Valid_6_delay_1_20;
  reg                 io_A_Valid_6_delay_2_19;
  reg                 io_A_Valid_6_delay_3_18;
  reg                 io_A_Valid_6_delay_4_17;
  reg                 io_A_Valid_6_delay_5_16;
  reg                 io_A_Valid_6_delay_6_15;
  reg                 io_A_Valid_6_delay_7_14;
  reg                 io_A_Valid_6_delay_8_13;
  reg                 io_A_Valid_6_delay_9_12;
  reg                 io_A_Valid_6_delay_10_11;
  reg                 io_A_Valid_6_delay_11_10;
  reg                 io_A_Valid_6_delay_12_9;
  reg                 io_A_Valid_6_delay_13_8;
  reg                 io_A_Valid_6_delay_14_7;
  reg                 io_A_Valid_6_delay_15_6;
  reg                 io_A_Valid_6_delay_16_5;
  reg                 io_A_Valid_6_delay_17_4;
  reg                 io_A_Valid_6_delay_18_3;
  reg                 io_A_Valid_6_delay_19_2;
  reg                 io_A_Valid_6_delay_20_1;
  reg                 io_A_Valid_6_delay_21;
  reg                 io_B_Valid_21_delay_1_5;
  reg                 io_B_Valid_21_delay_2_4;
  reg                 io_B_Valid_21_delay_3_3;
  reg                 io_B_Valid_21_delay_4_2;
  reg                 io_B_Valid_21_delay_5_1;
  reg                 io_B_Valid_21_delay_6;
  reg                 io_A_Valid_6_delay_1_21;
  reg                 io_A_Valid_6_delay_2_20;
  reg                 io_A_Valid_6_delay_3_19;
  reg                 io_A_Valid_6_delay_4_18;
  reg                 io_A_Valid_6_delay_5_17;
  reg                 io_A_Valid_6_delay_6_16;
  reg                 io_A_Valid_6_delay_7_15;
  reg                 io_A_Valid_6_delay_8_14;
  reg                 io_A_Valid_6_delay_9_13;
  reg                 io_A_Valid_6_delay_10_12;
  reg                 io_A_Valid_6_delay_11_11;
  reg                 io_A_Valid_6_delay_12_10;
  reg                 io_A_Valid_6_delay_13_9;
  reg                 io_A_Valid_6_delay_14_8;
  reg                 io_A_Valid_6_delay_15_7;
  reg                 io_A_Valid_6_delay_16_6;
  reg                 io_A_Valid_6_delay_17_5;
  reg                 io_A_Valid_6_delay_18_4;
  reg                 io_A_Valid_6_delay_19_3;
  reg                 io_A_Valid_6_delay_20_2;
  reg                 io_A_Valid_6_delay_21_1;
  reg                 io_A_Valid_6_delay_22;
  reg                 io_B_Valid_22_delay_1_5;
  reg                 io_B_Valid_22_delay_2_4;
  reg                 io_B_Valid_22_delay_3_3;
  reg                 io_B_Valid_22_delay_4_2;
  reg                 io_B_Valid_22_delay_5_1;
  reg                 io_B_Valid_22_delay_6;
  reg                 io_A_Valid_6_delay_1_22;
  reg                 io_A_Valid_6_delay_2_21;
  reg                 io_A_Valid_6_delay_3_20;
  reg                 io_A_Valid_6_delay_4_19;
  reg                 io_A_Valid_6_delay_5_18;
  reg                 io_A_Valid_6_delay_6_17;
  reg                 io_A_Valid_6_delay_7_16;
  reg                 io_A_Valid_6_delay_8_15;
  reg                 io_A_Valid_6_delay_9_14;
  reg                 io_A_Valid_6_delay_10_13;
  reg                 io_A_Valid_6_delay_11_12;
  reg                 io_A_Valid_6_delay_12_11;
  reg                 io_A_Valid_6_delay_13_10;
  reg                 io_A_Valid_6_delay_14_9;
  reg                 io_A_Valid_6_delay_15_8;
  reg                 io_A_Valid_6_delay_16_7;
  reg                 io_A_Valid_6_delay_17_6;
  reg                 io_A_Valid_6_delay_18_5;
  reg                 io_A_Valid_6_delay_19_4;
  reg                 io_A_Valid_6_delay_20_3;
  reg                 io_A_Valid_6_delay_21_2;
  reg                 io_A_Valid_6_delay_22_1;
  reg                 io_A_Valid_6_delay_23;
  reg                 io_B_Valid_23_delay_1_5;
  reg                 io_B_Valid_23_delay_2_4;
  reg                 io_B_Valid_23_delay_3_3;
  reg                 io_B_Valid_23_delay_4_2;
  reg                 io_B_Valid_23_delay_5_1;
  reg                 io_B_Valid_23_delay_6;
  reg                 io_A_Valid_6_delay_1_23;
  reg                 io_A_Valid_6_delay_2_22;
  reg                 io_A_Valid_6_delay_3_21;
  reg                 io_A_Valid_6_delay_4_20;
  reg                 io_A_Valid_6_delay_5_19;
  reg                 io_A_Valid_6_delay_6_18;
  reg                 io_A_Valid_6_delay_7_17;
  reg                 io_A_Valid_6_delay_8_16;
  reg                 io_A_Valid_6_delay_9_15;
  reg                 io_A_Valid_6_delay_10_14;
  reg                 io_A_Valid_6_delay_11_13;
  reg                 io_A_Valid_6_delay_12_12;
  reg                 io_A_Valid_6_delay_13_11;
  reg                 io_A_Valid_6_delay_14_10;
  reg                 io_A_Valid_6_delay_15_9;
  reg                 io_A_Valid_6_delay_16_8;
  reg                 io_A_Valid_6_delay_17_7;
  reg                 io_A_Valid_6_delay_18_6;
  reg                 io_A_Valid_6_delay_19_5;
  reg                 io_A_Valid_6_delay_20_4;
  reg                 io_A_Valid_6_delay_21_3;
  reg                 io_A_Valid_6_delay_22_2;
  reg                 io_A_Valid_6_delay_23_1;
  reg                 io_A_Valid_6_delay_24;
  reg                 io_B_Valid_24_delay_1_5;
  reg                 io_B_Valid_24_delay_2_4;
  reg                 io_B_Valid_24_delay_3_3;
  reg                 io_B_Valid_24_delay_4_2;
  reg                 io_B_Valid_24_delay_5_1;
  reg                 io_B_Valid_24_delay_6;
  reg                 io_A_Valid_6_delay_1_24;
  reg                 io_A_Valid_6_delay_2_23;
  reg                 io_A_Valid_6_delay_3_22;
  reg                 io_A_Valid_6_delay_4_21;
  reg                 io_A_Valid_6_delay_5_20;
  reg                 io_A_Valid_6_delay_6_19;
  reg                 io_A_Valid_6_delay_7_18;
  reg                 io_A_Valid_6_delay_8_17;
  reg                 io_A_Valid_6_delay_9_16;
  reg                 io_A_Valid_6_delay_10_15;
  reg                 io_A_Valid_6_delay_11_14;
  reg                 io_A_Valid_6_delay_12_13;
  reg                 io_A_Valid_6_delay_13_12;
  reg                 io_A_Valid_6_delay_14_11;
  reg                 io_A_Valid_6_delay_15_10;
  reg                 io_A_Valid_6_delay_16_9;
  reg                 io_A_Valid_6_delay_17_8;
  reg                 io_A_Valid_6_delay_18_7;
  reg                 io_A_Valid_6_delay_19_6;
  reg                 io_A_Valid_6_delay_20_5;
  reg                 io_A_Valid_6_delay_21_4;
  reg                 io_A_Valid_6_delay_22_3;
  reg                 io_A_Valid_6_delay_23_2;
  reg                 io_A_Valid_6_delay_24_1;
  reg                 io_A_Valid_6_delay_25;
  reg                 io_B_Valid_25_delay_1_5;
  reg                 io_B_Valid_25_delay_2_4;
  reg                 io_B_Valid_25_delay_3_3;
  reg                 io_B_Valid_25_delay_4_2;
  reg                 io_B_Valid_25_delay_5_1;
  reg                 io_B_Valid_25_delay_6;
  reg                 io_A_Valid_6_delay_1_25;
  reg                 io_A_Valid_6_delay_2_24;
  reg                 io_A_Valid_6_delay_3_23;
  reg                 io_A_Valid_6_delay_4_22;
  reg                 io_A_Valid_6_delay_5_21;
  reg                 io_A_Valid_6_delay_6_20;
  reg                 io_A_Valid_6_delay_7_19;
  reg                 io_A_Valid_6_delay_8_18;
  reg                 io_A_Valid_6_delay_9_17;
  reg                 io_A_Valid_6_delay_10_16;
  reg                 io_A_Valid_6_delay_11_15;
  reg                 io_A_Valid_6_delay_12_14;
  reg                 io_A_Valid_6_delay_13_13;
  reg                 io_A_Valid_6_delay_14_12;
  reg                 io_A_Valid_6_delay_15_11;
  reg                 io_A_Valid_6_delay_16_10;
  reg                 io_A_Valid_6_delay_17_9;
  reg                 io_A_Valid_6_delay_18_8;
  reg                 io_A_Valid_6_delay_19_7;
  reg                 io_A_Valid_6_delay_20_6;
  reg                 io_A_Valid_6_delay_21_5;
  reg                 io_A_Valid_6_delay_22_4;
  reg                 io_A_Valid_6_delay_23_3;
  reg                 io_A_Valid_6_delay_24_2;
  reg                 io_A_Valid_6_delay_25_1;
  reg                 io_A_Valid_6_delay_26;
  reg                 io_B_Valid_26_delay_1_5;
  reg                 io_B_Valid_26_delay_2_4;
  reg                 io_B_Valid_26_delay_3_3;
  reg                 io_B_Valid_26_delay_4_2;
  reg                 io_B_Valid_26_delay_5_1;
  reg                 io_B_Valid_26_delay_6;
  reg                 io_A_Valid_6_delay_1_26;
  reg                 io_A_Valid_6_delay_2_25;
  reg                 io_A_Valid_6_delay_3_24;
  reg                 io_A_Valid_6_delay_4_23;
  reg                 io_A_Valid_6_delay_5_22;
  reg                 io_A_Valid_6_delay_6_21;
  reg                 io_A_Valid_6_delay_7_20;
  reg                 io_A_Valid_6_delay_8_19;
  reg                 io_A_Valid_6_delay_9_18;
  reg                 io_A_Valid_6_delay_10_17;
  reg                 io_A_Valid_6_delay_11_16;
  reg                 io_A_Valid_6_delay_12_15;
  reg                 io_A_Valid_6_delay_13_14;
  reg                 io_A_Valid_6_delay_14_13;
  reg                 io_A_Valid_6_delay_15_12;
  reg                 io_A_Valid_6_delay_16_11;
  reg                 io_A_Valid_6_delay_17_10;
  reg                 io_A_Valid_6_delay_18_9;
  reg                 io_A_Valid_6_delay_19_8;
  reg                 io_A_Valid_6_delay_20_7;
  reg                 io_A_Valid_6_delay_21_6;
  reg                 io_A_Valid_6_delay_22_5;
  reg                 io_A_Valid_6_delay_23_4;
  reg                 io_A_Valid_6_delay_24_3;
  reg                 io_A_Valid_6_delay_25_2;
  reg                 io_A_Valid_6_delay_26_1;
  reg                 io_A_Valid_6_delay_27;
  reg                 io_B_Valid_27_delay_1_5;
  reg                 io_B_Valid_27_delay_2_4;
  reg                 io_B_Valid_27_delay_3_3;
  reg                 io_B_Valid_27_delay_4_2;
  reg                 io_B_Valid_27_delay_5_1;
  reg                 io_B_Valid_27_delay_6;
  reg                 io_A_Valid_6_delay_1_27;
  reg                 io_A_Valid_6_delay_2_26;
  reg                 io_A_Valid_6_delay_3_25;
  reg                 io_A_Valid_6_delay_4_24;
  reg                 io_A_Valid_6_delay_5_23;
  reg                 io_A_Valid_6_delay_6_22;
  reg                 io_A_Valid_6_delay_7_21;
  reg                 io_A_Valid_6_delay_8_20;
  reg                 io_A_Valid_6_delay_9_19;
  reg                 io_A_Valid_6_delay_10_18;
  reg                 io_A_Valid_6_delay_11_17;
  reg                 io_A_Valid_6_delay_12_16;
  reg                 io_A_Valid_6_delay_13_15;
  reg                 io_A_Valid_6_delay_14_14;
  reg                 io_A_Valid_6_delay_15_13;
  reg                 io_A_Valid_6_delay_16_12;
  reg                 io_A_Valid_6_delay_17_11;
  reg                 io_A_Valid_6_delay_18_10;
  reg                 io_A_Valid_6_delay_19_9;
  reg                 io_A_Valid_6_delay_20_8;
  reg                 io_A_Valid_6_delay_21_7;
  reg                 io_A_Valid_6_delay_22_6;
  reg                 io_A_Valid_6_delay_23_5;
  reg                 io_A_Valid_6_delay_24_4;
  reg                 io_A_Valid_6_delay_25_3;
  reg                 io_A_Valid_6_delay_26_2;
  reg                 io_A_Valid_6_delay_27_1;
  reg                 io_A_Valid_6_delay_28;
  reg                 io_B_Valid_28_delay_1_5;
  reg                 io_B_Valid_28_delay_2_4;
  reg                 io_B_Valid_28_delay_3_3;
  reg                 io_B_Valid_28_delay_4_2;
  reg                 io_B_Valid_28_delay_5_1;
  reg                 io_B_Valid_28_delay_6;
  reg                 io_A_Valid_6_delay_1_28;
  reg                 io_A_Valid_6_delay_2_27;
  reg                 io_A_Valid_6_delay_3_26;
  reg                 io_A_Valid_6_delay_4_25;
  reg                 io_A_Valid_6_delay_5_24;
  reg                 io_A_Valid_6_delay_6_23;
  reg                 io_A_Valid_6_delay_7_22;
  reg                 io_A_Valid_6_delay_8_21;
  reg                 io_A_Valid_6_delay_9_20;
  reg                 io_A_Valid_6_delay_10_19;
  reg                 io_A_Valid_6_delay_11_18;
  reg                 io_A_Valid_6_delay_12_17;
  reg                 io_A_Valid_6_delay_13_16;
  reg                 io_A_Valid_6_delay_14_15;
  reg                 io_A_Valid_6_delay_15_14;
  reg                 io_A_Valid_6_delay_16_13;
  reg                 io_A_Valid_6_delay_17_12;
  reg                 io_A_Valid_6_delay_18_11;
  reg                 io_A_Valid_6_delay_19_10;
  reg                 io_A_Valid_6_delay_20_9;
  reg                 io_A_Valid_6_delay_21_8;
  reg                 io_A_Valid_6_delay_22_7;
  reg                 io_A_Valid_6_delay_23_6;
  reg                 io_A_Valid_6_delay_24_5;
  reg                 io_A_Valid_6_delay_25_4;
  reg                 io_A_Valid_6_delay_26_3;
  reg                 io_A_Valid_6_delay_27_2;
  reg                 io_A_Valid_6_delay_28_1;
  reg                 io_A_Valid_6_delay_29;
  reg                 io_B_Valid_29_delay_1_5;
  reg                 io_B_Valid_29_delay_2_4;
  reg                 io_B_Valid_29_delay_3_3;
  reg                 io_B_Valid_29_delay_4_2;
  reg                 io_B_Valid_29_delay_5_1;
  reg                 io_B_Valid_29_delay_6;
  reg                 io_A_Valid_6_delay_1_29;
  reg                 io_A_Valid_6_delay_2_28;
  reg                 io_A_Valid_6_delay_3_27;
  reg                 io_A_Valid_6_delay_4_26;
  reg                 io_A_Valid_6_delay_5_25;
  reg                 io_A_Valid_6_delay_6_24;
  reg                 io_A_Valid_6_delay_7_23;
  reg                 io_A_Valid_6_delay_8_22;
  reg                 io_A_Valid_6_delay_9_21;
  reg                 io_A_Valid_6_delay_10_20;
  reg                 io_A_Valid_6_delay_11_19;
  reg                 io_A_Valid_6_delay_12_18;
  reg                 io_A_Valid_6_delay_13_17;
  reg                 io_A_Valid_6_delay_14_16;
  reg                 io_A_Valid_6_delay_15_15;
  reg                 io_A_Valid_6_delay_16_14;
  reg                 io_A_Valid_6_delay_17_13;
  reg                 io_A_Valid_6_delay_18_12;
  reg                 io_A_Valid_6_delay_19_11;
  reg                 io_A_Valid_6_delay_20_10;
  reg                 io_A_Valid_6_delay_21_9;
  reg                 io_A_Valid_6_delay_22_8;
  reg                 io_A_Valid_6_delay_23_7;
  reg                 io_A_Valid_6_delay_24_6;
  reg                 io_A_Valid_6_delay_25_5;
  reg                 io_A_Valid_6_delay_26_4;
  reg                 io_A_Valid_6_delay_27_3;
  reg                 io_A_Valid_6_delay_28_2;
  reg                 io_A_Valid_6_delay_29_1;
  reg                 io_A_Valid_6_delay_30;
  reg                 io_B_Valid_30_delay_1_5;
  reg                 io_B_Valid_30_delay_2_4;
  reg                 io_B_Valid_30_delay_3_3;
  reg                 io_B_Valid_30_delay_4_2;
  reg                 io_B_Valid_30_delay_5_1;
  reg                 io_B_Valid_30_delay_6;
  reg                 io_A_Valid_6_delay_1_30;
  reg                 io_A_Valid_6_delay_2_29;
  reg                 io_A_Valid_6_delay_3_28;
  reg                 io_A_Valid_6_delay_4_27;
  reg                 io_A_Valid_6_delay_5_26;
  reg                 io_A_Valid_6_delay_6_25;
  reg                 io_A_Valid_6_delay_7_24;
  reg                 io_A_Valid_6_delay_8_23;
  reg                 io_A_Valid_6_delay_9_22;
  reg                 io_A_Valid_6_delay_10_21;
  reg                 io_A_Valid_6_delay_11_20;
  reg                 io_A_Valid_6_delay_12_19;
  reg                 io_A_Valid_6_delay_13_18;
  reg                 io_A_Valid_6_delay_14_17;
  reg                 io_A_Valid_6_delay_15_16;
  reg                 io_A_Valid_6_delay_16_15;
  reg                 io_A_Valid_6_delay_17_14;
  reg                 io_A_Valid_6_delay_18_13;
  reg                 io_A_Valid_6_delay_19_12;
  reg                 io_A_Valid_6_delay_20_11;
  reg                 io_A_Valid_6_delay_21_10;
  reg                 io_A_Valid_6_delay_22_9;
  reg                 io_A_Valid_6_delay_23_8;
  reg                 io_A_Valid_6_delay_24_7;
  reg                 io_A_Valid_6_delay_25_6;
  reg                 io_A_Valid_6_delay_26_5;
  reg                 io_A_Valid_6_delay_27_4;
  reg                 io_A_Valid_6_delay_28_3;
  reg                 io_A_Valid_6_delay_29_2;
  reg                 io_A_Valid_6_delay_30_1;
  reg                 io_A_Valid_6_delay_31;
  reg                 io_B_Valid_31_delay_1_5;
  reg                 io_B_Valid_31_delay_2_4;
  reg                 io_B_Valid_31_delay_3_3;
  reg                 io_B_Valid_31_delay_4_2;
  reg                 io_B_Valid_31_delay_5_1;
  reg                 io_B_Valid_31_delay_6;
  reg                 io_A_Valid_6_delay_1_31;
  reg                 io_A_Valid_6_delay_2_30;
  reg                 io_A_Valid_6_delay_3_29;
  reg                 io_A_Valid_6_delay_4_28;
  reg                 io_A_Valid_6_delay_5_27;
  reg                 io_A_Valid_6_delay_6_26;
  reg                 io_A_Valid_6_delay_7_25;
  reg                 io_A_Valid_6_delay_8_24;
  reg                 io_A_Valid_6_delay_9_23;
  reg                 io_A_Valid_6_delay_10_22;
  reg                 io_A_Valid_6_delay_11_21;
  reg                 io_A_Valid_6_delay_12_20;
  reg                 io_A_Valid_6_delay_13_19;
  reg                 io_A_Valid_6_delay_14_18;
  reg                 io_A_Valid_6_delay_15_17;
  reg                 io_A_Valid_6_delay_16_16;
  reg                 io_A_Valid_6_delay_17_15;
  reg                 io_A_Valid_6_delay_18_14;
  reg                 io_A_Valid_6_delay_19_13;
  reg                 io_A_Valid_6_delay_20_12;
  reg                 io_A_Valid_6_delay_21_11;
  reg                 io_A_Valid_6_delay_22_10;
  reg                 io_A_Valid_6_delay_23_9;
  reg                 io_A_Valid_6_delay_24_8;
  reg                 io_A_Valid_6_delay_25_7;
  reg                 io_A_Valid_6_delay_26_6;
  reg                 io_A_Valid_6_delay_27_5;
  reg                 io_A_Valid_6_delay_28_4;
  reg                 io_A_Valid_6_delay_29_3;
  reg                 io_A_Valid_6_delay_30_2;
  reg                 io_A_Valid_6_delay_31_1;
  reg                 io_A_Valid_6_delay_32;
  reg                 io_B_Valid_32_delay_1_5;
  reg                 io_B_Valid_32_delay_2_4;
  reg                 io_B_Valid_32_delay_3_3;
  reg                 io_B_Valid_32_delay_4_2;
  reg                 io_B_Valid_32_delay_5_1;
  reg                 io_B_Valid_32_delay_6;
  reg                 io_A_Valid_6_delay_1_32;
  reg                 io_A_Valid_6_delay_2_31;
  reg                 io_A_Valid_6_delay_3_30;
  reg                 io_A_Valid_6_delay_4_29;
  reg                 io_A_Valid_6_delay_5_28;
  reg                 io_A_Valid_6_delay_6_27;
  reg                 io_A_Valid_6_delay_7_26;
  reg                 io_A_Valid_6_delay_8_25;
  reg                 io_A_Valid_6_delay_9_24;
  reg                 io_A_Valid_6_delay_10_23;
  reg                 io_A_Valid_6_delay_11_22;
  reg                 io_A_Valid_6_delay_12_21;
  reg                 io_A_Valid_6_delay_13_20;
  reg                 io_A_Valid_6_delay_14_19;
  reg                 io_A_Valid_6_delay_15_18;
  reg                 io_A_Valid_6_delay_16_17;
  reg                 io_A_Valid_6_delay_17_16;
  reg                 io_A_Valid_6_delay_18_15;
  reg                 io_A_Valid_6_delay_19_14;
  reg                 io_A_Valid_6_delay_20_13;
  reg                 io_A_Valid_6_delay_21_12;
  reg                 io_A_Valid_6_delay_22_11;
  reg                 io_A_Valid_6_delay_23_10;
  reg                 io_A_Valid_6_delay_24_9;
  reg                 io_A_Valid_6_delay_25_8;
  reg                 io_A_Valid_6_delay_26_7;
  reg                 io_A_Valid_6_delay_27_6;
  reg                 io_A_Valid_6_delay_28_5;
  reg                 io_A_Valid_6_delay_29_4;
  reg                 io_A_Valid_6_delay_30_3;
  reg                 io_A_Valid_6_delay_31_2;
  reg                 io_A_Valid_6_delay_32_1;
  reg                 io_A_Valid_6_delay_33;
  reg                 io_B_Valid_33_delay_1_5;
  reg                 io_B_Valid_33_delay_2_4;
  reg                 io_B_Valid_33_delay_3_3;
  reg                 io_B_Valid_33_delay_4_2;
  reg                 io_B_Valid_33_delay_5_1;
  reg                 io_B_Valid_33_delay_6;
  reg                 io_A_Valid_6_delay_1_33;
  reg                 io_A_Valid_6_delay_2_32;
  reg                 io_A_Valid_6_delay_3_31;
  reg                 io_A_Valid_6_delay_4_30;
  reg                 io_A_Valid_6_delay_5_29;
  reg                 io_A_Valid_6_delay_6_28;
  reg                 io_A_Valid_6_delay_7_27;
  reg                 io_A_Valid_6_delay_8_26;
  reg                 io_A_Valid_6_delay_9_25;
  reg                 io_A_Valid_6_delay_10_24;
  reg                 io_A_Valid_6_delay_11_23;
  reg                 io_A_Valid_6_delay_12_22;
  reg                 io_A_Valid_6_delay_13_21;
  reg                 io_A_Valid_6_delay_14_20;
  reg                 io_A_Valid_6_delay_15_19;
  reg                 io_A_Valid_6_delay_16_18;
  reg                 io_A_Valid_6_delay_17_17;
  reg                 io_A_Valid_6_delay_18_16;
  reg                 io_A_Valid_6_delay_19_15;
  reg                 io_A_Valid_6_delay_20_14;
  reg                 io_A_Valid_6_delay_21_13;
  reg                 io_A_Valid_6_delay_22_12;
  reg                 io_A_Valid_6_delay_23_11;
  reg                 io_A_Valid_6_delay_24_10;
  reg                 io_A_Valid_6_delay_25_9;
  reg                 io_A_Valid_6_delay_26_8;
  reg                 io_A_Valid_6_delay_27_7;
  reg                 io_A_Valid_6_delay_28_6;
  reg                 io_A_Valid_6_delay_29_5;
  reg                 io_A_Valid_6_delay_30_4;
  reg                 io_A_Valid_6_delay_31_3;
  reg                 io_A_Valid_6_delay_32_2;
  reg                 io_A_Valid_6_delay_33_1;
  reg                 io_A_Valid_6_delay_34;
  reg                 io_B_Valid_34_delay_1_5;
  reg                 io_B_Valid_34_delay_2_4;
  reg                 io_B_Valid_34_delay_3_3;
  reg                 io_B_Valid_34_delay_4_2;
  reg                 io_B_Valid_34_delay_5_1;
  reg                 io_B_Valid_34_delay_6;
  reg                 io_A_Valid_6_delay_1_34;
  reg                 io_A_Valid_6_delay_2_33;
  reg                 io_A_Valid_6_delay_3_32;
  reg                 io_A_Valid_6_delay_4_31;
  reg                 io_A_Valid_6_delay_5_30;
  reg                 io_A_Valid_6_delay_6_29;
  reg                 io_A_Valid_6_delay_7_28;
  reg                 io_A_Valid_6_delay_8_27;
  reg                 io_A_Valid_6_delay_9_26;
  reg                 io_A_Valid_6_delay_10_25;
  reg                 io_A_Valid_6_delay_11_24;
  reg                 io_A_Valid_6_delay_12_23;
  reg                 io_A_Valid_6_delay_13_22;
  reg                 io_A_Valid_6_delay_14_21;
  reg                 io_A_Valid_6_delay_15_20;
  reg                 io_A_Valid_6_delay_16_19;
  reg                 io_A_Valid_6_delay_17_18;
  reg                 io_A_Valid_6_delay_18_17;
  reg                 io_A_Valid_6_delay_19_16;
  reg                 io_A_Valid_6_delay_20_15;
  reg                 io_A_Valid_6_delay_21_14;
  reg                 io_A_Valid_6_delay_22_13;
  reg                 io_A_Valid_6_delay_23_12;
  reg                 io_A_Valid_6_delay_24_11;
  reg                 io_A_Valid_6_delay_25_10;
  reg                 io_A_Valid_6_delay_26_9;
  reg                 io_A_Valid_6_delay_27_8;
  reg                 io_A_Valid_6_delay_28_7;
  reg                 io_A_Valid_6_delay_29_6;
  reg                 io_A_Valid_6_delay_30_5;
  reg                 io_A_Valid_6_delay_31_4;
  reg                 io_A_Valid_6_delay_32_3;
  reg                 io_A_Valid_6_delay_33_2;
  reg                 io_A_Valid_6_delay_34_1;
  reg                 io_A_Valid_6_delay_35;
  reg                 io_B_Valid_35_delay_1_5;
  reg                 io_B_Valid_35_delay_2_4;
  reg                 io_B_Valid_35_delay_3_3;
  reg                 io_B_Valid_35_delay_4_2;
  reg                 io_B_Valid_35_delay_5_1;
  reg                 io_B_Valid_35_delay_6;
  reg                 io_A_Valid_6_delay_1_35;
  reg                 io_A_Valid_6_delay_2_34;
  reg                 io_A_Valid_6_delay_3_33;
  reg                 io_A_Valid_6_delay_4_32;
  reg                 io_A_Valid_6_delay_5_31;
  reg                 io_A_Valid_6_delay_6_30;
  reg                 io_A_Valid_6_delay_7_29;
  reg                 io_A_Valid_6_delay_8_28;
  reg                 io_A_Valid_6_delay_9_27;
  reg                 io_A_Valid_6_delay_10_26;
  reg                 io_A_Valid_6_delay_11_25;
  reg                 io_A_Valid_6_delay_12_24;
  reg                 io_A_Valid_6_delay_13_23;
  reg                 io_A_Valid_6_delay_14_22;
  reg                 io_A_Valid_6_delay_15_21;
  reg                 io_A_Valid_6_delay_16_20;
  reg                 io_A_Valid_6_delay_17_19;
  reg                 io_A_Valid_6_delay_18_18;
  reg                 io_A_Valid_6_delay_19_17;
  reg                 io_A_Valid_6_delay_20_16;
  reg                 io_A_Valid_6_delay_21_15;
  reg                 io_A_Valid_6_delay_22_14;
  reg                 io_A_Valid_6_delay_23_13;
  reg                 io_A_Valid_6_delay_24_12;
  reg                 io_A_Valid_6_delay_25_11;
  reg                 io_A_Valid_6_delay_26_10;
  reg                 io_A_Valid_6_delay_27_9;
  reg                 io_A_Valid_6_delay_28_8;
  reg                 io_A_Valid_6_delay_29_7;
  reg                 io_A_Valid_6_delay_30_6;
  reg                 io_A_Valid_6_delay_31_5;
  reg                 io_A_Valid_6_delay_32_4;
  reg                 io_A_Valid_6_delay_33_3;
  reg                 io_A_Valid_6_delay_34_2;
  reg                 io_A_Valid_6_delay_35_1;
  reg                 io_A_Valid_6_delay_36;
  reg                 io_B_Valid_36_delay_1_5;
  reg                 io_B_Valid_36_delay_2_4;
  reg                 io_B_Valid_36_delay_3_3;
  reg                 io_B_Valid_36_delay_4_2;
  reg                 io_B_Valid_36_delay_5_1;
  reg                 io_B_Valid_36_delay_6;
  reg                 io_A_Valid_6_delay_1_36;
  reg                 io_A_Valid_6_delay_2_35;
  reg                 io_A_Valid_6_delay_3_34;
  reg                 io_A_Valid_6_delay_4_33;
  reg                 io_A_Valid_6_delay_5_32;
  reg                 io_A_Valid_6_delay_6_31;
  reg                 io_A_Valid_6_delay_7_30;
  reg                 io_A_Valid_6_delay_8_29;
  reg                 io_A_Valid_6_delay_9_28;
  reg                 io_A_Valid_6_delay_10_27;
  reg                 io_A_Valid_6_delay_11_26;
  reg                 io_A_Valid_6_delay_12_25;
  reg                 io_A_Valid_6_delay_13_24;
  reg                 io_A_Valid_6_delay_14_23;
  reg                 io_A_Valid_6_delay_15_22;
  reg                 io_A_Valid_6_delay_16_21;
  reg                 io_A_Valid_6_delay_17_20;
  reg                 io_A_Valid_6_delay_18_19;
  reg                 io_A_Valid_6_delay_19_18;
  reg                 io_A_Valid_6_delay_20_17;
  reg                 io_A_Valid_6_delay_21_16;
  reg                 io_A_Valid_6_delay_22_15;
  reg                 io_A_Valid_6_delay_23_14;
  reg                 io_A_Valid_6_delay_24_13;
  reg                 io_A_Valid_6_delay_25_12;
  reg                 io_A_Valid_6_delay_26_11;
  reg                 io_A_Valid_6_delay_27_10;
  reg                 io_A_Valid_6_delay_28_9;
  reg                 io_A_Valid_6_delay_29_8;
  reg                 io_A_Valid_6_delay_30_7;
  reg                 io_A_Valid_6_delay_31_6;
  reg                 io_A_Valid_6_delay_32_5;
  reg                 io_A_Valid_6_delay_33_4;
  reg                 io_A_Valid_6_delay_34_3;
  reg                 io_A_Valid_6_delay_35_2;
  reg                 io_A_Valid_6_delay_36_1;
  reg                 io_A_Valid_6_delay_37;
  reg                 io_B_Valid_37_delay_1_5;
  reg                 io_B_Valid_37_delay_2_4;
  reg                 io_B_Valid_37_delay_3_3;
  reg                 io_B_Valid_37_delay_4_2;
  reg                 io_B_Valid_37_delay_5_1;
  reg                 io_B_Valid_37_delay_6;
  reg                 io_A_Valid_6_delay_1_37;
  reg                 io_A_Valid_6_delay_2_36;
  reg                 io_A_Valid_6_delay_3_35;
  reg                 io_A_Valid_6_delay_4_34;
  reg                 io_A_Valid_6_delay_5_33;
  reg                 io_A_Valid_6_delay_6_32;
  reg                 io_A_Valid_6_delay_7_31;
  reg                 io_A_Valid_6_delay_8_30;
  reg                 io_A_Valid_6_delay_9_29;
  reg                 io_A_Valid_6_delay_10_28;
  reg                 io_A_Valid_6_delay_11_27;
  reg                 io_A_Valid_6_delay_12_26;
  reg                 io_A_Valid_6_delay_13_25;
  reg                 io_A_Valid_6_delay_14_24;
  reg                 io_A_Valid_6_delay_15_23;
  reg                 io_A_Valid_6_delay_16_22;
  reg                 io_A_Valid_6_delay_17_21;
  reg                 io_A_Valid_6_delay_18_20;
  reg                 io_A_Valid_6_delay_19_19;
  reg                 io_A_Valid_6_delay_20_18;
  reg                 io_A_Valid_6_delay_21_17;
  reg                 io_A_Valid_6_delay_22_16;
  reg                 io_A_Valid_6_delay_23_15;
  reg                 io_A_Valid_6_delay_24_14;
  reg                 io_A_Valid_6_delay_25_13;
  reg                 io_A_Valid_6_delay_26_12;
  reg                 io_A_Valid_6_delay_27_11;
  reg                 io_A_Valid_6_delay_28_10;
  reg                 io_A_Valid_6_delay_29_9;
  reg                 io_A_Valid_6_delay_30_8;
  reg                 io_A_Valid_6_delay_31_7;
  reg                 io_A_Valid_6_delay_32_6;
  reg                 io_A_Valid_6_delay_33_5;
  reg                 io_A_Valid_6_delay_34_4;
  reg                 io_A_Valid_6_delay_35_3;
  reg                 io_A_Valid_6_delay_36_2;
  reg                 io_A_Valid_6_delay_37_1;
  reg                 io_A_Valid_6_delay_38;
  reg                 io_B_Valid_38_delay_1_5;
  reg                 io_B_Valid_38_delay_2_4;
  reg                 io_B_Valid_38_delay_3_3;
  reg                 io_B_Valid_38_delay_4_2;
  reg                 io_B_Valid_38_delay_5_1;
  reg                 io_B_Valid_38_delay_6;
  reg                 io_A_Valid_6_delay_1_38;
  reg                 io_A_Valid_6_delay_2_37;
  reg                 io_A_Valid_6_delay_3_36;
  reg                 io_A_Valid_6_delay_4_35;
  reg                 io_A_Valid_6_delay_5_34;
  reg                 io_A_Valid_6_delay_6_33;
  reg                 io_A_Valid_6_delay_7_32;
  reg                 io_A_Valid_6_delay_8_31;
  reg                 io_A_Valid_6_delay_9_30;
  reg                 io_A_Valid_6_delay_10_29;
  reg                 io_A_Valid_6_delay_11_28;
  reg                 io_A_Valid_6_delay_12_27;
  reg                 io_A_Valid_6_delay_13_26;
  reg                 io_A_Valid_6_delay_14_25;
  reg                 io_A_Valid_6_delay_15_24;
  reg                 io_A_Valid_6_delay_16_23;
  reg                 io_A_Valid_6_delay_17_22;
  reg                 io_A_Valid_6_delay_18_21;
  reg                 io_A_Valid_6_delay_19_20;
  reg                 io_A_Valid_6_delay_20_19;
  reg                 io_A_Valid_6_delay_21_18;
  reg                 io_A_Valid_6_delay_22_17;
  reg                 io_A_Valid_6_delay_23_16;
  reg                 io_A_Valid_6_delay_24_15;
  reg                 io_A_Valid_6_delay_25_14;
  reg                 io_A_Valid_6_delay_26_13;
  reg                 io_A_Valid_6_delay_27_12;
  reg                 io_A_Valid_6_delay_28_11;
  reg                 io_A_Valid_6_delay_29_10;
  reg                 io_A_Valid_6_delay_30_9;
  reg                 io_A_Valid_6_delay_31_8;
  reg                 io_A_Valid_6_delay_32_7;
  reg                 io_A_Valid_6_delay_33_6;
  reg                 io_A_Valid_6_delay_34_5;
  reg                 io_A_Valid_6_delay_35_4;
  reg                 io_A_Valid_6_delay_36_3;
  reg                 io_A_Valid_6_delay_37_2;
  reg                 io_A_Valid_6_delay_38_1;
  reg                 io_A_Valid_6_delay_39;
  reg                 io_B_Valid_39_delay_1_5;
  reg                 io_B_Valid_39_delay_2_4;
  reg                 io_B_Valid_39_delay_3_3;
  reg                 io_B_Valid_39_delay_4_2;
  reg                 io_B_Valid_39_delay_5_1;
  reg                 io_B_Valid_39_delay_6;
  reg                 io_A_Valid_6_delay_1_39;
  reg                 io_A_Valid_6_delay_2_38;
  reg                 io_A_Valid_6_delay_3_37;
  reg                 io_A_Valid_6_delay_4_36;
  reg                 io_A_Valid_6_delay_5_35;
  reg                 io_A_Valid_6_delay_6_34;
  reg                 io_A_Valid_6_delay_7_33;
  reg                 io_A_Valid_6_delay_8_32;
  reg                 io_A_Valid_6_delay_9_31;
  reg                 io_A_Valid_6_delay_10_30;
  reg                 io_A_Valid_6_delay_11_29;
  reg                 io_A_Valid_6_delay_12_28;
  reg                 io_A_Valid_6_delay_13_27;
  reg                 io_A_Valid_6_delay_14_26;
  reg                 io_A_Valid_6_delay_15_25;
  reg                 io_A_Valid_6_delay_16_24;
  reg                 io_A_Valid_6_delay_17_23;
  reg                 io_A_Valid_6_delay_18_22;
  reg                 io_A_Valid_6_delay_19_21;
  reg                 io_A_Valid_6_delay_20_20;
  reg                 io_A_Valid_6_delay_21_19;
  reg                 io_A_Valid_6_delay_22_18;
  reg                 io_A_Valid_6_delay_23_17;
  reg                 io_A_Valid_6_delay_24_16;
  reg                 io_A_Valid_6_delay_25_15;
  reg                 io_A_Valid_6_delay_26_14;
  reg                 io_A_Valid_6_delay_27_13;
  reg                 io_A_Valid_6_delay_28_12;
  reg                 io_A_Valid_6_delay_29_11;
  reg                 io_A_Valid_6_delay_30_10;
  reg                 io_A_Valid_6_delay_31_9;
  reg                 io_A_Valid_6_delay_32_8;
  reg                 io_A_Valid_6_delay_33_7;
  reg                 io_A_Valid_6_delay_34_6;
  reg                 io_A_Valid_6_delay_35_5;
  reg                 io_A_Valid_6_delay_36_4;
  reg                 io_A_Valid_6_delay_37_3;
  reg                 io_A_Valid_6_delay_38_2;
  reg                 io_A_Valid_6_delay_39_1;
  reg                 io_A_Valid_6_delay_40;
  reg                 io_B_Valid_40_delay_1_5;
  reg                 io_B_Valid_40_delay_2_4;
  reg                 io_B_Valid_40_delay_3_3;
  reg                 io_B_Valid_40_delay_4_2;
  reg                 io_B_Valid_40_delay_5_1;
  reg                 io_B_Valid_40_delay_6;
  reg                 io_A_Valid_6_delay_1_40;
  reg                 io_A_Valid_6_delay_2_39;
  reg                 io_A_Valid_6_delay_3_38;
  reg                 io_A_Valid_6_delay_4_37;
  reg                 io_A_Valid_6_delay_5_36;
  reg                 io_A_Valid_6_delay_6_35;
  reg                 io_A_Valid_6_delay_7_34;
  reg                 io_A_Valid_6_delay_8_33;
  reg                 io_A_Valid_6_delay_9_32;
  reg                 io_A_Valid_6_delay_10_31;
  reg                 io_A_Valid_6_delay_11_30;
  reg                 io_A_Valid_6_delay_12_29;
  reg                 io_A_Valid_6_delay_13_28;
  reg                 io_A_Valid_6_delay_14_27;
  reg                 io_A_Valid_6_delay_15_26;
  reg                 io_A_Valid_6_delay_16_25;
  reg                 io_A_Valid_6_delay_17_24;
  reg                 io_A_Valid_6_delay_18_23;
  reg                 io_A_Valid_6_delay_19_22;
  reg                 io_A_Valid_6_delay_20_21;
  reg                 io_A_Valid_6_delay_21_20;
  reg                 io_A_Valid_6_delay_22_19;
  reg                 io_A_Valid_6_delay_23_18;
  reg                 io_A_Valid_6_delay_24_17;
  reg                 io_A_Valid_6_delay_25_16;
  reg                 io_A_Valid_6_delay_26_15;
  reg                 io_A_Valid_6_delay_27_14;
  reg                 io_A_Valid_6_delay_28_13;
  reg                 io_A_Valid_6_delay_29_12;
  reg                 io_A_Valid_6_delay_30_11;
  reg                 io_A_Valid_6_delay_31_10;
  reg                 io_A_Valid_6_delay_32_9;
  reg                 io_A_Valid_6_delay_33_8;
  reg                 io_A_Valid_6_delay_34_7;
  reg                 io_A_Valid_6_delay_35_6;
  reg                 io_A_Valid_6_delay_36_5;
  reg                 io_A_Valid_6_delay_37_4;
  reg                 io_A_Valid_6_delay_38_3;
  reg                 io_A_Valid_6_delay_39_2;
  reg                 io_A_Valid_6_delay_40_1;
  reg                 io_A_Valid_6_delay_41;
  reg                 io_B_Valid_41_delay_1_5;
  reg                 io_B_Valid_41_delay_2_4;
  reg                 io_B_Valid_41_delay_3_3;
  reg                 io_B_Valid_41_delay_4_2;
  reg                 io_B_Valid_41_delay_5_1;
  reg                 io_B_Valid_41_delay_6;
  reg                 io_A_Valid_6_delay_1_41;
  reg                 io_A_Valid_6_delay_2_40;
  reg                 io_A_Valid_6_delay_3_39;
  reg                 io_A_Valid_6_delay_4_38;
  reg                 io_A_Valid_6_delay_5_37;
  reg                 io_A_Valid_6_delay_6_36;
  reg                 io_A_Valid_6_delay_7_35;
  reg                 io_A_Valid_6_delay_8_34;
  reg                 io_A_Valid_6_delay_9_33;
  reg                 io_A_Valid_6_delay_10_32;
  reg                 io_A_Valid_6_delay_11_31;
  reg                 io_A_Valid_6_delay_12_30;
  reg                 io_A_Valid_6_delay_13_29;
  reg                 io_A_Valid_6_delay_14_28;
  reg                 io_A_Valid_6_delay_15_27;
  reg                 io_A_Valid_6_delay_16_26;
  reg                 io_A_Valid_6_delay_17_25;
  reg                 io_A_Valid_6_delay_18_24;
  reg                 io_A_Valid_6_delay_19_23;
  reg                 io_A_Valid_6_delay_20_22;
  reg                 io_A_Valid_6_delay_21_21;
  reg                 io_A_Valid_6_delay_22_20;
  reg                 io_A_Valid_6_delay_23_19;
  reg                 io_A_Valid_6_delay_24_18;
  reg                 io_A_Valid_6_delay_25_17;
  reg                 io_A_Valid_6_delay_26_16;
  reg                 io_A_Valid_6_delay_27_15;
  reg                 io_A_Valid_6_delay_28_14;
  reg                 io_A_Valid_6_delay_29_13;
  reg                 io_A_Valid_6_delay_30_12;
  reg                 io_A_Valid_6_delay_31_11;
  reg                 io_A_Valid_6_delay_32_10;
  reg                 io_A_Valid_6_delay_33_9;
  reg                 io_A_Valid_6_delay_34_8;
  reg                 io_A_Valid_6_delay_35_7;
  reg                 io_A_Valid_6_delay_36_6;
  reg                 io_A_Valid_6_delay_37_5;
  reg                 io_A_Valid_6_delay_38_4;
  reg                 io_A_Valid_6_delay_39_3;
  reg                 io_A_Valid_6_delay_40_2;
  reg                 io_A_Valid_6_delay_41_1;
  reg                 io_A_Valid_6_delay_42;
  reg                 io_B_Valid_42_delay_1_5;
  reg                 io_B_Valid_42_delay_2_4;
  reg                 io_B_Valid_42_delay_3_3;
  reg                 io_B_Valid_42_delay_4_2;
  reg                 io_B_Valid_42_delay_5_1;
  reg                 io_B_Valid_42_delay_6;
  reg                 io_A_Valid_6_delay_1_42;
  reg                 io_A_Valid_6_delay_2_41;
  reg                 io_A_Valid_6_delay_3_40;
  reg                 io_A_Valid_6_delay_4_39;
  reg                 io_A_Valid_6_delay_5_38;
  reg                 io_A_Valid_6_delay_6_37;
  reg                 io_A_Valid_6_delay_7_36;
  reg                 io_A_Valid_6_delay_8_35;
  reg                 io_A_Valid_6_delay_9_34;
  reg                 io_A_Valid_6_delay_10_33;
  reg                 io_A_Valid_6_delay_11_32;
  reg                 io_A_Valid_6_delay_12_31;
  reg                 io_A_Valid_6_delay_13_30;
  reg                 io_A_Valid_6_delay_14_29;
  reg                 io_A_Valid_6_delay_15_28;
  reg                 io_A_Valid_6_delay_16_27;
  reg                 io_A_Valid_6_delay_17_26;
  reg                 io_A_Valid_6_delay_18_25;
  reg                 io_A_Valid_6_delay_19_24;
  reg                 io_A_Valid_6_delay_20_23;
  reg                 io_A_Valid_6_delay_21_22;
  reg                 io_A_Valid_6_delay_22_21;
  reg                 io_A_Valid_6_delay_23_20;
  reg                 io_A_Valid_6_delay_24_19;
  reg                 io_A_Valid_6_delay_25_18;
  reg                 io_A_Valid_6_delay_26_17;
  reg                 io_A_Valid_6_delay_27_16;
  reg                 io_A_Valid_6_delay_28_15;
  reg                 io_A_Valid_6_delay_29_14;
  reg                 io_A_Valid_6_delay_30_13;
  reg                 io_A_Valid_6_delay_31_12;
  reg                 io_A_Valid_6_delay_32_11;
  reg                 io_A_Valid_6_delay_33_10;
  reg                 io_A_Valid_6_delay_34_9;
  reg                 io_A_Valid_6_delay_35_8;
  reg                 io_A_Valid_6_delay_36_7;
  reg                 io_A_Valid_6_delay_37_6;
  reg                 io_A_Valid_6_delay_38_5;
  reg                 io_A_Valid_6_delay_39_4;
  reg                 io_A_Valid_6_delay_40_3;
  reg                 io_A_Valid_6_delay_41_2;
  reg                 io_A_Valid_6_delay_42_1;
  reg                 io_A_Valid_6_delay_43;
  reg                 io_B_Valid_43_delay_1_5;
  reg                 io_B_Valid_43_delay_2_4;
  reg                 io_B_Valid_43_delay_3_3;
  reg                 io_B_Valid_43_delay_4_2;
  reg                 io_B_Valid_43_delay_5_1;
  reg                 io_B_Valid_43_delay_6;
  reg                 io_A_Valid_6_delay_1_43;
  reg                 io_A_Valid_6_delay_2_42;
  reg                 io_A_Valid_6_delay_3_41;
  reg                 io_A_Valid_6_delay_4_40;
  reg                 io_A_Valid_6_delay_5_39;
  reg                 io_A_Valid_6_delay_6_38;
  reg                 io_A_Valid_6_delay_7_37;
  reg                 io_A_Valid_6_delay_8_36;
  reg                 io_A_Valid_6_delay_9_35;
  reg                 io_A_Valid_6_delay_10_34;
  reg                 io_A_Valid_6_delay_11_33;
  reg                 io_A_Valid_6_delay_12_32;
  reg                 io_A_Valid_6_delay_13_31;
  reg                 io_A_Valid_6_delay_14_30;
  reg                 io_A_Valid_6_delay_15_29;
  reg                 io_A_Valid_6_delay_16_28;
  reg                 io_A_Valid_6_delay_17_27;
  reg                 io_A_Valid_6_delay_18_26;
  reg                 io_A_Valid_6_delay_19_25;
  reg                 io_A_Valid_6_delay_20_24;
  reg                 io_A_Valid_6_delay_21_23;
  reg                 io_A_Valid_6_delay_22_22;
  reg                 io_A_Valid_6_delay_23_21;
  reg                 io_A_Valid_6_delay_24_20;
  reg                 io_A_Valid_6_delay_25_19;
  reg                 io_A_Valid_6_delay_26_18;
  reg                 io_A_Valid_6_delay_27_17;
  reg                 io_A_Valid_6_delay_28_16;
  reg                 io_A_Valid_6_delay_29_15;
  reg                 io_A_Valid_6_delay_30_14;
  reg                 io_A_Valid_6_delay_31_13;
  reg                 io_A_Valid_6_delay_32_12;
  reg                 io_A_Valid_6_delay_33_11;
  reg                 io_A_Valid_6_delay_34_10;
  reg                 io_A_Valid_6_delay_35_9;
  reg                 io_A_Valid_6_delay_36_8;
  reg                 io_A_Valid_6_delay_37_7;
  reg                 io_A_Valid_6_delay_38_6;
  reg                 io_A_Valid_6_delay_39_5;
  reg                 io_A_Valid_6_delay_40_4;
  reg                 io_A_Valid_6_delay_41_3;
  reg                 io_A_Valid_6_delay_42_2;
  reg                 io_A_Valid_6_delay_43_1;
  reg                 io_A_Valid_6_delay_44;
  reg                 io_B_Valid_44_delay_1_5;
  reg                 io_B_Valid_44_delay_2_4;
  reg                 io_B_Valid_44_delay_3_3;
  reg                 io_B_Valid_44_delay_4_2;
  reg                 io_B_Valid_44_delay_5_1;
  reg                 io_B_Valid_44_delay_6;
  reg                 io_A_Valid_6_delay_1_44;
  reg                 io_A_Valid_6_delay_2_43;
  reg                 io_A_Valid_6_delay_3_42;
  reg                 io_A_Valid_6_delay_4_41;
  reg                 io_A_Valid_6_delay_5_40;
  reg                 io_A_Valid_6_delay_6_39;
  reg                 io_A_Valid_6_delay_7_38;
  reg                 io_A_Valid_6_delay_8_37;
  reg                 io_A_Valid_6_delay_9_36;
  reg                 io_A_Valid_6_delay_10_35;
  reg                 io_A_Valid_6_delay_11_34;
  reg                 io_A_Valid_6_delay_12_33;
  reg                 io_A_Valid_6_delay_13_32;
  reg                 io_A_Valid_6_delay_14_31;
  reg                 io_A_Valid_6_delay_15_30;
  reg                 io_A_Valid_6_delay_16_29;
  reg                 io_A_Valid_6_delay_17_28;
  reg                 io_A_Valid_6_delay_18_27;
  reg                 io_A_Valid_6_delay_19_26;
  reg                 io_A_Valid_6_delay_20_25;
  reg                 io_A_Valid_6_delay_21_24;
  reg                 io_A_Valid_6_delay_22_23;
  reg                 io_A_Valid_6_delay_23_22;
  reg                 io_A_Valid_6_delay_24_21;
  reg                 io_A_Valid_6_delay_25_20;
  reg                 io_A_Valid_6_delay_26_19;
  reg                 io_A_Valid_6_delay_27_18;
  reg                 io_A_Valid_6_delay_28_17;
  reg                 io_A_Valid_6_delay_29_16;
  reg                 io_A_Valid_6_delay_30_15;
  reg                 io_A_Valid_6_delay_31_14;
  reg                 io_A_Valid_6_delay_32_13;
  reg                 io_A_Valid_6_delay_33_12;
  reg                 io_A_Valid_6_delay_34_11;
  reg                 io_A_Valid_6_delay_35_10;
  reg                 io_A_Valid_6_delay_36_9;
  reg                 io_A_Valid_6_delay_37_8;
  reg                 io_A_Valid_6_delay_38_7;
  reg                 io_A_Valid_6_delay_39_6;
  reg                 io_A_Valid_6_delay_40_5;
  reg                 io_A_Valid_6_delay_41_4;
  reg                 io_A_Valid_6_delay_42_3;
  reg                 io_A_Valid_6_delay_43_2;
  reg                 io_A_Valid_6_delay_44_1;
  reg                 io_A_Valid_6_delay_45;
  reg                 io_B_Valid_45_delay_1_5;
  reg                 io_B_Valid_45_delay_2_4;
  reg                 io_B_Valid_45_delay_3_3;
  reg                 io_B_Valid_45_delay_4_2;
  reg                 io_B_Valid_45_delay_5_1;
  reg                 io_B_Valid_45_delay_6;
  reg                 io_A_Valid_6_delay_1_45;
  reg                 io_A_Valid_6_delay_2_44;
  reg                 io_A_Valid_6_delay_3_43;
  reg                 io_A_Valid_6_delay_4_42;
  reg                 io_A_Valid_6_delay_5_41;
  reg                 io_A_Valid_6_delay_6_40;
  reg                 io_A_Valid_6_delay_7_39;
  reg                 io_A_Valid_6_delay_8_38;
  reg                 io_A_Valid_6_delay_9_37;
  reg                 io_A_Valid_6_delay_10_36;
  reg                 io_A_Valid_6_delay_11_35;
  reg                 io_A_Valid_6_delay_12_34;
  reg                 io_A_Valid_6_delay_13_33;
  reg                 io_A_Valid_6_delay_14_32;
  reg                 io_A_Valid_6_delay_15_31;
  reg                 io_A_Valid_6_delay_16_30;
  reg                 io_A_Valid_6_delay_17_29;
  reg                 io_A_Valid_6_delay_18_28;
  reg                 io_A_Valid_6_delay_19_27;
  reg                 io_A_Valid_6_delay_20_26;
  reg                 io_A_Valid_6_delay_21_25;
  reg                 io_A_Valid_6_delay_22_24;
  reg                 io_A_Valid_6_delay_23_23;
  reg                 io_A_Valid_6_delay_24_22;
  reg                 io_A_Valid_6_delay_25_21;
  reg                 io_A_Valid_6_delay_26_20;
  reg                 io_A_Valid_6_delay_27_19;
  reg                 io_A_Valid_6_delay_28_18;
  reg                 io_A_Valid_6_delay_29_17;
  reg                 io_A_Valid_6_delay_30_16;
  reg                 io_A_Valid_6_delay_31_15;
  reg                 io_A_Valid_6_delay_32_14;
  reg                 io_A_Valid_6_delay_33_13;
  reg                 io_A_Valid_6_delay_34_12;
  reg                 io_A_Valid_6_delay_35_11;
  reg                 io_A_Valid_6_delay_36_10;
  reg                 io_A_Valid_6_delay_37_9;
  reg                 io_A_Valid_6_delay_38_8;
  reg                 io_A_Valid_6_delay_39_7;
  reg                 io_A_Valid_6_delay_40_6;
  reg                 io_A_Valid_6_delay_41_5;
  reg                 io_A_Valid_6_delay_42_4;
  reg                 io_A_Valid_6_delay_43_3;
  reg                 io_A_Valid_6_delay_44_2;
  reg                 io_A_Valid_6_delay_45_1;
  reg                 io_A_Valid_6_delay_46;
  reg                 io_B_Valid_46_delay_1_5;
  reg                 io_B_Valid_46_delay_2_4;
  reg                 io_B_Valid_46_delay_3_3;
  reg                 io_B_Valid_46_delay_4_2;
  reg                 io_B_Valid_46_delay_5_1;
  reg                 io_B_Valid_46_delay_6;
  reg                 io_A_Valid_6_delay_1_46;
  reg                 io_A_Valid_6_delay_2_45;
  reg                 io_A_Valid_6_delay_3_44;
  reg                 io_A_Valid_6_delay_4_43;
  reg                 io_A_Valid_6_delay_5_42;
  reg                 io_A_Valid_6_delay_6_41;
  reg                 io_A_Valid_6_delay_7_40;
  reg                 io_A_Valid_6_delay_8_39;
  reg                 io_A_Valid_6_delay_9_38;
  reg                 io_A_Valid_6_delay_10_37;
  reg                 io_A_Valid_6_delay_11_36;
  reg                 io_A_Valid_6_delay_12_35;
  reg                 io_A_Valid_6_delay_13_34;
  reg                 io_A_Valid_6_delay_14_33;
  reg                 io_A_Valid_6_delay_15_32;
  reg                 io_A_Valid_6_delay_16_31;
  reg                 io_A_Valid_6_delay_17_30;
  reg                 io_A_Valid_6_delay_18_29;
  reg                 io_A_Valid_6_delay_19_28;
  reg                 io_A_Valid_6_delay_20_27;
  reg                 io_A_Valid_6_delay_21_26;
  reg                 io_A_Valid_6_delay_22_25;
  reg                 io_A_Valid_6_delay_23_24;
  reg                 io_A_Valid_6_delay_24_23;
  reg                 io_A_Valid_6_delay_25_22;
  reg                 io_A_Valid_6_delay_26_21;
  reg                 io_A_Valid_6_delay_27_20;
  reg                 io_A_Valid_6_delay_28_19;
  reg                 io_A_Valid_6_delay_29_18;
  reg                 io_A_Valid_6_delay_30_17;
  reg                 io_A_Valid_6_delay_31_16;
  reg                 io_A_Valid_6_delay_32_15;
  reg                 io_A_Valid_6_delay_33_14;
  reg                 io_A_Valid_6_delay_34_13;
  reg                 io_A_Valid_6_delay_35_12;
  reg                 io_A_Valid_6_delay_36_11;
  reg                 io_A_Valid_6_delay_37_10;
  reg                 io_A_Valid_6_delay_38_9;
  reg                 io_A_Valid_6_delay_39_8;
  reg                 io_A_Valid_6_delay_40_7;
  reg                 io_A_Valid_6_delay_41_6;
  reg                 io_A_Valid_6_delay_42_5;
  reg                 io_A_Valid_6_delay_43_4;
  reg                 io_A_Valid_6_delay_44_3;
  reg                 io_A_Valid_6_delay_45_2;
  reg                 io_A_Valid_6_delay_46_1;
  reg                 io_A_Valid_6_delay_47;
  reg                 io_B_Valid_47_delay_1_5;
  reg                 io_B_Valid_47_delay_2_4;
  reg                 io_B_Valid_47_delay_3_3;
  reg                 io_B_Valid_47_delay_4_2;
  reg                 io_B_Valid_47_delay_5_1;
  reg                 io_B_Valid_47_delay_6;
  reg                 io_A_Valid_6_delay_1_47;
  reg                 io_A_Valid_6_delay_2_46;
  reg                 io_A_Valid_6_delay_3_45;
  reg                 io_A_Valid_6_delay_4_44;
  reg                 io_A_Valid_6_delay_5_43;
  reg                 io_A_Valid_6_delay_6_42;
  reg                 io_A_Valid_6_delay_7_41;
  reg                 io_A_Valid_6_delay_8_40;
  reg                 io_A_Valid_6_delay_9_39;
  reg                 io_A_Valid_6_delay_10_38;
  reg                 io_A_Valid_6_delay_11_37;
  reg                 io_A_Valid_6_delay_12_36;
  reg                 io_A_Valid_6_delay_13_35;
  reg                 io_A_Valid_6_delay_14_34;
  reg                 io_A_Valid_6_delay_15_33;
  reg                 io_A_Valid_6_delay_16_32;
  reg                 io_A_Valid_6_delay_17_31;
  reg                 io_A_Valid_6_delay_18_30;
  reg                 io_A_Valid_6_delay_19_29;
  reg                 io_A_Valid_6_delay_20_28;
  reg                 io_A_Valid_6_delay_21_27;
  reg                 io_A_Valid_6_delay_22_26;
  reg                 io_A_Valid_6_delay_23_25;
  reg                 io_A_Valid_6_delay_24_24;
  reg                 io_A_Valid_6_delay_25_23;
  reg                 io_A_Valid_6_delay_26_22;
  reg                 io_A_Valid_6_delay_27_21;
  reg                 io_A_Valid_6_delay_28_20;
  reg                 io_A_Valid_6_delay_29_19;
  reg                 io_A_Valid_6_delay_30_18;
  reg                 io_A_Valid_6_delay_31_17;
  reg                 io_A_Valid_6_delay_32_16;
  reg                 io_A_Valid_6_delay_33_15;
  reg                 io_A_Valid_6_delay_34_14;
  reg                 io_A_Valid_6_delay_35_13;
  reg                 io_A_Valid_6_delay_36_12;
  reg                 io_A_Valid_6_delay_37_11;
  reg                 io_A_Valid_6_delay_38_10;
  reg                 io_A_Valid_6_delay_39_9;
  reg                 io_A_Valid_6_delay_40_8;
  reg                 io_A_Valid_6_delay_41_7;
  reg                 io_A_Valid_6_delay_42_6;
  reg                 io_A_Valid_6_delay_43_5;
  reg                 io_A_Valid_6_delay_44_4;
  reg                 io_A_Valid_6_delay_45_3;
  reg                 io_A_Valid_6_delay_46_2;
  reg                 io_A_Valid_6_delay_47_1;
  reg                 io_A_Valid_6_delay_48;
  reg                 io_B_Valid_48_delay_1_5;
  reg                 io_B_Valid_48_delay_2_4;
  reg                 io_B_Valid_48_delay_3_3;
  reg                 io_B_Valid_48_delay_4_2;
  reg                 io_B_Valid_48_delay_5_1;
  reg                 io_B_Valid_48_delay_6;
  reg                 io_A_Valid_6_delay_1_48;
  reg                 io_A_Valid_6_delay_2_47;
  reg                 io_A_Valid_6_delay_3_46;
  reg                 io_A_Valid_6_delay_4_45;
  reg                 io_A_Valid_6_delay_5_44;
  reg                 io_A_Valid_6_delay_6_43;
  reg                 io_A_Valid_6_delay_7_42;
  reg                 io_A_Valid_6_delay_8_41;
  reg                 io_A_Valid_6_delay_9_40;
  reg                 io_A_Valid_6_delay_10_39;
  reg                 io_A_Valid_6_delay_11_38;
  reg                 io_A_Valid_6_delay_12_37;
  reg                 io_A_Valid_6_delay_13_36;
  reg                 io_A_Valid_6_delay_14_35;
  reg                 io_A_Valid_6_delay_15_34;
  reg                 io_A_Valid_6_delay_16_33;
  reg                 io_A_Valid_6_delay_17_32;
  reg                 io_A_Valid_6_delay_18_31;
  reg                 io_A_Valid_6_delay_19_30;
  reg                 io_A_Valid_6_delay_20_29;
  reg                 io_A_Valid_6_delay_21_28;
  reg                 io_A_Valid_6_delay_22_27;
  reg                 io_A_Valid_6_delay_23_26;
  reg                 io_A_Valid_6_delay_24_25;
  reg                 io_A_Valid_6_delay_25_24;
  reg                 io_A_Valid_6_delay_26_23;
  reg                 io_A_Valid_6_delay_27_22;
  reg                 io_A_Valid_6_delay_28_21;
  reg                 io_A_Valid_6_delay_29_20;
  reg                 io_A_Valid_6_delay_30_19;
  reg                 io_A_Valid_6_delay_31_18;
  reg                 io_A_Valid_6_delay_32_17;
  reg                 io_A_Valid_6_delay_33_16;
  reg                 io_A_Valid_6_delay_34_15;
  reg                 io_A_Valid_6_delay_35_14;
  reg                 io_A_Valid_6_delay_36_13;
  reg                 io_A_Valid_6_delay_37_12;
  reg                 io_A_Valid_6_delay_38_11;
  reg                 io_A_Valid_6_delay_39_10;
  reg                 io_A_Valid_6_delay_40_9;
  reg                 io_A_Valid_6_delay_41_8;
  reg                 io_A_Valid_6_delay_42_7;
  reg                 io_A_Valid_6_delay_43_6;
  reg                 io_A_Valid_6_delay_44_5;
  reg                 io_A_Valid_6_delay_45_4;
  reg                 io_A_Valid_6_delay_46_3;
  reg                 io_A_Valid_6_delay_47_2;
  reg                 io_A_Valid_6_delay_48_1;
  reg                 io_A_Valid_6_delay_49;
  reg                 io_B_Valid_49_delay_1_5;
  reg                 io_B_Valid_49_delay_2_4;
  reg                 io_B_Valid_49_delay_3_3;
  reg                 io_B_Valid_49_delay_4_2;
  reg                 io_B_Valid_49_delay_5_1;
  reg                 io_B_Valid_49_delay_6;
  reg                 io_A_Valid_6_delay_1_49;
  reg                 io_A_Valid_6_delay_2_48;
  reg                 io_A_Valid_6_delay_3_47;
  reg                 io_A_Valid_6_delay_4_46;
  reg                 io_A_Valid_6_delay_5_45;
  reg                 io_A_Valid_6_delay_6_44;
  reg                 io_A_Valid_6_delay_7_43;
  reg                 io_A_Valid_6_delay_8_42;
  reg                 io_A_Valid_6_delay_9_41;
  reg                 io_A_Valid_6_delay_10_40;
  reg                 io_A_Valid_6_delay_11_39;
  reg                 io_A_Valid_6_delay_12_38;
  reg                 io_A_Valid_6_delay_13_37;
  reg                 io_A_Valid_6_delay_14_36;
  reg                 io_A_Valid_6_delay_15_35;
  reg                 io_A_Valid_6_delay_16_34;
  reg                 io_A_Valid_6_delay_17_33;
  reg                 io_A_Valid_6_delay_18_32;
  reg                 io_A_Valid_6_delay_19_31;
  reg                 io_A_Valid_6_delay_20_30;
  reg                 io_A_Valid_6_delay_21_29;
  reg                 io_A_Valid_6_delay_22_28;
  reg                 io_A_Valid_6_delay_23_27;
  reg                 io_A_Valid_6_delay_24_26;
  reg                 io_A_Valid_6_delay_25_25;
  reg                 io_A_Valid_6_delay_26_24;
  reg                 io_A_Valid_6_delay_27_23;
  reg                 io_A_Valid_6_delay_28_22;
  reg                 io_A_Valid_6_delay_29_21;
  reg                 io_A_Valid_6_delay_30_20;
  reg                 io_A_Valid_6_delay_31_19;
  reg                 io_A_Valid_6_delay_32_18;
  reg                 io_A_Valid_6_delay_33_17;
  reg                 io_A_Valid_6_delay_34_16;
  reg                 io_A_Valid_6_delay_35_15;
  reg                 io_A_Valid_6_delay_36_14;
  reg                 io_A_Valid_6_delay_37_13;
  reg                 io_A_Valid_6_delay_38_12;
  reg                 io_A_Valid_6_delay_39_11;
  reg                 io_A_Valid_6_delay_40_10;
  reg                 io_A_Valid_6_delay_41_9;
  reg                 io_A_Valid_6_delay_42_8;
  reg                 io_A_Valid_6_delay_43_7;
  reg                 io_A_Valid_6_delay_44_6;
  reg                 io_A_Valid_6_delay_45_5;
  reg                 io_A_Valid_6_delay_46_4;
  reg                 io_A_Valid_6_delay_47_3;
  reg                 io_A_Valid_6_delay_48_2;
  reg                 io_A_Valid_6_delay_49_1;
  reg                 io_A_Valid_6_delay_50;
  reg                 io_B_Valid_50_delay_1_5;
  reg                 io_B_Valid_50_delay_2_4;
  reg                 io_B_Valid_50_delay_3_3;
  reg                 io_B_Valid_50_delay_4_2;
  reg                 io_B_Valid_50_delay_5_1;
  reg                 io_B_Valid_50_delay_6;
  reg                 io_A_Valid_6_delay_1_50;
  reg                 io_A_Valid_6_delay_2_49;
  reg                 io_A_Valid_6_delay_3_48;
  reg                 io_A_Valid_6_delay_4_47;
  reg                 io_A_Valid_6_delay_5_46;
  reg                 io_A_Valid_6_delay_6_45;
  reg                 io_A_Valid_6_delay_7_44;
  reg                 io_A_Valid_6_delay_8_43;
  reg                 io_A_Valid_6_delay_9_42;
  reg                 io_A_Valid_6_delay_10_41;
  reg                 io_A_Valid_6_delay_11_40;
  reg                 io_A_Valid_6_delay_12_39;
  reg                 io_A_Valid_6_delay_13_38;
  reg                 io_A_Valid_6_delay_14_37;
  reg                 io_A_Valid_6_delay_15_36;
  reg                 io_A_Valid_6_delay_16_35;
  reg                 io_A_Valid_6_delay_17_34;
  reg                 io_A_Valid_6_delay_18_33;
  reg                 io_A_Valid_6_delay_19_32;
  reg                 io_A_Valid_6_delay_20_31;
  reg                 io_A_Valid_6_delay_21_30;
  reg                 io_A_Valid_6_delay_22_29;
  reg                 io_A_Valid_6_delay_23_28;
  reg                 io_A_Valid_6_delay_24_27;
  reg                 io_A_Valid_6_delay_25_26;
  reg                 io_A_Valid_6_delay_26_25;
  reg                 io_A_Valid_6_delay_27_24;
  reg                 io_A_Valid_6_delay_28_23;
  reg                 io_A_Valid_6_delay_29_22;
  reg                 io_A_Valid_6_delay_30_21;
  reg                 io_A_Valid_6_delay_31_20;
  reg                 io_A_Valid_6_delay_32_19;
  reg                 io_A_Valid_6_delay_33_18;
  reg                 io_A_Valid_6_delay_34_17;
  reg                 io_A_Valid_6_delay_35_16;
  reg                 io_A_Valid_6_delay_36_15;
  reg                 io_A_Valid_6_delay_37_14;
  reg                 io_A_Valid_6_delay_38_13;
  reg                 io_A_Valid_6_delay_39_12;
  reg                 io_A_Valid_6_delay_40_11;
  reg                 io_A_Valid_6_delay_41_10;
  reg                 io_A_Valid_6_delay_42_9;
  reg                 io_A_Valid_6_delay_43_8;
  reg                 io_A_Valid_6_delay_44_7;
  reg                 io_A_Valid_6_delay_45_6;
  reg                 io_A_Valid_6_delay_46_5;
  reg                 io_A_Valid_6_delay_47_4;
  reg                 io_A_Valid_6_delay_48_3;
  reg                 io_A_Valid_6_delay_49_2;
  reg                 io_A_Valid_6_delay_50_1;
  reg                 io_A_Valid_6_delay_51;
  reg                 io_B_Valid_51_delay_1_5;
  reg                 io_B_Valid_51_delay_2_4;
  reg                 io_B_Valid_51_delay_3_3;
  reg                 io_B_Valid_51_delay_4_2;
  reg                 io_B_Valid_51_delay_5_1;
  reg                 io_B_Valid_51_delay_6;
  reg                 io_A_Valid_6_delay_1_51;
  reg                 io_A_Valid_6_delay_2_50;
  reg                 io_A_Valid_6_delay_3_49;
  reg                 io_A_Valid_6_delay_4_48;
  reg                 io_A_Valid_6_delay_5_47;
  reg                 io_A_Valid_6_delay_6_46;
  reg                 io_A_Valid_6_delay_7_45;
  reg                 io_A_Valid_6_delay_8_44;
  reg                 io_A_Valid_6_delay_9_43;
  reg                 io_A_Valid_6_delay_10_42;
  reg                 io_A_Valid_6_delay_11_41;
  reg                 io_A_Valid_6_delay_12_40;
  reg                 io_A_Valid_6_delay_13_39;
  reg                 io_A_Valid_6_delay_14_38;
  reg                 io_A_Valid_6_delay_15_37;
  reg                 io_A_Valid_6_delay_16_36;
  reg                 io_A_Valid_6_delay_17_35;
  reg                 io_A_Valid_6_delay_18_34;
  reg                 io_A_Valid_6_delay_19_33;
  reg                 io_A_Valid_6_delay_20_32;
  reg                 io_A_Valid_6_delay_21_31;
  reg                 io_A_Valid_6_delay_22_30;
  reg                 io_A_Valid_6_delay_23_29;
  reg                 io_A_Valid_6_delay_24_28;
  reg                 io_A_Valid_6_delay_25_27;
  reg                 io_A_Valid_6_delay_26_26;
  reg                 io_A_Valid_6_delay_27_25;
  reg                 io_A_Valid_6_delay_28_24;
  reg                 io_A_Valid_6_delay_29_23;
  reg                 io_A_Valid_6_delay_30_22;
  reg                 io_A_Valid_6_delay_31_21;
  reg                 io_A_Valid_6_delay_32_20;
  reg                 io_A_Valid_6_delay_33_19;
  reg                 io_A_Valid_6_delay_34_18;
  reg                 io_A_Valid_6_delay_35_17;
  reg                 io_A_Valid_6_delay_36_16;
  reg                 io_A_Valid_6_delay_37_15;
  reg                 io_A_Valid_6_delay_38_14;
  reg                 io_A_Valid_6_delay_39_13;
  reg                 io_A_Valid_6_delay_40_12;
  reg                 io_A_Valid_6_delay_41_11;
  reg                 io_A_Valid_6_delay_42_10;
  reg                 io_A_Valid_6_delay_43_9;
  reg                 io_A_Valid_6_delay_44_8;
  reg                 io_A_Valid_6_delay_45_7;
  reg                 io_A_Valid_6_delay_46_6;
  reg                 io_A_Valid_6_delay_47_5;
  reg                 io_A_Valid_6_delay_48_4;
  reg                 io_A_Valid_6_delay_49_3;
  reg                 io_A_Valid_6_delay_50_2;
  reg                 io_A_Valid_6_delay_51_1;
  reg                 io_A_Valid_6_delay_52;
  reg                 io_B_Valid_52_delay_1_5;
  reg                 io_B_Valid_52_delay_2_4;
  reg                 io_B_Valid_52_delay_3_3;
  reg                 io_B_Valid_52_delay_4_2;
  reg                 io_B_Valid_52_delay_5_1;
  reg                 io_B_Valid_52_delay_6;
  reg                 io_A_Valid_6_delay_1_52;
  reg                 io_A_Valid_6_delay_2_51;
  reg                 io_A_Valid_6_delay_3_50;
  reg                 io_A_Valid_6_delay_4_49;
  reg                 io_A_Valid_6_delay_5_48;
  reg                 io_A_Valid_6_delay_6_47;
  reg                 io_A_Valid_6_delay_7_46;
  reg                 io_A_Valid_6_delay_8_45;
  reg                 io_A_Valid_6_delay_9_44;
  reg                 io_A_Valid_6_delay_10_43;
  reg                 io_A_Valid_6_delay_11_42;
  reg                 io_A_Valid_6_delay_12_41;
  reg                 io_A_Valid_6_delay_13_40;
  reg                 io_A_Valid_6_delay_14_39;
  reg                 io_A_Valid_6_delay_15_38;
  reg                 io_A_Valid_6_delay_16_37;
  reg                 io_A_Valid_6_delay_17_36;
  reg                 io_A_Valid_6_delay_18_35;
  reg                 io_A_Valid_6_delay_19_34;
  reg                 io_A_Valid_6_delay_20_33;
  reg                 io_A_Valid_6_delay_21_32;
  reg                 io_A_Valid_6_delay_22_31;
  reg                 io_A_Valid_6_delay_23_30;
  reg                 io_A_Valid_6_delay_24_29;
  reg                 io_A_Valid_6_delay_25_28;
  reg                 io_A_Valid_6_delay_26_27;
  reg                 io_A_Valid_6_delay_27_26;
  reg                 io_A_Valid_6_delay_28_25;
  reg                 io_A_Valid_6_delay_29_24;
  reg                 io_A_Valid_6_delay_30_23;
  reg                 io_A_Valid_6_delay_31_22;
  reg                 io_A_Valid_6_delay_32_21;
  reg                 io_A_Valid_6_delay_33_20;
  reg                 io_A_Valid_6_delay_34_19;
  reg                 io_A_Valid_6_delay_35_18;
  reg                 io_A_Valid_6_delay_36_17;
  reg                 io_A_Valid_6_delay_37_16;
  reg                 io_A_Valid_6_delay_38_15;
  reg                 io_A_Valid_6_delay_39_14;
  reg                 io_A_Valid_6_delay_40_13;
  reg                 io_A_Valid_6_delay_41_12;
  reg                 io_A_Valid_6_delay_42_11;
  reg                 io_A_Valid_6_delay_43_10;
  reg                 io_A_Valid_6_delay_44_9;
  reg                 io_A_Valid_6_delay_45_8;
  reg                 io_A_Valid_6_delay_46_7;
  reg                 io_A_Valid_6_delay_47_6;
  reg                 io_A_Valid_6_delay_48_5;
  reg                 io_A_Valid_6_delay_49_4;
  reg                 io_A_Valid_6_delay_50_3;
  reg                 io_A_Valid_6_delay_51_2;
  reg                 io_A_Valid_6_delay_52_1;
  reg                 io_A_Valid_6_delay_53;
  reg                 io_B_Valid_53_delay_1_5;
  reg                 io_B_Valid_53_delay_2_4;
  reg                 io_B_Valid_53_delay_3_3;
  reg                 io_B_Valid_53_delay_4_2;
  reg                 io_B_Valid_53_delay_5_1;
  reg                 io_B_Valid_53_delay_6;
  reg                 io_A_Valid_6_delay_1_53;
  reg                 io_A_Valid_6_delay_2_52;
  reg                 io_A_Valid_6_delay_3_51;
  reg                 io_A_Valid_6_delay_4_50;
  reg                 io_A_Valid_6_delay_5_49;
  reg                 io_A_Valid_6_delay_6_48;
  reg                 io_A_Valid_6_delay_7_47;
  reg                 io_A_Valid_6_delay_8_46;
  reg                 io_A_Valid_6_delay_9_45;
  reg                 io_A_Valid_6_delay_10_44;
  reg                 io_A_Valid_6_delay_11_43;
  reg                 io_A_Valid_6_delay_12_42;
  reg                 io_A_Valid_6_delay_13_41;
  reg                 io_A_Valid_6_delay_14_40;
  reg                 io_A_Valid_6_delay_15_39;
  reg                 io_A_Valid_6_delay_16_38;
  reg                 io_A_Valid_6_delay_17_37;
  reg                 io_A_Valid_6_delay_18_36;
  reg                 io_A_Valid_6_delay_19_35;
  reg                 io_A_Valid_6_delay_20_34;
  reg                 io_A_Valid_6_delay_21_33;
  reg                 io_A_Valid_6_delay_22_32;
  reg                 io_A_Valid_6_delay_23_31;
  reg                 io_A_Valid_6_delay_24_30;
  reg                 io_A_Valid_6_delay_25_29;
  reg                 io_A_Valid_6_delay_26_28;
  reg                 io_A_Valid_6_delay_27_27;
  reg                 io_A_Valid_6_delay_28_26;
  reg                 io_A_Valid_6_delay_29_25;
  reg                 io_A_Valid_6_delay_30_24;
  reg                 io_A_Valid_6_delay_31_23;
  reg                 io_A_Valid_6_delay_32_22;
  reg                 io_A_Valid_6_delay_33_21;
  reg                 io_A_Valid_6_delay_34_20;
  reg                 io_A_Valid_6_delay_35_19;
  reg                 io_A_Valid_6_delay_36_18;
  reg                 io_A_Valid_6_delay_37_17;
  reg                 io_A_Valid_6_delay_38_16;
  reg                 io_A_Valid_6_delay_39_15;
  reg                 io_A_Valid_6_delay_40_14;
  reg                 io_A_Valid_6_delay_41_13;
  reg                 io_A_Valid_6_delay_42_12;
  reg                 io_A_Valid_6_delay_43_11;
  reg                 io_A_Valid_6_delay_44_10;
  reg                 io_A_Valid_6_delay_45_9;
  reg                 io_A_Valid_6_delay_46_8;
  reg                 io_A_Valid_6_delay_47_7;
  reg                 io_A_Valid_6_delay_48_6;
  reg                 io_A_Valid_6_delay_49_5;
  reg                 io_A_Valid_6_delay_50_4;
  reg                 io_A_Valid_6_delay_51_3;
  reg                 io_A_Valid_6_delay_52_2;
  reg                 io_A_Valid_6_delay_53_1;
  reg                 io_A_Valid_6_delay_54;
  reg                 io_B_Valid_54_delay_1_5;
  reg                 io_B_Valid_54_delay_2_4;
  reg                 io_B_Valid_54_delay_3_3;
  reg                 io_B_Valid_54_delay_4_2;
  reg                 io_B_Valid_54_delay_5_1;
  reg                 io_B_Valid_54_delay_6;
  reg                 io_A_Valid_6_delay_1_54;
  reg                 io_A_Valid_6_delay_2_53;
  reg                 io_A_Valid_6_delay_3_52;
  reg                 io_A_Valid_6_delay_4_51;
  reg                 io_A_Valid_6_delay_5_50;
  reg                 io_A_Valid_6_delay_6_49;
  reg                 io_A_Valid_6_delay_7_48;
  reg                 io_A_Valid_6_delay_8_47;
  reg                 io_A_Valid_6_delay_9_46;
  reg                 io_A_Valid_6_delay_10_45;
  reg                 io_A_Valid_6_delay_11_44;
  reg                 io_A_Valid_6_delay_12_43;
  reg                 io_A_Valid_6_delay_13_42;
  reg                 io_A_Valid_6_delay_14_41;
  reg                 io_A_Valid_6_delay_15_40;
  reg                 io_A_Valid_6_delay_16_39;
  reg                 io_A_Valid_6_delay_17_38;
  reg                 io_A_Valid_6_delay_18_37;
  reg                 io_A_Valid_6_delay_19_36;
  reg                 io_A_Valid_6_delay_20_35;
  reg                 io_A_Valid_6_delay_21_34;
  reg                 io_A_Valid_6_delay_22_33;
  reg                 io_A_Valid_6_delay_23_32;
  reg                 io_A_Valid_6_delay_24_31;
  reg                 io_A_Valid_6_delay_25_30;
  reg                 io_A_Valid_6_delay_26_29;
  reg                 io_A_Valid_6_delay_27_28;
  reg                 io_A_Valid_6_delay_28_27;
  reg                 io_A_Valid_6_delay_29_26;
  reg                 io_A_Valid_6_delay_30_25;
  reg                 io_A_Valid_6_delay_31_24;
  reg                 io_A_Valid_6_delay_32_23;
  reg                 io_A_Valid_6_delay_33_22;
  reg                 io_A_Valid_6_delay_34_21;
  reg                 io_A_Valid_6_delay_35_20;
  reg                 io_A_Valid_6_delay_36_19;
  reg                 io_A_Valid_6_delay_37_18;
  reg                 io_A_Valid_6_delay_38_17;
  reg                 io_A_Valid_6_delay_39_16;
  reg                 io_A_Valid_6_delay_40_15;
  reg                 io_A_Valid_6_delay_41_14;
  reg                 io_A_Valid_6_delay_42_13;
  reg                 io_A_Valid_6_delay_43_12;
  reg                 io_A_Valid_6_delay_44_11;
  reg                 io_A_Valid_6_delay_45_10;
  reg                 io_A_Valid_6_delay_46_9;
  reg                 io_A_Valid_6_delay_47_8;
  reg                 io_A_Valid_6_delay_48_7;
  reg                 io_A_Valid_6_delay_49_6;
  reg                 io_A_Valid_6_delay_50_5;
  reg                 io_A_Valid_6_delay_51_4;
  reg                 io_A_Valid_6_delay_52_3;
  reg                 io_A_Valid_6_delay_53_2;
  reg                 io_A_Valid_6_delay_54_1;
  reg                 io_A_Valid_6_delay_55;
  reg                 io_B_Valid_55_delay_1_5;
  reg                 io_B_Valid_55_delay_2_4;
  reg                 io_B_Valid_55_delay_3_3;
  reg                 io_B_Valid_55_delay_4_2;
  reg                 io_B_Valid_55_delay_5_1;
  reg                 io_B_Valid_55_delay_6;
  reg                 io_A_Valid_6_delay_1_55;
  reg                 io_A_Valid_6_delay_2_54;
  reg                 io_A_Valid_6_delay_3_53;
  reg                 io_A_Valid_6_delay_4_52;
  reg                 io_A_Valid_6_delay_5_51;
  reg                 io_A_Valid_6_delay_6_50;
  reg                 io_A_Valid_6_delay_7_49;
  reg                 io_A_Valid_6_delay_8_48;
  reg                 io_A_Valid_6_delay_9_47;
  reg                 io_A_Valid_6_delay_10_46;
  reg                 io_A_Valid_6_delay_11_45;
  reg                 io_A_Valid_6_delay_12_44;
  reg                 io_A_Valid_6_delay_13_43;
  reg                 io_A_Valid_6_delay_14_42;
  reg                 io_A_Valid_6_delay_15_41;
  reg                 io_A_Valid_6_delay_16_40;
  reg                 io_A_Valid_6_delay_17_39;
  reg                 io_A_Valid_6_delay_18_38;
  reg                 io_A_Valid_6_delay_19_37;
  reg                 io_A_Valid_6_delay_20_36;
  reg                 io_A_Valid_6_delay_21_35;
  reg                 io_A_Valid_6_delay_22_34;
  reg                 io_A_Valid_6_delay_23_33;
  reg                 io_A_Valid_6_delay_24_32;
  reg                 io_A_Valid_6_delay_25_31;
  reg                 io_A_Valid_6_delay_26_30;
  reg                 io_A_Valid_6_delay_27_29;
  reg                 io_A_Valid_6_delay_28_28;
  reg                 io_A_Valid_6_delay_29_27;
  reg                 io_A_Valid_6_delay_30_26;
  reg                 io_A_Valid_6_delay_31_25;
  reg                 io_A_Valid_6_delay_32_24;
  reg                 io_A_Valid_6_delay_33_23;
  reg                 io_A_Valid_6_delay_34_22;
  reg                 io_A_Valid_6_delay_35_21;
  reg                 io_A_Valid_6_delay_36_20;
  reg                 io_A_Valid_6_delay_37_19;
  reg                 io_A_Valid_6_delay_38_18;
  reg                 io_A_Valid_6_delay_39_17;
  reg                 io_A_Valid_6_delay_40_16;
  reg                 io_A_Valid_6_delay_41_15;
  reg                 io_A_Valid_6_delay_42_14;
  reg                 io_A_Valid_6_delay_43_13;
  reg                 io_A_Valid_6_delay_44_12;
  reg                 io_A_Valid_6_delay_45_11;
  reg                 io_A_Valid_6_delay_46_10;
  reg                 io_A_Valid_6_delay_47_9;
  reg                 io_A_Valid_6_delay_48_8;
  reg                 io_A_Valid_6_delay_49_7;
  reg                 io_A_Valid_6_delay_50_6;
  reg                 io_A_Valid_6_delay_51_5;
  reg                 io_A_Valid_6_delay_52_4;
  reg                 io_A_Valid_6_delay_53_3;
  reg                 io_A_Valid_6_delay_54_2;
  reg                 io_A_Valid_6_delay_55_1;
  reg                 io_A_Valid_6_delay_56;
  reg                 io_B_Valid_56_delay_1_5;
  reg                 io_B_Valid_56_delay_2_4;
  reg                 io_B_Valid_56_delay_3_3;
  reg                 io_B_Valid_56_delay_4_2;
  reg                 io_B_Valid_56_delay_5_1;
  reg                 io_B_Valid_56_delay_6;
  reg                 io_A_Valid_6_delay_1_56;
  reg                 io_A_Valid_6_delay_2_55;
  reg                 io_A_Valid_6_delay_3_54;
  reg                 io_A_Valid_6_delay_4_53;
  reg                 io_A_Valid_6_delay_5_52;
  reg                 io_A_Valid_6_delay_6_51;
  reg                 io_A_Valid_6_delay_7_50;
  reg                 io_A_Valid_6_delay_8_49;
  reg                 io_A_Valid_6_delay_9_48;
  reg                 io_A_Valid_6_delay_10_47;
  reg                 io_A_Valid_6_delay_11_46;
  reg                 io_A_Valid_6_delay_12_45;
  reg                 io_A_Valid_6_delay_13_44;
  reg                 io_A_Valid_6_delay_14_43;
  reg                 io_A_Valid_6_delay_15_42;
  reg                 io_A_Valid_6_delay_16_41;
  reg                 io_A_Valid_6_delay_17_40;
  reg                 io_A_Valid_6_delay_18_39;
  reg                 io_A_Valid_6_delay_19_38;
  reg                 io_A_Valid_6_delay_20_37;
  reg                 io_A_Valid_6_delay_21_36;
  reg                 io_A_Valid_6_delay_22_35;
  reg                 io_A_Valid_6_delay_23_34;
  reg                 io_A_Valid_6_delay_24_33;
  reg                 io_A_Valid_6_delay_25_32;
  reg                 io_A_Valid_6_delay_26_31;
  reg                 io_A_Valid_6_delay_27_30;
  reg                 io_A_Valid_6_delay_28_29;
  reg                 io_A_Valid_6_delay_29_28;
  reg                 io_A_Valid_6_delay_30_27;
  reg                 io_A_Valid_6_delay_31_26;
  reg                 io_A_Valid_6_delay_32_25;
  reg                 io_A_Valid_6_delay_33_24;
  reg                 io_A_Valid_6_delay_34_23;
  reg                 io_A_Valid_6_delay_35_22;
  reg                 io_A_Valid_6_delay_36_21;
  reg                 io_A_Valid_6_delay_37_20;
  reg                 io_A_Valid_6_delay_38_19;
  reg                 io_A_Valid_6_delay_39_18;
  reg                 io_A_Valid_6_delay_40_17;
  reg                 io_A_Valid_6_delay_41_16;
  reg                 io_A_Valid_6_delay_42_15;
  reg                 io_A_Valid_6_delay_43_14;
  reg                 io_A_Valid_6_delay_44_13;
  reg                 io_A_Valid_6_delay_45_12;
  reg                 io_A_Valid_6_delay_46_11;
  reg                 io_A_Valid_6_delay_47_10;
  reg                 io_A_Valid_6_delay_48_9;
  reg                 io_A_Valid_6_delay_49_8;
  reg                 io_A_Valid_6_delay_50_7;
  reg                 io_A_Valid_6_delay_51_6;
  reg                 io_A_Valid_6_delay_52_5;
  reg                 io_A_Valid_6_delay_53_4;
  reg                 io_A_Valid_6_delay_54_3;
  reg                 io_A_Valid_6_delay_55_2;
  reg                 io_A_Valid_6_delay_56_1;
  reg                 io_A_Valid_6_delay_57;
  reg                 io_B_Valid_57_delay_1_5;
  reg                 io_B_Valid_57_delay_2_4;
  reg                 io_B_Valid_57_delay_3_3;
  reg                 io_B_Valid_57_delay_4_2;
  reg                 io_B_Valid_57_delay_5_1;
  reg                 io_B_Valid_57_delay_6;
  reg                 io_A_Valid_6_delay_1_57;
  reg                 io_A_Valid_6_delay_2_56;
  reg                 io_A_Valid_6_delay_3_55;
  reg                 io_A_Valid_6_delay_4_54;
  reg                 io_A_Valid_6_delay_5_53;
  reg                 io_A_Valid_6_delay_6_52;
  reg                 io_A_Valid_6_delay_7_51;
  reg                 io_A_Valid_6_delay_8_50;
  reg                 io_A_Valid_6_delay_9_49;
  reg                 io_A_Valid_6_delay_10_48;
  reg                 io_A_Valid_6_delay_11_47;
  reg                 io_A_Valid_6_delay_12_46;
  reg                 io_A_Valid_6_delay_13_45;
  reg                 io_A_Valid_6_delay_14_44;
  reg                 io_A_Valid_6_delay_15_43;
  reg                 io_A_Valid_6_delay_16_42;
  reg                 io_A_Valid_6_delay_17_41;
  reg                 io_A_Valid_6_delay_18_40;
  reg                 io_A_Valid_6_delay_19_39;
  reg                 io_A_Valid_6_delay_20_38;
  reg                 io_A_Valid_6_delay_21_37;
  reg                 io_A_Valid_6_delay_22_36;
  reg                 io_A_Valid_6_delay_23_35;
  reg                 io_A_Valid_6_delay_24_34;
  reg                 io_A_Valid_6_delay_25_33;
  reg                 io_A_Valid_6_delay_26_32;
  reg                 io_A_Valid_6_delay_27_31;
  reg                 io_A_Valid_6_delay_28_30;
  reg                 io_A_Valid_6_delay_29_29;
  reg                 io_A_Valid_6_delay_30_28;
  reg                 io_A_Valid_6_delay_31_27;
  reg                 io_A_Valid_6_delay_32_26;
  reg                 io_A_Valid_6_delay_33_25;
  reg                 io_A_Valid_6_delay_34_24;
  reg                 io_A_Valid_6_delay_35_23;
  reg                 io_A_Valid_6_delay_36_22;
  reg                 io_A_Valid_6_delay_37_21;
  reg                 io_A_Valid_6_delay_38_20;
  reg                 io_A_Valid_6_delay_39_19;
  reg                 io_A_Valid_6_delay_40_18;
  reg                 io_A_Valid_6_delay_41_17;
  reg                 io_A_Valid_6_delay_42_16;
  reg                 io_A_Valid_6_delay_43_15;
  reg                 io_A_Valid_6_delay_44_14;
  reg                 io_A_Valid_6_delay_45_13;
  reg                 io_A_Valid_6_delay_46_12;
  reg                 io_A_Valid_6_delay_47_11;
  reg                 io_A_Valid_6_delay_48_10;
  reg                 io_A_Valid_6_delay_49_9;
  reg                 io_A_Valid_6_delay_50_8;
  reg                 io_A_Valid_6_delay_51_7;
  reg                 io_A_Valid_6_delay_52_6;
  reg                 io_A_Valid_6_delay_53_5;
  reg                 io_A_Valid_6_delay_54_4;
  reg                 io_A_Valid_6_delay_55_3;
  reg                 io_A_Valid_6_delay_56_2;
  reg                 io_A_Valid_6_delay_57_1;
  reg                 io_A_Valid_6_delay_58;
  reg                 io_B_Valid_58_delay_1_5;
  reg                 io_B_Valid_58_delay_2_4;
  reg                 io_B_Valid_58_delay_3_3;
  reg                 io_B_Valid_58_delay_4_2;
  reg                 io_B_Valid_58_delay_5_1;
  reg                 io_B_Valid_58_delay_6;
  reg                 io_A_Valid_6_delay_1_58;
  reg                 io_A_Valid_6_delay_2_57;
  reg                 io_A_Valid_6_delay_3_56;
  reg                 io_A_Valid_6_delay_4_55;
  reg                 io_A_Valid_6_delay_5_54;
  reg                 io_A_Valid_6_delay_6_53;
  reg                 io_A_Valid_6_delay_7_52;
  reg                 io_A_Valid_6_delay_8_51;
  reg                 io_A_Valid_6_delay_9_50;
  reg                 io_A_Valid_6_delay_10_49;
  reg                 io_A_Valid_6_delay_11_48;
  reg                 io_A_Valid_6_delay_12_47;
  reg                 io_A_Valid_6_delay_13_46;
  reg                 io_A_Valid_6_delay_14_45;
  reg                 io_A_Valid_6_delay_15_44;
  reg                 io_A_Valid_6_delay_16_43;
  reg                 io_A_Valid_6_delay_17_42;
  reg                 io_A_Valid_6_delay_18_41;
  reg                 io_A_Valid_6_delay_19_40;
  reg                 io_A_Valid_6_delay_20_39;
  reg                 io_A_Valid_6_delay_21_38;
  reg                 io_A_Valid_6_delay_22_37;
  reg                 io_A_Valid_6_delay_23_36;
  reg                 io_A_Valid_6_delay_24_35;
  reg                 io_A_Valid_6_delay_25_34;
  reg                 io_A_Valid_6_delay_26_33;
  reg                 io_A_Valid_6_delay_27_32;
  reg                 io_A_Valid_6_delay_28_31;
  reg                 io_A_Valid_6_delay_29_30;
  reg                 io_A_Valid_6_delay_30_29;
  reg                 io_A_Valid_6_delay_31_28;
  reg                 io_A_Valid_6_delay_32_27;
  reg                 io_A_Valid_6_delay_33_26;
  reg                 io_A_Valid_6_delay_34_25;
  reg                 io_A_Valid_6_delay_35_24;
  reg                 io_A_Valid_6_delay_36_23;
  reg                 io_A_Valid_6_delay_37_22;
  reg                 io_A_Valid_6_delay_38_21;
  reg                 io_A_Valid_6_delay_39_20;
  reg                 io_A_Valid_6_delay_40_19;
  reg                 io_A_Valid_6_delay_41_18;
  reg                 io_A_Valid_6_delay_42_17;
  reg                 io_A_Valid_6_delay_43_16;
  reg                 io_A_Valid_6_delay_44_15;
  reg                 io_A_Valid_6_delay_45_14;
  reg                 io_A_Valid_6_delay_46_13;
  reg                 io_A_Valid_6_delay_47_12;
  reg                 io_A_Valid_6_delay_48_11;
  reg                 io_A_Valid_6_delay_49_10;
  reg                 io_A_Valid_6_delay_50_9;
  reg                 io_A_Valid_6_delay_51_8;
  reg                 io_A_Valid_6_delay_52_7;
  reg                 io_A_Valid_6_delay_53_6;
  reg                 io_A_Valid_6_delay_54_5;
  reg                 io_A_Valid_6_delay_55_4;
  reg                 io_A_Valid_6_delay_56_3;
  reg                 io_A_Valid_6_delay_57_2;
  reg                 io_A_Valid_6_delay_58_1;
  reg                 io_A_Valid_6_delay_59;
  reg                 io_B_Valid_59_delay_1_5;
  reg                 io_B_Valid_59_delay_2_4;
  reg                 io_B_Valid_59_delay_3_3;
  reg                 io_B_Valid_59_delay_4_2;
  reg                 io_B_Valid_59_delay_5_1;
  reg                 io_B_Valid_59_delay_6;
  reg                 io_A_Valid_6_delay_1_59;
  reg                 io_A_Valid_6_delay_2_58;
  reg                 io_A_Valid_6_delay_3_57;
  reg                 io_A_Valid_6_delay_4_56;
  reg                 io_A_Valid_6_delay_5_55;
  reg                 io_A_Valid_6_delay_6_54;
  reg                 io_A_Valid_6_delay_7_53;
  reg                 io_A_Valid_6_delay_8_52;
  reg                 io_A_Valid_6_delay_9_51;
  reg                 io_A_Valid_6_delay_10_50;
  reg                 io_A_Valid_6_delay_11_49;
  reg                 io_A_Valid_6_delay_12_48;
  reg                 io_A_Valid_6_delay_13_47;
  reg                 io_A_Valid_6_delay_14_46;
  reg                 io_A_Valid_6_delay_15_45;
  reg                 io_A_Valid_6_delay_16_44;
  reg                 io_A_Valid_6_delay_17_43;
  reg                 io_A_Valid_6_delay_18_42;
  reg                 io_A_Valid_6_delay_19_41;
  reg                 io_A_Valid_6_delay_20_40;
  reg                 io_A_Valid_6_delay_21_39;
  reg                 io_A_Valid_6_delay_22_38;
  reg                 io_A_Valid_6_delay_23_37;
  reg                 io_A_Valid_6_delay_24_36;
  reg                 io_A_Valid_6_delay_25_35;
  reg                 io_A_Valid_6_delay_26_34;
  reg                 io_A_Valid_6_delay_27_33;
  reg                 io_A_Valid_6_delay_28_32;
  reg                 io_A_Valid_6_delay_29_31;
  reg                 io_A_Valid_6_delay_30_30;
  reg                 io_A_Valid_6_delay_31_29;
  reg                 io_A_Valid_6_delay_32_28;
  reg                 io_A_Valid_6_delay_33_27;
  reg                 io_A_Valid_6_delay_34_26;
  reg                 io_A_Valid_6_delay_35_25;
  reg                 io_A_Valid_6_delay_36_24;
  reg                 io_A_Valid_6_delay_37_23;
  reg                 io_A_Valid_6_delay_38_22;
  reg                 io_A_Valid_6_delay_39_21;
  reg                 io_A_Valid_6_delay_40_20;
  reg                 io_A_Valid_6_delay_41_19;
  reg                 io_A_Valid_6_delay_42_18;
  reg                 io_A_Valid_6_delay_43_17;
  reg                 io_A_Valid_6_delay_44_16;
  reg                 io_A_Valid_6_delay_45_15;
  reg                 io_A_Valid_6_delay_46_14;
  reg                 io_A_Valid_6_delay_47_13;
  reg                 io_A_Valid_6_delay_48_12;
  reg                 io_A_Valid_6_delay_49_11;
  reg                 io_A_Valid_6_delay_50_10;
  reg                 io_A_Valid_6_delay_51_9;
  reg                 io_A_Valid_6_delay_52_8;
  reg                 io_A_Valid_6_delay_53_7;
  reg                 io_A_Valid_6_delay_54_6;
  reg                 io_A_Valid_6_delay_55_5;
  reg                 io_A_Valid_6_delay_56_4;
  reg                 io_A_Valid_6_delay_57_3;
  reg                 io_A_Valid_6_delay_58_2;
  reg                 io_A_Valid_6_delay_59_1;
  reg                 io_A_Valid_6_delay_60;
  reg                 io_B_Valid_60_delay_1_5;
  reg                 io_B_Valid_60_delay_2_4;
  reg                 io_B_Valid_60_delay_3_3;
  reg                 io_B_Valid_60_delay_4_2;
  reg                 io_B_Valid_60_delay_5_1;
  reg                 io_B_Valid_60_delay_6;
  reg                 io_A_Valid_6_delay_1_60;
  reg                 io_A_Valid_6_delay_2_59;
  reg                 io_A_Valid_6_delay_3_58;
  reg                 io_A_Valid_6_delay_4_57;
  reg                 io_A_Valid_6_delay_5_56;
  reg                 io_A_Valid_6_delay_6_55;
  reg                 io_A_Valid_6_delay_7_54;
  reg                 io_A_Valid_6_delay_8_53;
  reg                 io_A_Valid_6_delay_9_52;
  reg                 io_A_Valid_6_delay_10_51;
  reg                 io_A_Valid_6_delay_11_50;
  reg                 io_A_Valid_6_delay_12_49;
  reg                 io_A_Valid_6_delay_13_48;
  reg                 io_A_Valid_6_delay_14_47;
  reg                 io_A_Valid_6_delay_15_46;
  reg                 io_A_Valid_6_delay_16_45;
  reg                 io_A_Valid_6_delay_17_44;
  reg                 io_A_Valid_6_delay_18_43;
  reg                 io_A_Valid_6_delay_19_42;
  reg                 io_A_Valid_6_delay_20_41;
  reg                 io_A_Valid_6_delay_21_40;
  reg                 io_A_Valid_6_delay_22_39;
  reg                 io_A_Valid_6_delay_23_38;
  reg                 io_A_Valid_6_delay_24_37;
  reg                 io_A_Valid_6_delay_25_36;
  reg                 io_A_Valid_6_delay_26_35;
  reg                 io_A_Valid_6_delay_27_34;
  reg                 io_A_Valid_6_delay_28_33;
  reg                 io_A_Valid_6_delay_29_32;
  reg                 io_A_Valid_6_delay_30_31;
  reg                 io_A_Valid_6_delay_31_30;
  reg                 io_A_Valid_6_delay_32_29;
  reg                 io_A_Valid_6_delay_33_28;
  reg                 io_A_Valid_6_delay_34_27;
  reg                 io_A_Valid_6_delay_35_26;
  reg                 io_A_Valid_6_delay_36_25;
  reg                 io_A_Valid_6_delay_37_24;
  reg                 io_A_Valid_6_delay_38_23;
  reg                 io_A_Valid_6_delay_39_22;
  reg                 io_A_Valid_6_delay_40_21;
  reg                 io_A_Valid_6_delay_41_20;
  reg                 io_A_Valid_6_delay_42_19;
  reg                 io_A_Valid_6_delay_43_18;
  reg                 io_A_Valid_6_delay_44_17;
  reg                 io_A_Valid_6_delay_45_16;
  reg                 io_A_Valid_6_delay_46_15;
  reg                 io_A_Valid_6_delay_47_14;
  reg                 io_A_Valid_6_delay_48_13;
  reg                 io_A_Valid_6_delay_49_12;
  reg                 io_A_Valid_6_delay_50_11;
  reg                 io_A_Valid_6_delay_51_10;
  reg                 io_A_Valid_6_delay_52_9;
  reg                 io_A_Valid_6_delay_53_8;
  reg                 io_A_Valid_6_delay_54_7;
  reg                 io_A_Valid_6_delay_55_6;
  reg                 io_A_Valid_6_delay_56_5;
  reg                 io_A_Valid_6_delay_57_4;
  reg                 io_A_Valid_6_delay_58_3;
  reg                 io_A_Valid_6_delay_59_2;
  reg                 io_A_Valid_6_delay_60_1;
  reg                 io_A_Valid_6_delay_61;
  reg                 io_B_Valid_61_delay_1_5;
  reg                 io_B_Valid_61_delay_2_4;
  reg                 io_B_Valid_61_delay_3_3;
  reg                 io_B_Valid_61_delay_4_2;
  reg                 io_B_Valid_61_delay_5_1;
  reg                 io_B_Valid_61_delay_6;
  reg                 io_A_Valid_6_delay_1_61;
  reg                 io_A_Valid_6_delay_2_60;
  reg                 io_A_Valid_6_delay_3_59;
  reg                 io_A_Valid_6_delay_4_58;
  reg                 io_A_Valid_6_delay_5_57;
  reg                 io_A_Valid_6_delay_6_56;
  reg                 io_A_Valid_6_delay_7_55;
  reg                 io_A_Valid_6_delay_8_54;
  reg                 io_A_Valid_6_delay_9_53;
  reg                 io_A_Valid_6_delay_10_52;
  reg                 io_A_Valid_6_delay_11_51;
  reg                 io_A_Valid_6_delay_12_50;
  reg                 io_A_Valid_6_delay_13_49;
  reg                 io_A_Valid_6_delay_14_48;
  reg                 io_A_Valid_6_delay_15_47;
  reg                 io_A_Valid_6_delay_16_46;
  reg                 io_A_Valid_6_delay_17_45;
  reg                 io_A_Valid_6_delay_18_44;
  reg                 io_A_Valid_6_delay_19_43;
  reg                 io_A_Valid_6_delay_20_42;
  reg                 io_A_Valid_6_delay_21_41;
  reg                 io_A_Valid_6_delay_22_40;
  reg                 io_A_Valid_6_delay_23_39;
  reg                 io_A_Valid_6_delay_24_38;
  reg                 io_A_Valid_6_delay_25_37;
  reg                 io_A_Valid_6_delay_26_36;
  reg                 io_A_Valid_6_delay_27_35;
  reg                 io_A_Valid_6_delay_28_34;
  reg                 io_A_Valid_6_delay_29_33;
  reg                 io_A_Valid_6_delay_30_32;
  reg                 io_A_Valid_6_delay_31_31;
  reg                 io_A_Valid_6_delay_32_30;
  reg                 io_A_Valid_6_delay_33_29;
  reg                 io_A_Valid_6_delay_34_28;
  reg                 io_A_Valid_6_delay_35_27;
  reg                 io_A_Valid_6_delay_36_26;
  reg                 io_A_Valid_6_delay_37_25;
  reg                 io_A_Valid_6_delay_38_24;
  reg                 io_A_Valid_6_delay_39_23;
  reg                 io_A_Valid_6_delay_40_22;
  reg                 io_A_Valid_6_delay_41_21;
  reg                 io_A_Valid_6_delay_42_20;
  reg                 io_A_Valid_6_delay_43_19;
  reg                 io_A_Valid_6_delay_44_18;
  reg                 io_A_Valid_6_delay_45_17;
  reg                 io_A_Valid_6_delay_46_16;
  reg                 io_A_Valid_6_delay_47_15;
  reg                 io_A_Valid_6_delay_48_14;
  reg                 io_A_Valid_6_delay_49_13;
  reg                 io_A_Valid_6_delay_50_12;
  reg                 io_A_Valid_6_delay_51_11;
  reg                 io_A_Valid_6_delay_52_10;
  reg                 io_A_Valid_6_delay_53_9;
  reg                 io_A_Valid_6_delay_54_8;
  reg                 io_A_Valid_6_delay_55_7;
  reg                 io_A_Valid_6_delay_56_6;
  reg                 io_A_Valid_6_delay_57_5;
  reg                 io_A_Valid_6_delay_58_4;
  reg                 io_A_Valid_6_delay_59_3;
  reg                 io_A_Valid_6_delay_60_2;
  reg                 io_A_Valid_6_delay_61_1;
  reg                 io_A_Valid_6_delay_62;
  reg                 io_B_Valid_62_delay_1_5;
  reg                 io_B_Valid_62_delay_2_4;
  reg                 io_B_Valid_62_delay_3_3;
  reg                 io_B_Valid_62_delay_4_2;
  reg                 io_B_Valid_62_delay_5_1;
  reg                 io_B_Valid_62_delay_6;
  reg                 io_A_Valid_6_delay_1_62;
  reg                 io_A_Valid_6_delay_2_61;
  reg                 io_A_Valid_6_delay_3_60;
  reg                 io_A_Valid_6_delay_4_59;
  reg                 io_A_Valid_6_delay_5_58;
  reg                 io_A_Valid_6_delay_6_57;
  reg                 io_A_Valid_6_delay_7_56;
  reg                 io_A_Valid_6_delay_8_55;
  reg                 io_A_Valid_6_delay_9_54;
  reg                 io_A_Valid_6_delay_10_53;
  reg                 io_A_Valid_6_delay_11_52;
  reg                 io_A_Valid_6_delay_12_51;
  reg                 io_A_Valid_6_delay_13_50;
  reg                 io_A_Valid_6_delay_14_49;
  reg                 io_A_Valid_6_delay_15_48;
  reg                 io_A_Valid_6_delay_16_47;
  reg                 io_A_Valid_6_delay_17_46;
  reg                 io_A_Valid_6_delay_18_45;
  reg                 io_A_Valid_6_delay_19_44;
  reg                 io_A_Valid_6_delay_20_43;
  reg                 io_A_Valid_6_delay_21_42;
  reg                 io_A_Valid_6_delay_22_41;
  reg                 io_A_Valid_6_delay_23_40;
  reg                 io_A_Valid_6_delay_24_39;
  reg                 io_A_Valid_6_delay_25_38;
  reg                 io_A_Valid_6_delay_26_37;
  reg                 io_A_Valid_6_delay_27_36;
  reg                 io_A_Valid_6_delay_28_35;
  reg                 io_A_Valid_6_delay_29_34;
  reg                 io_A_Valid_6_delay_30_33;
  reg                 io_A_Valid_6_delay_31_32;
  reg                 io_A_Valid_6_delay_32_31;
  reg                 io_A_Valid_6_delay_33_30;
  reg                 io_A_Valid_6_delay_34_29;
  reg                 io_A_Valid_6_delay_35_28;
  reg                 io_A_Valid_6_delay_36_27;
  reg                 io_A_Valid_6_delay_37_26;
  reg                 io_A_Valid_6_delay_38_25;
  reg                 io_A_Valid_6_delay_39_24;
  reg                 io_A_Valid_6_delay_40_23;
  reg                 io_A_Valid_6_delay_41_22;
  reg                 io_A_Valid_6_delay_42_21;
  reg                 io_A_Valid_6_delay_43_20;
  reg                 io_A_Valid_6_delay_44_19;
  reg                 io_A_Valid_6_delay_45_18;
  reg                 io_A_Valid_6_delay_46_17;
  reg                 io_A_Valid_6_delay_47_16;
  reg                 io_A_Valid_6_delay_48_15;
  reg                 io_A_Valid_6_delay_49_14;
  reg                 io_A_Valid_6_delay_50_13;
  reg                 io_A_Valid_6_delay_51_12;
  reg                 io_A_Valid_6_delay_52_11;
  reg                 io_A_Valid_6_delay_53_10;
  reg                 io_A_Valid_6_delay_54_9;
  reg                 io_A_Valid_6_delay_55_8;
  reg                 io_A_Valid_6_delay_56_7;
  reg                 io_A_Valid_6_delay_57_6;
  reg                 io_A_Valid_6_delay_58_5;
  reg                 io_A_Valid_6_delay_59_4;
  reg                 io_A_Valid_6_delay_60_3;
  reg                 io_A_Valid_6_delay_61_2;
  reg                 io_A_Valid_6_delay_62_1;
  reg                 io_A_Valid_6_delay_63;
  reg                 io_B_Valid_63_delay_1_5;
  reg                 io_B_Valid_63_delay_2_4;
  reg                 io_B_Valid_63_delay_3_3;
  reg                 io_B_Valid_63_delay_4_2;
  reg                 io_B_Valid_63_delay_5_1;
  reg                 io_B_Valid_63_delay_6;
  reg        [15:0]   io_signCount_regNextWhen_7;
  reg                 io_B_Valid_0_delay_1_6;
  reg                 io_B_Valid_0_delay_2_5;
  reg                 io_B_Valid_0_delay_3_4;
  reg                 io_B_Valid_0_delay_4_3;
  reg                 io_B_Valid_0_delay_5_2;
  reg                 io_B_Valid_0_delay_6_1;
  reg                 io_B_Valid_0_delay_7;
  reg                 io_A_Valid_7_delay_1;
  reg                 io_B_Valid_1_delay_1_6;
  reg                 io_B_Valid_1_delay_2_5;
  reg                 io_B_Valid_1_delay_3_4;
  reg                 io_B_Valid_1_delay_4_3;
  reg                 io_B_Valid_1_delay_5_2;
  reg                 io_B_Valid_1_delay_6_1;
  reg                 io_B_Valid_1_delay_7;
  reg                 io_A_Valid_7_delay_1_1;
  reg                 io_A_Valid_7_delay_2;
  reg                 io_B_Valid_2_delay_1_6;
  reg                 io_B_Valid_2_delay_2_5;
  reg                 io_B_Valid_2_delay_3_4;
  reg                 io_B_Valid_2_delay_4_3;
  reg                 io_B_Valid_2_delay_5_2;
  reg                 io_B_Valid_2_delay_6_1;
  reg                 io_B_Valid_2_delay_7;
  reg                 io_A_Valid_7_delay_1_2;
  reg                 io_A_Valid_7_delay_2_1;
  reg                 io_A_Valid_7_delay_3;
  reg                 io_B_Valid_3_delay_1_6;
  reg                 io_B_Valid_3_delay_2_5;
  reg                 io_B_Valid_3_delay_3_4;
  reg                 io_B_Valid_3_delay_4_3;
  reg                 io_B_Valid_3_delay_5_2;
  reg                 io_B_Valid_3_delay_6_1;
  reg                 io_B_Valid_3_delay_7;
  reg                 io_A_Valid_7_delay_1_3;
  reg                 io_A_Valid_7_delay_2_2;
  reg                 io_A_Valid_7_delay_3_1;
  reg                 io_A_Valid_7_delay_4;
  reg                 io_B_Valid_4_delay_1_6;
  reg                 io_B_Valid_4_delay_2_5;
  reg                 io_B_Valid_4_delay_3_4;
  reg                 io_B_Valid_4_delay_4_3;
  reg                 io_B_Valid_4_delay_5_2;
  reg                 io_B_Valid_4_delay_6_1;
  reg                 io_B_Valid_4_delay_7;
  reg                 io_A_Valid_7_delay_1_4;
  reg                 io_A_Valid_7_delay_2_3;
  reg                 io_A_Valid_7_delay_3_2;
  reg                 io_A_Valid_7_delay_4_1;
  reg                 io_A_Valid_7_delay_5;
  reg                 io_B_Valid_5_delay_1_6;
  reg                 io_B_Valid_5_delay_2_5;
  reg                 io_B_Valid_5_delay_3_4;
  reg                 io_B_Valid_5_delay_4_3;
  reg                 io_B_Valid_5_delay_5_2;
  reg                 io_B_Valid_5_delay_6_1;
  reg                 io_B_Valid_5_delay_7;
  reg                 io_A_Valid_7_delay_1_5;
  reg                 io_A_Valid_7_delay_2_4;
  reg                 io_A_Valid_7_delay_3_3;
  reg                 io_A_Valid_7_delay_4_2;
  reg                 io_A_Valid_7_delay_5_1;
  reg                 io_A_Valid_7_delay_6;
  reg                 io_B_Valid_6_delay_1_6;
  reg                 io_B_Valid_6_delay_2_5;
  reg                 io_B_Valid_6_delay_3_4;
  reg                 io_B_Valid_6_delay_4_3;
  reg                 io_B_Valid_6_delay_5_2;
  reg                 io_B_Valid_6_delay_6_1;
  reg                 io_B_Valid_6_delay_7;
  reg                 io_A_Valid_7_delay_1_6;
  reg                 io_A_Valid_7_delay_2_5;
  reg                 io_A_Valid_7_delay_3_4;
  reg                 io_A_Valid_7_delay_4_3;
  reg                 io_A_Valid_7_delay_5_2;
  reg                 io_A_Valid_7_delay_6_1;
  reg                 io_A_Valid_7_delay_7;
  reg                 io_B_Valid_7_delay_1_6;
  reg                 io_B_Valid_7_delay_2_5;
  reg                 io_B_Valid_7_delay_3_4;
  reg                 io_B_Valid_7_delay_4_3;
  reg                 io_B_Valid_7_delay_5_2;
  reg                 io_B_Valid_7_delay_6_1;
  reg                 io_B_Valid_7_delay_7;
  reg                 io_A_Valid_7_delay_1_7;
  reg                 io_A_Valid_7_delay_2_6;
  reg                 io_A_Valid_7_delay_3_5;
  reg                 io_A_Valid_7_delay_4_4;
  reg                 io_A_Valid_7_delay_5_3;
  reg                 io_A_Valid_7_delay_6_2;
  reg                 io_A_Valid_7_delay_7_1;
  reg                 io_A_Valid_7_delay_8;
  reg                 io_B_Valid_8_delay_1_6;
  reg                 io_B_Valid_8_delay_2_5;
  reg                 io_B_Valid_8_delay_3_4;
  reg                 io_B_Valid_8_delay_4_3;
  reg                 io_B_Valid_8_delay_5_2;
  reg                 io_B_Valid_8_delay_6_1;
  reg                 io_B_Valid_8_delay_7;
  reg                 io_A_Valid_7_delay_1_8;
  reg                 io_A_Valid_7_delay_2_7;
  reg                 io_A_Valid_7_delay_3_6;
  reg                 io_A_Valid_7_delay_4_5;
  reg                 io_A_Valid_7_delay_5_4;
  reg                 io_A_Valid_7_delay_6_3;
  reg                 io_A_Valid_7_delay_7_2;
  reg                 io_A_Valid_7_delay_8_1;
  reg                 io_A_Valid_7_delay_9;
  reg                 io_B_Valid_9_delay_1_6;
  reg                 io_B_Valid_9_delay_2_5;
  reg                 io_B_Valid_9_delay_3_4;
  reg                 io_B_Valid_9_delay_4_3;
  reg                 io_B_Valid_9_delay_5_2;
  reg                 io_B_Valid_9_delay_6_1;
  reg                 io_B_Valid_9_delay_7;
  reg                 io_A_Valid_7_delay_1_9;
  reg                 io_A_Valid_7_delay_2_8;
  reg                 io_A_Valid_7_delay_3_7;
  reg                 io_A_Valid_7_delay_4_6;
  reg                 io_A_Valid_7_delay_5_5;
  reg                 io_A_Valid_7_delay_6_4;
  reg                 io_A_Valid_7_delay_7_3;
  reg                 io_A_Valid_7_delay_8_2;
  reg                 io_A_Valid_7_delay_9_1;
  reg                 io_A_Valid_7_delay_10;
  reg                 io_B_Valid_10_delay_1_6;
  reg                 io_B_Valid_10_delay_2_5;
  reg                 io_B_Valid_10_delay_3_4;
  reg                 io_B_Valid_10_delay_4_3;
  reg                 io_B_Valid_10_delay_5_2;
  reg                 io_B_Valid_10_delay_6_1;
  reg                 io_B_Valid_10_delay_7;
  reg                 io_A_Valid_7_delay_1_10;
  reg                 io_A_Valid_7_delay_2_9;
  reg                 io_A_Valid_7_delay_3_8;
  reg                 io_A_Valid_7_delay_4_7;
  reg                 io_A_Valid_7_delay_5_6;
  reg                 io_A_Valid_7_delay_6_5;
  reg                 io_A_Valid_7_delay_7_4;
  reg                 io_A_Valid_7_delay_8_3;
  reg                 io_A_Valid_7_delay_9_2;
  reg                 io_A_Valid_7_delay_10_1;
  reg                 io_A_Valid_7_delay_11;
  reg                 io_B_Valid_11_delay_1_6;
  reg                 io_B_Valid_11_delay_2_5;
  reg                 io_B_Valid_11_delay_3_4;
  reg                 io_B_Valid_11_delay_4_3;
  reg                 io_B_Valid_11_delay_5_2;
  reg                 io_B_Valid_11_delay_6_1;
  reg                 io_B_Valid_11_delay_7;
  reg                 io_A_Valid_7_delay_1_11;
  reg                 io_A_Valid_7_delay_2_10;
  reg                 io_A_Valid_7_delay_3_9;
  reg                 io_A_Valid_7_delay_4_8;
  reg                 io_A_Valid_7_delay_5_7;
  reg                 io_A_Valid_7_delay_6_6;
  reg                 io_A_Valid_7_delay_7_5;
  reg                 io_A_Valid_7_delay_8_4;
  reg                 io_A_Valid_7_delay_9_3;
  reg                 io_A_Valid_7_delay_10_2;
  reg                 io_A_Valid_7_delay_11_1;
  reg                 io_A_Valid_7_delay_12;
  reg                 io_B_Valid_12_delay_1_6;
  reg                 io_B_Valid_12_delay_2_5;
  reg                 io_B_Valid_12_delay_3_4;
  reg                 io_B_Valid_12_delay_4_3;
  reg                 io_B_Valid_12_delay_5_2;
  reg                 io_B_Valid_12_delay_6_1;
  reg                 io_B_Valid_12_delay_7;
  reg                 io_A_Valid_7_delay_1_12;
  reg                 io_A_Valid_7_delay_2_11;
  reg                 io_A_Valid_7_delay_3_10;
  reg                 io_A_Valid_7_delay_4_9;
  reg                 io_A_Valid_7_delay_5_8;
  reg                 io_A_Valid_7_delay_6_7;
  reg                 io_A_Valid_7_delay_7_6;
  reg                 io_A_Valid_7_delay_8_5;
  reg                 io_A_Valid_7_delay_9_4;
  reg                 io_A_Valid_7_delay_10_3;
  reg                 io_A_Valid_7_delay_11_2;
  reg                 io_A_Valid_7_delay_12_1;
  reg                 io_A_Valid_7_delay_13;
  reg                 io_B_Valid_13_delay_1_6;
  reg                 io_B_Valid_13_delay_2_5;
  reg                 io_B_Valid_13_delay_3_4;
  reg                 io_B_Valid_13_delay_4_3;
  reg                 io_B_Valid_13_delay_5_2;
  reg                 io_B_Valid_13_delay_6_1;
  reg                 io_B_Valid_13_delay_7;
  reg                 io_A_Valid_7_delay_1_13;
  reg                 io_A_Valid_7_delay_2_12;
  reg                 io_A_Valid_7_delay_3_11;
  reg                 io_A_Valid_7_delay_4_10;
  reg                 io_A_Valid_7_delay_5_9;
  reg                 io_A_Valid_7_delay_6_8;
  reg                 io_A_Valid_7_delay_7_7;
  reg                 io_A_Valid_7_delay_8_6;
  reg                 io_A_Valid_7_delay_9_5;
  reg                 io_A_Valid_7_delay_10_4;
  reg                 io_A_Valid_7_delay_11_3;
  reg                 io_A_Valid_7_delay_12_2;
  reg                 io_A_Valid_7_delay_13_1;
  reg                 io_A_Valid_7_delay_14;
  reg                 io_B_Valid_14_delay_1_6;
  reg                 io_B_Valid_14_delay_2_5;
  reg                 io_B_Valid_14_delay_3_4;
  reg                 io_B_Valid_14_delay_4_3;
  reg                 io_B_Valid_14_delay_5_2;
  reg                 io_B_Valid_14_delay_6_1;
  reg                 io_B_Valid_14_delay_7;
  reg                 io_A_Valid_7_delay_1_14;
  reg                 io_A_Valid_7_delay_2_13;
  reg                 io_A_Valid_7_delay_3_12;
  reg                 io_A_Valid_7_delay_4_11;
  reg                 io_A_Valid_7_delay_5_10;
  reg                 io_A_Valid_7_delay_6_9;
  reg                 io_A_Valid_7_delay_7_8;
  reg                 io_A_Valid_7_delay_8_7;
  reg                 io_A_Valid_7_delay_9_6;
  reg                 io_A_Valid_7_delay_10_5;
  reg                 io_A_Valid_7_delay_11_4;
  reg                 io_A_Valid_7_delay_12_3;
  reg                 io_A_Valid_7_delay_13_2;
  reg                 io_A_Valid_7_delay_14_1;
  reg                 io_A_Valid_7_delay_15;
  reg                 io_B_Valid_15_delay_1_6;
  reg                 io_B_Valid_15_delay_2_5;
  reg                 io_B_Valid_15_delay_3_4;
  reg                 io_B_Valid_15_delay_4_3;
  reg                 io_B_Valid_15_delay_5_2;
  reg                 io_B_Valid_15_delay_6_1;
  reg                 io_B_Valid_15_delay_7;
  reg                 io_A_Valid_7_delay_1_15;
  reg                 io_A_Valid_7_delay_2_14;
  reg                 io_A_Valid_7_delay_3_13;
  reg                 io_A_Valid_7_delay_4_12;
  reg                 io_A_Valid_7_delay_5_11;
  reg                 io_A_Valid_7_delay_6_10;
  reg                 io_A_Valid_7_delay_7_9;
  reg                 io_A_Valid_7_delay_8_8;
  reg                 io_A_Valid_7_delay_9_7;
  reg                 io_A_Valid_7_delay_10_6;
  reg                 io_A_Valid_7_delay_11_5;
  reg                 io_A_Valid_7_delay_12_4;
  reg                 io_A_Valid_7_delay_13_3;
  reg                 io_A_Valid_7_delay_14_2;
  reg                 io_A_Valid_7_delay_15_1;
  reg                 io_A_Valid_7_delay_16;
  reg                 io_B_Valid_16_delay_1_6;
  reg                 io_B_Valid_16_delay_2_5;
  reg                 io_B_Valid_16_delay_3_4;
  reg                 io_B_Valid_16_delay_4_3;
  reg                 io_B_Valid_16_delay_5_2;
  reg                 io_B_Valid_16_delay_6_1;
  reg                 io_B_Valid_16_delay_7;
  reg                 io_A_Valid_7_delay_1_16;
  reg                 io_A_Valid_7_delay_2_15;
  reg                 io_A_Valid_7_delay_3_14;
  reg                 io_A_Valid_7_delay_4_13;
  reg                 io_A_Valid_7_delay_5_12;
  reg                 io_A_Valid_7_delay_6_11;
  reg                 io_A_Valid_7_delay_7_10;
  reg                 io_A_Valid_7_delay_8_9;
  reg                 io_A_Valid_7_delay_9_8;
  reg                 io_A_Valid_7_delay_10_7;
  reg                 io_A_Valid_7_delay_11_6;
  reg                 io_A_Valid_7_delay_12_5;
  reg                 io_A_Valid_7_delay_13_4;
  reg                 io_A_Valid_7_delay_14_3;
  reg                 io_A_Valid_7_delay_15_2;
  reg                 io_A_Valid_7_delay_16_1;
  reg                 io_A_Valid_7_delay_17;
  reg                 io_B_Valid_17_delay_1_6;
  reg                 io_B_Valid_17_delay_2_5;
  reg                 io_B_Valid_17_delay_3_4;
  reg                 io_B_Valid_17_delay_4_3;
  reg                 io_B_Valid_17_delay_5_2;
  reg                 io_B_Valid_17_delay_6_1;
  reg                 io_B_Valid_17_delay_7;
  reg                 io_A_Valid_7_delay_1_17;
  reg                 io_A_Valid_7_delay_2_16;
  reg                 io_A_Valid_7_delay_3_15;
  reg                 io_A_Valid_7_delay_4_14;
  reg                 io_A_Valid_7_delay_5_13;
  reg                 io_A_Valid_7_delay_6_12;
  reg                 io_A_Valid_7_delay_7_11;
  reg                 io_A_Valid_7_delay_8_10;
  reg                 io_A_Valid_7_delay_9_9;
  reg                 io_A_Valid_7_delay_10_8;
  reg                 io_A_Valid_7_delay_11_7;
  reg                 io_A_Valid_7_delay_12_6;
  reg                 io_A_Valid_7_delay_13_5;
  reg                 io_A_Valid_7_delay_14_4;
  reg                 io_A_Valid_7_delay_15_3;
  reg                 io_A_Valid_7_delay_16_2;
  reg                 io_A_Valid_7_delay_17_1;
  reg                 io_A_Valid_7_delay_18;
  reg                 io_B_Valid_18_delay_1_6;
  reg                 io_B_Valid_18_delay_2_5;
  reg                 io_B_Valid_18_delay_3_4;
  reg                 io_B_Valid_18_delay_4_3;
  reg                 io_B_Valid_18_delay_5_2;
  reg                 io_B_Valid_18_delay_6_1;
  reg                 io_B_Valid_18_delay_7;
  reg                 io_A_Valid_7_delay_1_18;
  reg                 io_A_Valid_7_delay_2_17;
  reg                 io_A_Valid_7_delay_3_16;
  reg                 io_A_Valid_7_delay_4_15;
  reg                 io_A_Valid_7_delay_5_14;
  reg                 io_A_Valid_7_delay_6_13;
  reg                 io_A_Valid_7_delay_7_12;
  reg                 io_A_Valid_7_delay_8_11;
  reg                 io_A_Valid_7_delay_9_10;
  reg                 io_A_Valid_7_delay_10_9;
  reg                 io_A_Valid_7_delay_11_8;
  reg                 io_A_Valid_7_delay_12_7;
  reg                 io_A_Valid_7_delay_13_6;
  reg                 io_A_Valid_7_delay_14_5;
  reg                 io_A_Valid_7_delay_15_4;
  reg                 io_A_Valid_7_delay_16_3;
  reg                 io_A_Valid_7_delay_17_2;
  reg                 io_A_Valid_7_delay_18_1;
  reg                 io_A_Valid_7_delay_19;
  reg                 io_B_Valid_19_delay_1_6;
  reg                 io_B_Valid_19_delay_2_5;
  reg                 io_B_Valid_19_delay_3_4;
  reg                 io_B_Valid_19_delay_4_3;
  reg                 io_B_Valid_19_delay_5_2;
  reg                 io_B_Valid_19_delay_6_1;
  reg                 io_B_Valid_19_delay_7;
  reg                 io_A_Valid_7_delay_1_19;
  reg                 io_A_Valid_7_delay_2_18;
  reg                 io_A_Valid_7_delay_3_17;
  reg                 io_A_Valid_7_delay_4_16;
  reg                 io_A_Valid_7_delay_5_15;
  reg                 io_A_Valid_7_delay_6_14;
  reg                 io_A_Valid_7_delay_7_13;
  reg                 io_A_Valid_7_delay_8_12;
  reg                 io_A_Valid_7_delay_9_11;
  reg                 io_A_Valid_7_delay_10_10;
  reg                 io_A_Valid_7_delay_11_9;
  reg                 io_A_Valid_7_delay_12_8;
  reg                 io_A_Valid_7_delay_13_7;
  reg                 io_A_Valid_7_delay_14_6;
  reg                 io_A_Valid_7_delay_15_5;
  reg                 io_A_Valid_7_delay_16_4;
  reg                 io_A_Valid_7_delay_17_3;
  reg                 io_A_Valid_7_delay_18_2;
  reg                 io_A_Valid_7_delay_19_1;
  reg                 io_A_Valid_7_delay_20;
  reg                 io_B_Valid_20_delay_1_6;
  reg                 io_B_Valid_20_delay_2_5;
  reg                 io_B_Valid_20_delay_3_4;
  reg                 io_B_Valid_20_delay_4_3;
  reg                 io_B_Valid_20_delay_5_2;
  reg                 io_B_Valid_20_delay_6_1;
  reg                 io_B_Valid_20_delay_7;
  reg                 io_A_Valid_7_delay_1_20;
  reg                 io_A_Valid_7_delay_2_19;
  reg                 io_A_Valid_7_delay_3_18;
  reg                 io_A_Valid_7_delay_4_17;
  reg                 io_A_Valid_7_delay_5_16;
  reg                 io_A_Valid_7_delay_6_15;
  reg                 io_A_Valid_7_delay_7_14;
  reg                 io_A_Valid_7_delay_8_13;
  reg                 io_A_Valid_7_delay_9_12;
  reg                 io_A_Valid_7_delay_10_11;
  reg                 io_A_Valid_7_delay_11_10;
  reg                 io_A_Valid_7_delay_12_9;
  reg                 io_A_Valid_7_delay_13_8;
  reg                 io_A_Valid_7_delay_14_7;
  reg                 io_A_Valid_7_delay_15_6;
  reg                 io_A_Valid_7_delay_16_5;
  reg                 io_A_Valid_7_delay_17_4;
  reg                 io_A_Valid_7_delay_18_3;
  reg                 io_A_Valid_7_delay_19_2;
  reg                 io_A_Valid_7_delay_20_1;
  reg                 io_A_Valid_7_delay_21;
  reg                 io_B_Valid_21_delay_1_6;
  reg                 io_B_Valid_21_delay_2_5;
  reg                 io_B_Valid_21_delay_3_4;
  reg                 io_B_Valid_21_delay_4_3;
  reg                 io_B_Valid_21_delay_5_2;
  reg                 io_B_Valid_21_delay_6_1;
  reg                 io_B_Valid_21_delay_7;
  reg                 io_A_Valid_7_delay_1_21;
  reg                 io_A_Valid_7_delay_2_20;
  reg                 io_A_Valid_7_delay_3_19;
  reg                 io_A_Valid_7_delay_4_18;
  reg                 io_A_Valid_7_delay_5_17;
  reg                 io_A_Valid_7_delay_6_16;
  reg                 io_A_Valid_7_delay_7_15;
  reg                 io_A_Valid_7_delay_8_14;
  reg                 io_A_Valid_7_delay_9_13;
  reg                 io_A_Valid_7_delay_10_12;
  reg                 io_A_Valid_7_delay_11_11;
  reg                 io_A_Valid_7_delay_12_10;
  reg                 io_A_Valid_7_delay_13_9;
  reg                 io_A_Valid_7_delay_14_8;
  reg                 io_A_Valid_7_delay_15_7;
  reg                 io_A_Valid_7_delay_16_6;
  reg                 io_A_Valid_7_delay_17_5;
  reg                 io_A_Valid_7_delay_18_4;
  reg                 io_A_Valid_7_delay_19_3;
  reg                 io_A_Valid_7_delay_20_2;
  reg                 io_A_Valid_7_delay_21_1;
  reg                 io_A_Valid_7_delay_22;
  reg                 io_B_Valid_22_delay_1_6;
  reg                 io_B_Valid_22_delay_2_5;
  reg                 io_B_Valid_22_delay_3_4;
  reg                 io_B_Valid_22_delay_4_3;
  reg                 io_B_Valid_22_delay_5_2;
  reg                 io_B_Valid_22_delay_6_1;
  reg                 io_B_Valid_22_delay_7;
  reg                 io_A_Valid_7_delay_1_22;
  reg                 io_A_Valid_7_delay_2_21;
  reg                 io_A_Valid_7_delay_3_20;
  reg                 io_A_Valid_7_delay_4_19;
  reg                 io_A_Valid_7_delay_5_18;
  reg                 io_A_Valid_7_delay_6_17;
  reg                 io_A_Valid_7_delay_7_16;
  reg                 io_A_Valid_7_delay_8_15;
  reg                 io_A_Valid_7_delay_9_14;
  reg                 io_A_Valid_7_delay_10_13;
  reg                 io_A_Valid_7_delay_11_12;
  reg                 io_A_Valid_7_delay_12_11;
  reg                 io_A_Valid_7_delay_13_10;
  reg                 io_A_Valid_7_delay_14_9;
  reg                 io_A_Valid_7_delay_15_8;
  reg                 io_A_Valid_7_delay_16_7;
  reg                 io_A_Valid_7_delay_17_6;
  reg                 io_A_Valid_7_delay_18_5;
  reg                 io_A_Valid_7_delay_19_4;
  reg                 io_A_Valid_7_delay_20_3;
  reg                 io_A_Valid_7_delay_21_2;
  reg                 io_A_Valid_7_delay_22_1;
  reg                 io_A_Valid_7_delay_23;
  reg                 io_B_Valid_23_delay_1_6;
  reg                 io_B_Valid_23_delay_2_5;
  reg                 io_B_Valid_23_delay_3_4;
  reg                 io_B_Valid_23_delay_4_3;
  reg                 io_B_Valid_23_delay_5_2;
  reg                 io_B_Valid_23_delay_6_1;
  reg                 io_B_Valid_23_delay_7;
  reg                 io_A_Valid_7_delay_1_23;
  reg                 io_A_Valid_7_delay_2_22;
  reg                 io_A_Valid_7_delay_3_21;
  reg                 io_A_Valid_7_delay_4_20;
  reg                 io_A_Valid_7_delay_5_19;
  reg                 io_A_Valid_7_delay_6_18;
  reg                 io_A_Valid_7_delay_7_17;
  reg                 io_A_Valid_7_delay_8_16;
  reg                 io_A_Valid_7_delay_9_15;
  reg                 io_A_Valid_7_delay_10_14;
  reg                 io_A_Valid_7_delay_11_13;
  reg                 io_A_Valid_7_delay_12_12;
  reg                 io_A_Valid_7_delay_13_11;
  reg                 io_A_Valid_7_delay_14_10;
  reg                 io_A_Valid_7_delay_15_9;
  reg                 io_A_Valid_7_delay_16_8;
  reg                 io_A_Valid_7_delay_17_7;
  reg                 io_A_Valid_7_delay_18_6;
  reg                 io_A_Valid_7_delay_19_5;
  reg                 io_A_Valid_7_delay_20_4;
  reg                 io_A_Valid_7_delay_21_3;
  reg                 io_A_Valid_7_delay_22_2;
  reg                 io_A_Valid_7_delay_23_1;
  reg                 io_A_Valid_7_delay_24;
  reg                 io_B_Valid_24_delay_1_6;
  reg                 io_B_Valid_24_delay_2_5;
  reg                 io_B_Valid_24_delay_3_4;
  reg                 io_B_Valid_24_delay_4_3;
  reg                 io_B_Valid_24_delay_5_2;
  reg                 io_B_Valid_24_delay_6_1;
  reg                 io_B_Valid_24_delay_7;
  reg                 io_A_Valid_7_delay_1_24;
  reg                 io_A_Valid_7_delay_2_23;
  reg                 io_A_Valid_7_delay_3_22;
  reg                 io_A_Valid_7_delay_4_21;
  reg                 io_A_Valid_7_delay_5_20;
  reg                 io_A_Valid_7_delay_6_19;
  reg                 io_A_Valid_7_delay_7_18;
  reg                 io_A_Valid_7_delay_8_17;
  reg                 io_A_Valid_7_delay_9_16;
  reg                 io_A_Valid_7_delay_10_15;
  reg                 io_A_Valid_7_delay_11_14;
  reg                 io_A_Valid_7_delay_12_13;
  reg                 io_A_Valid_7_delay_13_12;
  reg                 io_A_Valid_7_delay_14_11;
  reg                 io_A_Valid_7_delay_15_10;
  reg                 io_A_Valid_7_delay_16_9;
  reg                 io_A_Valid_7_delay_17_8;
  reg                 io_A_Valid_7_delay_18_7;
  reg                 io_A_Valid_7_delay_19_6;
  reg                 io_A_Valid_7_delay_20_5;
  reg                 io_A_Valid_7_delay_21_4;
  reg                 io_A_Valid_7_delay_22_3;
  reg                 io_A_Valid_7_delay_23_2;
  reg                 io_A_Valid_7_delay_24_1;
  reg                 io_A_Valid_7_delay_25;
  reg                 io_B_Valid_25_delay_1_6;
  reg                 io_B_Valid_25_delay_2_5;
  reg                 io_B_Valid_25_delay_3_4;
  reg                 io_B_Valid_25_delay_4_3;
  reg                 io_B_Valid_25_delay_5_2;
  reg                 io_B_Valid_25_delay_6_1;
  reg                 io_B_Valid_25_delay_7;
  reg                 io_A_Valid_7_delay_1_25;
  reg                 io_A_Valid_7_delay_2_24;
  reg                 io_A_Valid_7_delay_3_23;
  reg                 io_A_Valid_7_delay_4_22;
  reg                 io_A_Valid_7_delay_5_21;
  reg                 io_A_Valid_7_delay_6_20;
  reg                 io_A_Valid_7_delay_7_19;
  reg                 io_A_Valid_7_delay_8_18;
  reg                 io_A_Valid_7_delay_9_17;
  reg                 io_A_Valid_7_delay_10_16;
  reg                 io_A_Valid_7_delay_11_15;
  reg                 io_A_Valid_7_delay_12_14;
  reg                 io_A_Valid_7_delay_13_13;
  reg                 io_A_Valid_7_delay_14_12;
  reg                 io_A_Valid_7_delay_15_11;
  reg                 io_A_Valid_7_delay_16_10;
  reg                 io_A_Valid_7_delay_17_9;
  reg                 io_A_Valid_7_delay_18_8;
  reg                 io_A_Valid_7_delay_19_7;
  reg                 io_A_Valid_7_delay_20_6;
  reg                 io_A_Valid_7_delay_21_5;
  reg                 io_A_Valid_7_delay_22_4;
  reg                 io_A_Valid_7_delay_23_3;
  reg                 io_A_Valid_7_delay_24_2;
  reg                 io_A_Valid_7_delay_25_1;
  reg                 io_A_Valid_7_delay_26;
  reg                 io_B_Valid_26_delay_1_6;
  reg                 io_B_Valid_26_delay_2_5;
  reg                 io_B_Valid_26_delay_3_4;
  reg                 io_B_Valid_26_delay_4_3;
  reg                 io_B_Valid_26_delay_5_2;
  reg                 io_B_Valid_26_delay_6_1;
  reg                 io_B_Valid_26_delay_7;
  reg                 io_A_Valid_7_delay_1_26;
  reg                 io_A_Valid_7_delay_2_25;
  reg                 io_A_Valid_7_delay_3_24;
  reg                 io_A_Valid_7_delay_4_23;
  reg                 io_A_Valid_7_delay_5_22;
  reg                 io_A_Valid_7_delay_6_21;
  reg                 io_A_Valid_7_delay_7_20;
  reg                 io_A_Valid_7_delay_8_19;
  reg                 io_A_Valid_7_delay_9_18;
  reg                 io_A_Valid_7_delay_10_17;
  reg                 io_A_Valid_7_delay_11_16;
  reg                 io_A_Valid_7_delay_12_15;
  reg                 io_A_Valid_7_delay_13_14;
  reg                 io_A_Valid_7_delay_14_13;
  reg                 io_A_Valid_7_delay_15_12;
  reg                 io_A_Valid_7_delay_16_11;
  reg                 io_A_Valid_7_delay_17_10;
  reg                 io_A_Valid_7_delay_18_9;
  reg                 io_A_Valid_7_delay_19_8;
  reg                 io_A_Valid_7_delay_20_7;
  reg                 io_A_Valid_7_delay_21_6;
  reg                 io_A_Valid_7_delay_22_5;
  reg                 io_A_Valid_7_delay_23_4;
  reg                 io_A_Valid_7_delay_24_3;
  reg                 io_A_Valid_7_delay_25_2;
  reg                 io_A_Valid_7_delay_26_1;
  reg                 io_A_Valid_7_delay_27;
  reg                 io_B_Valid_27_delay_1_6;
  reg                 io_B_Valid_27_delay_2_5;
  reg                 io_B_Valid_27_delay_3_4;
  reg                 io_B_Valid_27_delay_4_3;
  reg                 io_B_Valid_27_delay_5_2;
  reg                 io_B_Valid_27_delay_6_1;
  reg                 io_B_Valid_27_delay_7;
  reg                 io_A_Valid_7_delay_1_27;
  reg                 io_A_Valid_7_delay_2_26;
  reg                 io_A_Valid_7_delay_3_25;
  reg                 io_A_Valid_7_delay_4_24;
  reg                 io_A_Valid_7_delay_5_23;
  reg                 io_A_Valid_7_delay_6_22;
  reg                 io_A_Valid_7_delay_7_21;
  reg                 io_A_Valid_7_delay_8_20;
  reg                 io_A_Valid_7_delay_9_19;
  reg                 io_A_Valid_7_delay_10_18;
  reg                 io_A_Valid_7_delay_11_17;
  reg                 io_A_Valid_7_delay_12_16;
  reg                 io_A_Valid_7_delay_13_15;
  reg                 io_A_Valid_7_delay_14_14;
  reg                 io_A_Valid_7_delay_15_13;
  reg                 io_A_Valid_7_delay_16_12;
  reg                 io_A_Valid_7_delay_17_11;
  reg                 io_A_Valid_7_delay_18_10;
  reg                 io_A_Valid_7_delay_19_9;
  reg                 io_A_Valid_7_delay_20_8;
  reg                 io_A_Valid_7_delay_21_7;
  reg                 io_A_Valid_7_delay_22_6;
  reg                 io_A_Valid_7_delay_23_5;
  reg                 io_A_Valid_7_delay_24_4;
  reg                 io_A_Valid_7_delay_25_3;
  reg                 io_A_Valid_7_delay_26_2;
  reg                 io_A_Valid_7_delay_27_1;
  reg                 io_A_Valid_7_delay_28;
  reg                 io_B_Valid_28_delay_1_6;
  reg                 io_B_Valid_28_delay_2_5;
  reg                 io_B_Valid_28_delay_3_4;
  reg                 io_B_Valid_28_delay_4_3;
  reg                 io_B_Valid_28_delay_5_2;
  reg                 io_B_Valid_28_delay_6_1;
  reg                 io_B_Valid_28_delay_7;
  reg                 io_A_Valid_7_delay_1_28;
  reg                 io_A_Valid_7_delay_2_27;
  reg                 io_A_Valid_7_delay_3_26;
  reg                 io_A_Valid_7_delay_4_25;
  reg                 io_A_Valid_7_delay_5_24;
  reg                 io_A_Valid_7_delay_6_23;
  reg                 io_A_Valid_7_delay_7_22;
  reg                 io_A_Valid_7_delay_8_21;
  reg                 io_A_Valid_7_delay_9_20;
  reg                 io_A_Valid_7_delay_10_19;
  reg                 io_A_Valid_7_delay_11_18;
  reg                 io_A_Valid_7_delay_12_17;
  reg                 io_A_Valid_7_delay_13_16;
  reg                 io_A_Valid_7_delay_14_15;
  reg                 io_A_Valid_7_delay_15_14;
  reg                 io_A_Valid_7_delay_16_13;
  reg                 io_A_Valid_7_delay_17_12;
  reg                 io_A_Valid_7_delay_18_11;
  reg                 io_A_Valid_7_delay_19_10;
  reg                 io_A_Valid_7_delay_20_9;
  reg                 io_A_Valid_7_delay_21_8;
  reg                 io_A_Valid_7_delay_22_7;
  reg                 io_A_Valid_7_delay_23_6;
  reg                 io_A_Valid_7_delay_24_5;
  reg                 io_A_Valid_7_delay_25_4;
  reg                 io_A_Valid_7_delay_26_3;
  reg                 io_A_Valid_7_delay_27_2;
  reg                 io_A_Valid_7_delay_28_1;
  reg                 io_A_Valid_7_delay_29;
  reg                 io_B_Valid_29_delay_1_6;
  reg                 io_B_Valid_29_delay_2_5;
  reg                 io_B_Valid_29_delay_3_4;
  reg                 io_B_Valid_29_delay_4_3;
  reg                 io_B_Valid_29_delay_5_2;
  reg                 io_B_Valid_29_delay_6_1;
  reg                 io_B_Valid_29_delay_7;
  reg                 io_A_Valid_7_delay_1_29;
  reg                 io_A_Valid_7_delay_2_28;
  reg                 io_A_Valid_7_delay_3_27;
  reg                 io_A_Valid_7_delay_4_26;
  reg                 io_A_Valid_7_delay_5_25;
  reg                 io_A_Valid_7_delay_6_24;
  reg                 io_A_Valid_7_delay_7_23;
  reg                 io_A_Valid_7_delay_8_22;
  reg                 io_A_Valid_7_delay_9_21;
  reg                 io_A_Valid_7_delay_10_20;
  reg                 io_A_Valid_7_delay_11_19;
  reg                 io_A_Valid_7_delay_12_18;
  reg                 io_A_Valid_7_delay_13_17;
  reg                 io_A_Valid_7_delay_14_16;
  reg                 io_A_Valid_7_delay_15_15;
  reg                 io_A_Valid_7_delay_16_14;
  reg                 io_A_Valid_7_delay_17_13;
  reg                 io_A_Valid_7_delay_18_12;
  reg                 io_A_Valid_7_delay_19_11;
  reg                 io_A_Valid_7_delay_20_10;
  reg                 io_A_Valid_7_delay_21_9;
  reg                 io_A_Valid_7_delay_22_8;
  reg                 io_A_Valid_7_delay_23_7;
  reg                 io_A_Valid_7_delay_24_6;
  reg                 io_A_Valid_7_delay_25_5;
  reg                 io_A_Valid_7_delay_26_4;
  reg                 io_A_Valid_7_delay_27_3;
  reg                 io_A_Valid_7_delay_28_2;
  reg                 io_A_Valid_7_delay_29_1;
  reg                 io_A_Valid_7_delay_30;
  reg                 io_B_Valid_30_delay_1_6;
  reg                 io_B_Valid_30_delay_2_5;
  reg                 io_B_Valid_30_delay_3_4;
  reg                 io_B_Valid_30_delay_4_3;
  reg                 io_B_Valid_30_delay_5_2;
  reg                 io_B_Valid_30_delay_6_1;
  reg                 io_B_Valid_30_delay_7;
  reg                 io_A_Valid_7_delay_1_30;
  reg                 io_A_Valid_7_delay_2_29;
  reg                 io_A_Valid_7_delay_3_28;
  reg                 io_A_Valid_7_delay_4_27;
  reg                 io_A_Valid_7_delay_5_26;
  reg                 io_A_Valid_7_delay_6_25;
  reg                 io_A_Valid_7_delay_7_24;
  reg                 io_A_Valid_7_delay_8_23;
  reg                 io_A_Valid_7_delay_9_22;
  reg                 io_A_Valid_7_delay_10_21;
  reg                 io_A_Valid_7_delay_11_20;
  reg                 io_A_Valid_7_delay_12_19;
  reg                 io_A_Valid_7_delay_13_18;
  reg                 io_A_Valid_7_delay_14_17;
  reg                 io_A_Valid_7_delay_15_16;
  reg                 io_A_Valid_7_delay_16_15;
  reg                 io_A_Valid_7_delay_17_14;
  reg                 io_A_Valid_7_delay_18_13;
  reg                 io_A_Valid_7_delay_19_12;
  reg                 io_A_Valid_7_delay_20_11;
  reg                 io_A_Valid_7_delay_21_10;
  reg                 io_A_Valid_7_delay_22_9;
  reg                 io_A_Valid_7_delay_23_8;
  reg                 io_A_Valid_7_delay_24_7;
  reg                 io_A_Valid_7_delay_25_6;
  reg                 io_A_Valid_7_delay_26_5;
  reg                 io_A_Valid_7_delay_27_4;
  reg                 io_A_Valid_7_delay_28_3;
  reg                 io_A_Valid_7_delay_29_2;
  reg                 io_A_Valid_7_delay_30_1;
  reg                 io_A_Valid_7_delay_31;
  reg                 io_B_Valid_31_delay_1_6;
  reg                 io_B_Valid_31_delay_2_5;
  reg                 io_B_Valid_31_delay_3_4;
  reg                 io_B_Valid_31_delay_4_3;
  reg                 io_B_Valid_31_delay_5_2;
  reg                 io_B_Valid_31_delay_6_1;
  reg                 io_B_Valid_31_delay_7;
  reg                 io_A_Valid_7_delay_1_31;
  reg                 io_A_Valid_7_delay_2_30;
  reg                 io_A_Valid_7_delay_3_29;
  reg                 io_A_Valid_7_delay_4_28;
  reg                 io_A_Valid_7_delay_5_27;
  reg                 io_A_Valid_7_delay_6_26;
  reg                 io_A_Valid_7_delay_7_25;
  reg                 io_A_Valid_7_delay_8_24;
  reg                 io_A_Valid_7_delay_9_23;
  reg                 io_A_Valid_7_delay_10_22;
  reg                 io_A_Valid_7_delay_11_21;
  reg                 io_A_Valid_7_delay_12_20;
  reg                 io_A_Valid_7_delay_13_19;
  reg                 io_A_Valid_7_delay_14_18;
  reg                 io_A_Valid_7_delay_15_17;
  reg                 io_A_Valid_7_delay_16_16;
  reg                 io_A_Valid_7_delay_17_15;
  reg                 io_A_Valid_7_delay_18_14;
  reg                 io_A_Valid_7_delay_19_13;
  reg                 io_A_Valid_7_delay_20_12;
  reg                 io_A_Valid_7_delay_21_11;
  reg                 io_A_Valid_7_delay_22_10;
  reg                 io_A_Valid_7_delay_23_9;
  reg                 io_A_Valid_7_delay_24_8;
  reg                 io_A_Valid_7_delay_25_7;
  reg                 io_A_Valid_7_delay_26_6;
  reg                 io_A_Valid_7_delay_27_5;
  reg                 io_A_Valid_7_delay_28_4;
  reg                 io_A_Valid_7_delay_29_3;
  reg                 io_A_Valid_7_delay_30_2;
  reg                 io_A_Valid_7_delay_31_1;
  reg                 io_A_Valid_7_delay_32;
  reg                 io_B_Valid_32_delay_1_6;
  reg                 io_B_Valid_32_delay_2_5;
  reg                 io_B_Valid_32_delay_3_4;
  reg                 io_B_Valid_32_delay_4_3;
  reg                 io_B_Valid_32_delay_5_2;
  reg                 io_B_Valid_32_delay_6_1;
  reg                 io_B_Valid_32_delay_7;
  reg                 io_A_Valid_7_delay_1_32;
  reg                 io_A_Valid_7_delay_2_31;
  reg                 io_A_Valid_7_delay_3_30;
  reg                 io_A_Valid_7_delay_4_29;
  reg                 io_A_Valid_7_delay_5_28;
  reg                 io_A_Valid_7_delay_6_27;
  reg                 io_A_Valid_7_delay_7_26;
  reg                 io_A_Valid_7_delay_8_25;
  reg                 io_A_Valid_7_delay_9_24;
  reg                 io_A_Valid_7_delay_10_23;
  reg                 io_A_Valid_7_delay_11_22;
  reg                 io_A_Valid_7_delay_12_21;
  reg                 io_A_Valid_7_delay_13_20;
  reg                 io_A_Valid_7_delay_14_19;
  reg                 io_A_Valid_7_delay_15_18;
  reg                 io_A_Valid_7_delay_16_17;
  reg                 io_A_Valid_7_delay_17_16;
  reg                 io_A_Valid_7_delay_18_15;
  reg                 io_A_Valid_7_delay_19_14;
  reg                 io_A_Valid_7_delay_20_13;
  reg                 io_A_Valid_7_delay_21_12;
  reg                 io_A_Valid_7_delay_22_11;
  reg                 io_A_Valid_7_delay_23_10;
  reg                 io_A_Valid_7_delay_24_9;
  reg                 io_A_Valid_7_delay_25_8;
  reg                 io_A_Valid_7_delay_26_7;
  reg                 io_A_Valid_7_delay_27_6;
  reg                 io_A_Valid_7_delay_28_5;
  reg                 io_A_Valid_7_delay_29_4;
  reg                 io_A_Valid_7_delay_30_3;
  reg                 io_A_Valid_7_delay_31_2;
  reg                 io_A_Valid_7_delay_32_1;
  reg                 io_A_Valid_7_delay_33;
  reg                 io_B_Valid_33_delay_1_6;
  reg                 io_B_Valid_33_delay_2_5;
  reg                 io_B_Valid_33_delay_3_4;
  reg                 io_B_Valid_33_delay_4_3;
  reg                 io_B_Valid_33_delay_5_2;
  reg                 io_B_Valid_33_delay_6_1;
  reg                 io_B_Valid_33_delay_7;
  reg                 io_A_Valid_7_delay_1_33;
  reg                 io_A_Valid_7_delay_2_32;
  reg                 io_A_Valid_7_delay_3_31;
  reg                 io_A_Valid_7_delay_4_30;
  reg                 io_A_Valid_7_delay_5_29;
  reg                 io_A_Valid_7_delay_6_28;
  reg                 io_A_Valid_7_delay_7_27;
  reg                 io_A_Valid_7_delay_8_26;
  reg                 io_A_Valid_7_delay_9_25;
  reg                 io_A_Valid_7_delay_10_24;
  reg                 io_A_Valid_7_delay_11_23;
  reg                 io_A_Valid_7_delay_12_22;
  reg                 io_A_Valid_7_delay_13_21;
  reg                 io_A_Valid_7_delay_14_20;
  reg                 io_A_Valid_7_delay_15_19;
  reg                 io_A_Valid_7_delay_16_18;
  reg                 io_A_Valid_7_delay_17_17;
  reg                 io_A_Valid_7_delay_18_16;
  reg                 io_A_Valid_7_delay_19_15;
  reg                 io_A_Valid_7_delay_20_14;
  reg                 io_A_Valid_7_delay_21_13;
  reg                 io_A_Valid_7_delay_22_12;
  reg                 io_A_Valid_7_delay_23_11;
  reg                 io_A_Valid_7_delay_24_10;
  reg                 io_A_Valid_7_delay_25_9;
  reg                 io_A_Valid_7_delay_26_8;
  reg                 io_A_Valid_7_delay_27_7;
  reg                 io_A_Valid_7_delay_28_6;
  reg                 io_A_Valid_7_delay_29_5;
  reg                 io_A_Valid_7_delay_30_4;
  reg                 io_A_Valid_7_delay_31_3;
  reg                 io_A_Valid_7_delay_32_2;
  reg                 io_A_Valid_7_delay_33_1;
  reg                 io_A_Valid_7_delay_34;
  reg                 io_B_Valid_34_delay_1_6;
  reg                 io_B_Valid_34_delay_2_5;
  reg                 io_B_Valid_34_delay_3_4;
  reg                 io_B_Valid_34_delay_4_3;
  reg                 io_B_Valid_34_delay_5_2;
  reg                 io_B_Valid_34_delay_6_1;
  reg                 io_B_Valid_34_delay_7;
  reg                 io_A_Valid_7_delay_1_34;
  reg                 io_A_Valid_7_delay_2_33;
  reg                 io_A_Valid_7_delay_3_32;
  reg                 io_A_Valid_7_delay_4_31;
  reg                 io_A_Valid_7_delay_5_30;
  reg                 io_A_Valid_7_delay_6_29;
  reg                 io_A_Valid_7_delay_7_28;
  reg                 io_A_Valid_7_delay_8_27;
  reg                 io_A_Valid_7_delay_9_26;
  reg                 io_A_Valid_7_delay_10_25;
  reg                 io_A_Valid_7_delay_11_24;
  reg                 io_A_Valid_7_delay_12_23;
  reg                 io_A_Valid_7_delay_13_22;
  reg                 io_A_Valid_7_delay_14_21;
  reg                 io_A_Valid_7_delay_15_20;
  reg                 io_A_Valid_7_delay_16_19;
  reg                 io_A_Valid_7_delay_17_18;
  reg                 io_A_Valid_7_delay_18_17;
  reg                 io_A_Valid_7_delay_19_16;
  reg                 io_A_Valid_7_delay_20_15;
  reg                 io_A_Valid_7_delay_21_14;
  reg                 io_A_Valid_7_delay_22_13;
  reg                 io_A_Valid_7_delay_23_12;
  reg                 io_A_Valid_7_delay_24_11;
  reg                 io_A_Valid_7_delay_25_10;
  reg                 io_A_Valid_7_delay_26_9;
  reg                 io_A_Valid_7_delay_27_8;
  reg                 io_A_Valid_7_delay_28_7;
  reg                 io_A_Valid_7_delay_29_6;
  reg                 io_A_Valid_7_delay_30_5;
  reg                 io_A_Valid_7_delay_31_4;
  reg                 io_A_Valid_7_delay_32_3;
  reg                 io_A_Valid_7_delay_33_2;
  reg                 io_A_Valid_7_delay_34_1;
  reg                 io_A_Valid_7_delay_35;
  reg                 io_B_Valid_35_delay_1_6;
  reg                 io_B_Valid_35_delay_2_5;
  reg                 io_B_Valid_35_delay_3_4;
  reg                 io_B_Valid_35_delay_4_3;
  reg                 io_B_Valid_35_delay_5_2;
  reg                 io_B_Valid_35_delay_6_1;
  reg                 io_B_Valid_35_delay_7;
  reg                 io_A_Valid_7_delay_1_35;
  reg                 io_A_Valid_7_delay_2_34;
  reg                 io_A_Valid_7_delay_3_33;
  reg                 io_A_Valid_7_delay_4_32;
  reg                 io_A_Valid_7_delay_5_31;
  reg                 io_A_Valid_7_delay_6_30;
  reg                 io_A_Valid_7_delay_7_29;
  reg                 io_A_Valid_7_delay_8_28;
  reg                 io_A_Valid_7_delay_9_27;
  reg                 io_A_Valid_7_delay_10_26;
  reg                 io_A_Valid_7_delay_11_25;
  reg                 io_A_Valid_7_delay_12_24;
  reg                 io_A_Valid_7_delay_13_23;
  reg                 io_A_Valid_7_delay_14_22;
  reg                 io_A_Valid_7_delay_15_21;
  reg                 io_A_Valid_7_delay_16_20;
  reg                 io_A_Valid_7_delay_17_19;
  reg                 io_A_Valid_7_delay_18_18;
  reg                 io_A_Valid_7_delay_19_17;
  reg                 io_A_Valid_7_delay_20_16;
  reg                 io_A_Valid_7_delay_21_15;
  reg                 io_A_Valid_7_delay_22_14;
  reg                 io_A_Valid_7_delay_23_13;
  reg                 io_A_Valid_7_delay_24_12;
  reg                 io_A_Valid_7_delay_25_11;
  reg                 io_A_Valid_7_delay_26_10;
  reg                 io_A_Valid_7_delay_27_9;
  reg                 io_A_Valid_7_delay_28_8;
  reg                 io_A_Valid_7_delay_29_7;
  reg                 io_A_Valid_7_delay_30_6;
  reg                 io_A_Valid_7_delay_31_5;
  reg                 io_A_Valid_7_delay_32_4;
  reg                 io_A_Valid_7_delay_33_3;
  reg                 io_A_Valid_7_delay_34_2;
  reg                 io_A_Valid_7_delay_35_1;
  reg                 io_A_Valid_7_delay_36;
  reg                 io_B_Valid_36_delay_1_6;
  reg                 io_B_Valid_36_delay_2_5;
  reg                 io_B_Valid_36_delay_3_4;
  reg                 io_B_Valid_36_delay_4_3;
  reg                 io_B_Valid_36_delay_5_2;
  reg                 io_B_Valid_36_delay_6_1;
  reg                 io_B_Valid_36_delay_7;
  reg                 io_A_Valid_7_delay_1_36;
  reg                 io_A_Valid_7_delay_2_35;
  reg                 io_A_Valid_7_delay_3_34;
  reg                 io_A_Valid_7_delay_4_33;
  reg                 io_A_Valid_7_delay_5_32;
  reg                 io_A_Valid_7_delay_6_31;
  reg                 io_A_Valid_7_delay_7_30;
  reg                 io_A_Valid_7_delay_8_29;
  reg                 io_A_Valid_7_delay_9_28;
  reg                 io_A_Valid_7_delay_10_27;
  reg                 io_A_Valid_7_delay_11_26;
  reg                 io_A_Valid_7_delay_12_25;
  reg                 io_A_Valid_7_delay_13_24;
  reg                 io_A_Valid_7_delay_14_23;
  reg                 io_A_Valid_7_delay_15_22;
  reg                 io_A_Valid_7_delay_16_21;
  reg                 io_A_Valid_7_delay_17_20;
  reg                 io_A_Valid_7_delay_18_19;
  reg                 io_A_Valid_7_delay_19_18;
  reg                 io_A_Valid_7_delay_20_17;
  reg                 io_A_Valid_7_delay_21_16;
  reg                 io_A_Valid_7_delay_22_15;
  reg                 io_A_Valid_7_delay_23_14;
  reg                 io_A_Valid_7_delay_24_13;
  reg                 io_A_Valid_7_delay_25_12;
  reg                 io_A_Valid_7_delay_26_11;
  reg                 io_A_Valid_7_delay_27_10;
  reg                 io_A_Valid_7_delay_28_9;
  reg                 io_A_Valid_7_delay_29_8;
  reg                 io_A_Valid_7_delay_30_7;
  reg                 io_A_Valid_7_delay_31_6;
  reg                 io_A_Valid_7_delay_32_5;
  reg                 io_A_Valid_7_delay_33_4;
  reg                 io_A_Valid_7_delay_34_3;
  reg                 io_A_Valid_7_delay_35_2;
  reg                 io_A_Valid_7_delay_36_1;
  reg                 io_A_Valid_7_delay_37;
  reg                 io_B_Valid_37_delay_1_6;
  reg                 io_B_Valid_37_delay_2_5;
  reg                 io_B_Valid_37_delay_3_4;
  reg                 io_B_Valid_37_delay_4_3;
  reg                 io_B_Valid_37_delay_5_2;
  reg                 io_B_Valid_37_delay_6_1;
  reg                 io_B_Valid_37_delay_7;
  reg                 io_A_Valid_7_delay_1_37;
  reg                 io_A_Valid_7_delay_2_36;
  reg                 io_A_Valid_7_delay_3_35;
  reg                 io_A_Valid_7_delay_4_34;
  reg                 io_A_Valid_7_delay_5_33;
  reg                 io_A_Valid_7_delay_6_32;
  reg                 io_A_Valid_7_delay_7_31;
  reg                 io_A_Valid_7_delay_8_30;
  reg                 io_A_Valid_7_delay_9_29;
  reg                 io_A_Valid_7_delay_10_28;
  reg                 io_A_Valid_7_delay_11_27;
  reg                 io_A_Valid_7_delay_12_26;
  reg                 io_A_Valid_7_delay_13_25;
  reg                 io_A_Valid_7_delay_14_24;
  reg                 io_A_Valid_7_delay_15_23;
  reg                 io_A_Valid_7_delay_16_22;
  reg                 io_A_Valid_7_delay_17_21;
  reg                 io_A_Valid_7_delay_18_20;
  reg                 io_A_Valid_7_delay_19_19;
  reg                 io_A_Valid_7_delay_20_18;
  reg                 io_A_Valid_7_delay_21_17;
  reg                 io_A_Valid_7_delay_22_16;
  reg                 io_A_Valid_7_delay_23_15;
  reg                 io_A_Valid_7_delay_24_14;
  reg                 io_A_Valid_7_delay_25_13;
  reg                 io_A_Valid_7_delay_26_12;
  reg                 io_A_Valid_7_delay_27_11;
  reg                 io_A_Valid_7_delay_28_10;
  reg                 io_A_Valid_7_delay_29_9;
  reg                 io_A_Valid_7_delay_30_8;
  reg                 io_A_Valid_7_delay_31_7;
  reg                 io_A_Valid_7_delay_32_6;
  reg                 io_A_Valid_7_delay_33_5;
  reg                 io_A_Valid_7_delay_34_4;
  reg                 io_A_Valid_7_delay_35_3;
  reg                 io_A_Valid_7_delay_36_2;
  reg                 io_A_Valid_7_delay_37_1;
  reg                 io_A_Valid_7_delay_38;
  reg                 io_B_Valid_38_delay_1_6;
  reg                 io_B_Valid_38_delay_2_5;
  reg                 io_B_Valid_38_delay_3_4;
  reg                 io_B_Valid_38_delay_4_3;
  reg                 io_B_Valid_38_delay_5_2;
  reg                 io_B_Valid_38_delay_6_1;
  reg                 io_B_Valid_38_delay_7;
  reg                 io_A_Valid_7_delay_1_38;
  reg                 io_A_Valid_7_delay_2_37;
  reg                 io_A_Valid_7_delay_3_36;
  reg                 io_A_Valid_7_delay_4_35;
  reg                 io_A_Valid_7_delay_5_34;
  reg                 io_A_Valid_7_delay_6_33;
  reg                 io_A_Valid_7_delay_7_32;
  reg                 io_A_Valid_7_delay_8_31;
  reg                 io_A_Valid_7_delay_9_30;
  reg                 io_A_Valid_7_delay_10_29;
  reg                 io_A_Valid_7_delay_11_28;
  reg                 io_A_Valid_7_delay_12_27;
  reg                 io_A_Valid_7_delay_13_26;
  reg                 io_A_Valid_7_delay_14_25;
  reg                 io_A_Valid_7_delay_15_24;
  reg                 io_A_Valid_7_delay_16_23;
  reg                 io_A_Valid_7_delay_17_22;
  reg                 io_A_Valid_7_delay_18_21;
  reg                 io_A_Valid_7_delay_19_20;
  reg                 io_A_Valid_7_delay_20_19;
  reg                 io_A_Valid_7_delay_21_18;
  reg                 io_A_Valid_7_delay_22_17;
  reg                 io_A_Valid_7_delay_23_16;
  reg                 io_A_Valid_7_delay_24_15;
  reg                 io_A_Valid_7_delay_25_14;
  reg                 io_A_Valid_7_delay_26_13;
  reg                 io_A_Valid_7_delay_27_12;
  reg                 io_A_Valid_7_delay_28_11;
  reg                 io_A_Valid_7_delay_29_10;
  reg                 io_A_Valid_7_delay_30_9;
  reg                 io_A_Valid_7_delay_31_8;
  reg                 io_A_Valid_7_delay_32_7;
  reg                 io_A_Valid_7_delay_33_6;
  reg                 io_A_Valid_7_delay_34_5;
  reg                 io_A_Valid_7_delay_35_4;
  reg                 io_A_Valid_7_delay_36_3;
  reg                 io_A_Valid_7_delay_37_2;
  reg                 io_A_Valid_7_delay_38_1;
  reg                 io_A_Valid_7_delay_39;
  reg                 io_B_Valid_39_delay_1_6;
  reg                 io_B_Valid_39_delay_2_5;
  reg                 io_B_Valid_39_delay_3_4;
  reg                 io_B_Valid_39_delay_4_3;
  reg                 io_B_Valid_39_delay_5_2;
  reg                 io_B_Valid_39_delay_6_1;
  reg                 io_B_Valid_39_delay_7;
  reg                 io_A_Valid_7_delay_1_39;
  reg                 io_A_Valid_7_delay_2_38;
  reg                 io_A_Valid_7_delay_3_37;
  reg                 io_A_Valid_7_delay_4_36;
  reg                 io_A_Valid_7_delay_5_35;
  reg                 io_A_Valid_7_delay_6_34;
  reg                 io_A_Valid_7_delay_7_33;
  reg                 io_A_Valid_7_delay_8_32;
  reg                 io_A_Valid_7_delay_9_31;
  reg                 io_A_Valid_7_delay_10_30;
  reg                 io_A_Valid_7_delay_11_29;
  reg                 io_A_Valid_7_delay_12_28;
  reg                 io_A_Valid_7_delay_13_27;
  reg                 io_A_Valid_7_delay_14_26;
  reg                 io_A_Valid_7_delay_15_25;
  reg                 io_A_Valid_7_delay_16_24;
  reg                 io_A_Valid_7_delay_17_23;
  reg                 io_A_Valid_7_delay_18_22;
  reg                 io_A_Valid_7_delay_19_21;
  reg                 io_A_Valid_7_delay_20_20;
  reg                 io_A_Valid_7_delay_21_19;
  reg                 io_A_Valid_7_delay_22_18;
  reg                 io_A_Valid_7_delay_23_17;
  reg                 io_A_Valid_7_delay_24_16;
  reg                 io_A_Valid_7_delay_25_15;
  reg                 io_A_Valid_7_delay_26_14;
  reg                 io_A_Valid_7_delay_27_13;
  reg                 io_A_Valid_7_delay_28_12;
  reg                 io_A_Valid_7_delay_29_11;
  reg                 io_A_Valid_7_delay_30_10;
  reg                 io_A_Valid_7_delay_31_9;
  reg                 io_A_Valid_7_delay_32_8;
  reg                 io_A_Valid_7_delay_33_7;
  reg                 io_A_Valid_7_delay_34_6;
  reg                 io_A_Valid_7_delay_35_5;
  reg                 io_A_Valid_7_delay_36_4;
  reg                 io_A_Valid_7_delay_37_3;
  reg                 io_A_Valid_7_delay_38_2;
  reg                 io_A_Valid_7_delay_39_1;
  reg                 io_A_Valid_7_delay_40;
  reg                 io_B_Valid_40_delay_1_6;
  reg                 io_B_Valid_40_delay_2_5;
  reg                 io_B_Valid_40_delay_3_4;
  reg                 io_B_Valid_40_delay_4_3;
  reg                 io_B_Valid_40_delay_5_2;
  reg                 io_B_Valid_40_delay_6_1;
  reg                 io_B_Valid_40_delay_7;
  reg                 io_A_Valid_7_delay_1_40;
  reg                 io_A_Valid_7_delay_2_39;
  reg                 io_A_Valid_7_delay_3_38;
  reg                 io_A_Valid_7_delay_4_37;
  reg                 io_A_Valid_7_delay_5_36;
  reg                 io_A_Valid_7_delay_6_35;
  reg                 io_A_Valid_7_delay_7_34;
  reg                 io_A_Valid_7_delay_8_33;
  reg                 io_A_Valid_7_delay_9_32;
  reg                 io_A_Valid_7_delay_10_31;
  reg                 io_A_Valid_7_delay_11_30;
  reg                 io_A_Valid_7_delay_12_29;
  reg                 io_A_Valid_7_delay_13_28;
  reg                 io_A_Valid_7_delay_14_27;
  reg                 io_A_Valid_7_delay_15_26;
  reg                 io_A_Valid_7_delay_16_25;
  reg                 io_A_Valid_7_delay_17_24;
  reg                 io_A_Valid_7_delay_18_23;
  reg                 io_A_Valid_7_delay_19_22;
  reg                 io_A_Valid_7_delay_20_21;
  reg                 io_A_Valid_7_delay_21_20;
  reg                 io_A_Valid_7_delay_22_19;
  reg                 io_A_Valid_7_delay_23_18;
  reg                 io_A_Valid_7_delay_24_17;
  reg                 io_A_Valid_7_delay_25_16;
  reg                 io_A_Valid_7_delay_26_15;
  reg                 io_A_Valid_7_delay_27_14;
  reg                 io_A_Valid_7_delay_28_13;
  reg                 io_A_Valid_7_delay_29_12;
  reg                 io_A_Valid_7_delay_30_11;
  reg                 io_A_Valid_7_delay_31_10;
  reg                 io_A_Valid_7_delay_32_9;
  reg                 io_A_Valid_7_delay_33_8;
  reg                 io_A_Valid_7_delay_34_7;
  reg                 io_A_Valid_7_delay_35_6;
  reg                 io_A_Valid_7_delay_36_5;
  reg                 io_A_Valid_7_delay_37_4;
  reg                 io_A_Valid_7_delay_38_3;
  reg                 io_A_Valid_7_delay_39_2;
  reg                 io_A_Valid_7_delay_40_1;
  reg                 io_A_Valid_7_delay_41;
  reg                 io_B_Valid_41_delay_1_6;
  reg                 io_B_Valid_41_delay_2_5;
  reg                 io_B_Valid_41_delay_3_4;
  reg                 io_B_Valid_41_delay_4_3;
  reg                 io_B_Valid_41_delay_5_2;
  reg                 io_B_Valid_41_delay_6_1;
  reg                 io_B_Valid_41_delay_7;
  reg                 io_A_Valid_7_delay_1_41;
  reg                 io_A_Valid_7_delay_2_40;
  reg                 io_A_Valid_7_delay_3_39;
  reg                 io_A_Valid_7_delay_4_38;
  reg                 io_A_Valid_7_delay_5_37;
  reg                 io_A_Valid_7_delay_6_36;
  reg                 io_A_Valid_7_delay_7_35;
  reg                 io_A_Valid_7_delay_8_34;
  reg                 io_A_Valid_7_delay_9_33;
  reg                 io_A_Valid_7_delay_10_32;
  reg                 io_A_Valid_7_delay_11_31;
  reg                 io_A_Valid_7_delay_12_30;
  reg                 io_A_Valid_7_delay_13_29;
  reg                 io_A_Valid_7_delay_14_28;
  reg                 io_A_Valid_7_delay_15_27;
  reg                 io_A_Valid_7_delay_16_26;
  reg                 io_A_Valid_7_delay_17_25;
  reg                 io_A_Valid_7_delay_18_24;
  reg                 io_A_Valid_7_delay_19_23;
  reg                 io_A_Valid_7_delay_20_22;
  reg                 io_A_Valid_7_delay_21_21;
  reg                 io_A_Valid_7_delay_22_20;
  reg                 io_A_Valid_7_delay_23_19;
  reg                 io_A_Valid_7_delay_24_18;
  reg                 io_A_Valid_7_delay_25_17;
  reg                 io_A_Valid_7_delay_26_16;
  reg                 io_A_Valid_7_delay_27_15;
  reg                 io_A_Valid_7_delay_28_14;
  reg                 io_A_Valid_7_delay_29_13;
  reg                 io_A_Valid_7_delay_30_12;
  reg                 io_A_Valid_7_delay_31_11;
  reg                 io_A_Valid_7_delay_32_10;
  reg                 io_A_Valid_7_delay_33_9;
  reg                 io_A_Valid_7_delay_34_8;
  reg                 io_A_Valid_7_delay_35_7;
  reg                 io_A_Valid_7_delay_36_6;
  reg                 io_A_Valid_7_delay_37_5;
  reg                 io_A_Valid_7_delay_38_4;
  reg                 io_A_Valid_7_delay_39_3;
  reg                 io_A_Valid_7_delay_40_2;
  reg                 io_A_Valid_7_delay_41_1;
  reg                 io_A_Valid_7_delay_42;
  reg                 io_B_Valid_42_delay_1_6;
  reg                 io_B_Valid_42_delay_2_5;
  reg                 io_B_Valid_42_delay_3_4;
  reg                 io_B_Valid_42_delay_4_3;
  reg                 io_B_Valid_42_delay_5_2;
  reg                 io_B_Valid_42_delay_6_1;
  reg                 io_B_Valid_42_delay_7;
  reg                 io_A_Valid_7_delay_1_42;
  reg                 io_A_Valid_7_delay_2_41;
  reg                 io_A_Valid_7_delay_3_40;
  reg                 io_A_Valid_7_delay_4_39;
  reg                 io_A_Valid_7_delay_5_38;
  reg                 io_A_Valid_7_delay_6_37;
  reg                 io_A_Valid_7_delay_7_36;
  reg                 io_A_Valid_7_delay_8_35;
  reg                 io_A_Valid_7_delay_9_34;
  reg                 io_A_Valid_7_delay_10_33;
  reg                 io_A_Valid_7_delay_11_32;
  reg                 io_A_Valid_7_delay_12_31;
  reg                 io_A_Valid_7_delay_13_30;
  reg                 io_A_Valid_7_delay_14_29;
  reg                 io_A_Valid_7_delay_15_28;
  reg                 io_A_Valid_7_delay_16_27;
  reg                 io_A_Valid_7_delay_17_26;
  reg                 io_A_Valid_7_delay_18_25;
  reg                 io_A_Valid_7_delay_19_24;
  reg                 io_A_Valid_7_delay_20_23;
  reg                 io_A_Valid_7_delay_21_22;
  reg                 io_A_Valid_7_delay_22_21;
  reg                 io_A_Valid_7_delay_23_20;
  reg                 io_A_Valid_7_delay_24_19;
  reg                 io_A_Valid_7_delay_25_18;
  reg                 io_A_Valid_7_delay_26_17;
  reg                 io_A_Valid_7_delay_27_16;
  reg                 io_A_Valid_7_delay_28_15;
  reg                 io_A_Valid_7_delay_29_14;
  reg                 io_A_Valid_7_delay_30_13;
  reg                 io_A_Valid_7_delay_31_12;
  reg                 io_A_Valid_7_delay_32_11;
  reg                 io_A_Valid_7_delay_33_10;
  reg                 io_A_Valid_7_delay_34_9;
  reg                 io_A_Valid_7_delay_35_8;
  reg                 io_A_Valid_7_delay_36_7;
  reg                 io_A_Valid_7_delay_37_6;
  reg                 io_A_Valid_7_delay_38_5;
  reg                 io_A_Valid_7_delay_39_4;
  reg                 io_A_Valid_7_delay_40_3;
  reg                 io_A_Valid_7_delay_41_2;
  reg                 io_A_Valid_7_delay_42_1;
  reg                 io_A_Valid_7_delay_43;
  reg                 io_B_Valid_43_delay_1_6;
  reg                 io_B_Valid_43_delay_2_5;
  reg                 io_B_Valid_43_delay_3_4;
  reg                 io_B_Valid_43_delay_4_3;
  reg                 io_B_Valid_43_delay_5_2;
  reg                 io_B_Valid_43_delay_6_1;
  reg                 io_B_Valid_43_delay_7;
  reg                 io_A_Valid_7_delay_1_43;
  reg                 io_A_Valid_7_delay_2_42;
  reg                 io_A_Valid_7_delay_3_41;
  reg                 io_A_Valid_7_delay_4_40;
  reg                 io_A_Valid_7_delay_5_39;
  reg                 io_A_Valid_7_delay_6_38;
  reg                 io_A_Valid_7_delay_7_37;
  reg                 io_A_Valid_7_delay_8_36;
  reg                 io_A_Valid_7_delay_9_35;
  reg                 io_A_Valid_7_delay_10_34;
  reg                 io_A_Valid_7_delay_11_33;
  reg                 io_A_Valid_7_delay_12_32;
  reg                 io_A_Valid_7_delay_13_31;
  reg                 io_A_Valid_7_delay_14_30;
  reg                 io_A_Valid_7_delay_15_29;
  reg                 io_A_Valid_7_delay_16_28;
  reg                 io_A_Valid_7_delay_17_27;
  reg                 io_A_Valid_7_delay_18_26;
  reg                 io_A_Valid_7_delay_19_25;
  reg                 io_A_Valid_7_delay_20_24;
  reg                 io_A_Valid_7_delay_21_23;
  reg                 io_A_Valid_7_delay_22_22;
  reg                 io_A_Valid_7_delay_23_21;
  reg                 io_A_Valid_7_delay_24_20;
  reg                 io_A_Valid_7_delay_25_19;
  reg                 io_A_Valid_7_delay_26_18;
  reg                 io_A_Valid_7_delay_27_17;
  reg                 io_A_Valid_7_delay_28_16;
  reg                 io_A_Valid_7_delay_29_15;
  reg                 io_A_Valid_7_delay_30_14;
  reg                 io_A_Valid_7_delay_31_13;
  reg                 io_A_Valid_7_delay_32_12;
  reg                 io_A_Valid_7_delay_33_11;
  reg                 io_A_Valid_7_delay_34_10;
  reg                 io_A_Valid_7_delay_35_9;
  reg                 io_A_Valid_7_delay_36_8;
  reg                 io_A_Valid_7_delay_37_7;
  reg                 io_A_Valid_7_delay_38_6;
  reg                 io_A_Valid_7_delay_39_5;
  reg                 io_A_Valid_7_delay_40_4;
  reg                 io_A_Valid_7_delay_41_3;
  reg                 io_A_Valid_7_delay_42_2;
  reg                 io_A_Valid_7_delay_43_1;
  reg                 io_A_Valid_7_delay_44;
  reg                 io_B_Valid_44_delay_1_6;
  reg                 io_B_Valid_44_delay_2_5;
  reg                 io_B_Valid_44_delay_3_4;
  reg                 io_B_Valid_44_delay_4_3;
  reg                 io_B_Valid_44_delay_5_2;
  reg                 io_B_Valid_44_delay_6_1;
  reg                 io_B_Valid_44_delay_7;
  reg                 io_A_Valid_7_delay_1_44;
  reg                 io_A_Valid_7_delay_2_43;
  reg                 io_A_Valid_7_delay_3_42;
  reg                 io_A_Valid_7_delay_4_41;
  reg                 io_A_Valid_7_delay_5_40;
  reg                 io_A_Valid_7_delay_6_39;
  reg                 io_A_Valid_7_delay_7_38;
  reg                 io_A_Valid_7_delay_8_37;
  reg                 io_A_Valid_7_delay_9_36;
  reg                 io_A_Valid_7_delay_10_35;
  reg                 io_A_Valid_7_delay_11_34;
  reg                 io_A_Valid_7_delay_12_33;
  reg                 io_A_Valid_7_delay_13_32;
  reg                 io_A_Valid_7_delay_14_31;
  reg                 io_A_Valid_7_delay_15_30;
  reg                 io_A_Valid_7_delay_16_29;
  reg                 io_A_Valid_7_delay_17_28;
  reg                 io_A_Valid_7_delay_18_27;
  reg                 io_A_Valid_7_delay_19_26;
  reg                 io_A_Valid_7_delay_20_25;
  reg                 io_A_Valid_7_delay_21_24;
  reg                 io_A_Valid_7_delay_22_23;
  reg                 io_A_Valid_7_delay_23_22;
  reg                 io_A_Valid_7_delay_24_21;
  reg                 io_A_Valid_7_delay_25_20;
  reg                 io_A_Valid_7_delay_26_19;
  reg                 io_A_Valid_7_delay_27_18;
  reg                 io_A_Valid_7_delay_28_17;
  reg                 io_A_Valid_7_delay_29_16;
  reg                 io_A_Valid_7_delay_30_15;
  reg                 io_A_Valid_7_delay_31_14;
  reg                 io_A_Valid_7_delay_32_13;
  reg                 io_A_Valid_7_delay_33_12;
  reg                 io_A_Valid_7_delay_34_11;
  reg                 io_A_Valid_7_delay_35_10;
  reg                 io_A_Valid_7_delay_36_9;
  reg                 io_A_Valid_7_delay_37_8;
  reg                 io_A_Valid_7_delay_38_7;
  reg                 io_A_Valid_7_delay_39_6;
  reg                 io_A_Valid_7_delay_40_5;
  reg                 io_A_Valid_7_delay_41_4;
  reg                 io_A_Valid_7_delay_42_3;
  reg                 io_A_Valid_7_delay_43_2;
  reg                 io_A_Valid_7_delay_44_1;
  reg                 io_A_Valid_7_delay_45;
  reg                 io_B_Valid_45_delay_1_6;
  reg                 io_B_Valid_45_delay_2_5;
  reg                 io_B_Valid_45_delay_3_4;
  reg                 io_B_Valid_45_delay_4_3;
  reg                 io_B_Valid_45_delay_5_2;
  reg                 io_B_Valid_45_delay_6_1;
  reg                 io_B_Valid_45_delay_7;
  reg                 io_A_Valid_7_delay_1_45;
  reg                 io_A_Valid_7_delay_2_44;
  reg                 io_A_Valid_7_delay_3_43;
  reg                 io_A_Valid_7_delay_4_42;
  reg                 io_A_Valid_7_delay_5_41;
  reg                 io_A_Valid_7_delay_6_40;
  reg                 io_A_Valid_7_delay_7_39;
  reg                 io_A_Valid_7_delay_8_38;
  reg                 io_A_Valid_7_delay_9_37;
  reg                 io_A_Valid_7_delay_10_36;
  reg                 io_A_Valid_7_delay_11_35;
  reg                 io_A_Valid_7_delay_12_34;
  reg                 io_A_Valid_7_delay_13_33;
  reg                 io_A_Valid_7_delay_14_32;
  reg                 io_A_Valid_7_delay_15_31;
  reg                 io_A_Valid_7_delay_16_30;
  reg                 io_A_Valid_7_delay_17_29;
  reg                 io_A_Valid_7_delay_18_28;
  reg                 io_A_Valid_7_delay_19_27;
  reg                 io_A_Valid_7_delay_20_26;
  reg                 io_A_Valid_7_delay_21_25;
  reg                 io_A_Valid_7_delay_22_24;
  reg                 io_A_Valid_7_delay_23_23;
  reg                 io_A_Valid_7_delay_24_22;
  reg                 io_A_Valid_7_delay_25_21;
  reg                 io_A_Valid_7_delay_26_20;
  reg                 io_A_Valid_7_delay_27_19;
  reg                 io_A_Valid_7_delay_28_18;
  reg                 io_A_Valid_7_delay_29_17;
  reg                 io_A_Valid_7_delay_30_16;
  reg                 io_A_Valid_7_delay_31_15;
  reg                 io_A_Valid_7_delay_32_14;
  reg                 io_A_Valid_7_delay_33_13;
  reg                 io_A_Valid_7_delay_34_12;
  reg                 io_A_Valid_7_delay_35_11;
  reg                 io_A_Valid_7_delay_36_10;
  reg                 io_A_Valid_7_delay_37_9;
  reg                 io_A_Valid_7_delay_38_8;
  reg                 io_A_Valid_7_delay_39_7;
  reg                 io_A_Valid_7_delay_40_6;
  reg                 io_A_Valid_7_delay_41_5;
  reg                 io_A_Valid_7_delay_42_4;
  reg                 io_A_Valid_7_delay_43_3;
  reg                 io_A_Valid_7_delay_44_2;
  reg                 io_A_Valid_7_delay_45_1;
  reg                 io_A_Valid_7_delay_46;
  reg                 io_B_Valid_46_delay_1_6;
  reg                 io_B_Valid_46_delay_2_5;
  reg                 io_B_Valid_46_delay_3_4;
  reg                 io_B_Valid_46_delay_4_3;
  reg                 io_B_Valid_46_delay_5_2;
  reg                 io_B_Valid_46_delay_6_1;
  reg                 io_B_Valid_46_delay_7;
  reg                 io_A_Valid_7_delay_1_46;
  reg                 io_A_Valid_7_delay_2_45;
  reg                 io_A_Valid_7_delay_3_44;
  reg                 io_A_Valid_7_delay_4_43;
  reg                 io_A_Valid_7_delay_5_42;
  reg                 io_A_Valid_7_delay_6_41;
  reg                 io_A_Valid_7_delay_7_40;
  reg                 io_A_Valid_7_delay_8_39;
  reg                 io_A_Valid_7_delay_9_38;
  reg                 io_A_Valid_7_delay_10_37;
  reg                 io_A_Valid_7_delay_11_36;
  reg                 io_A_Valid_7_delay_12_35;
  reg                 io_A_Valid_7_delay_13_34;
  reg                 io_A_Valid_7_delay_14_33;
  reg                 io_A_Valid_7_delay_15_32;
  reg                 io_A_Valid_7_delay_16_31;
  reg                 io_A_Valid_7_delay_17_30;
  reg                 io_A_Valid_7_delay_18_29;
  reg                 io_A_Valid_7_delay_19_28;
  reg                 io_A_Valid_7_delay_20_27;
  reg                 io_A_Valid_7_delay_21_26;
  reg                 io_A_Valid_7_delay_22_25;
  reg                 io_A_Valid_7_delay_23_24;
  reg                 io_A_Valid_7_delay_24_23;
  reg                 io_A_Valid_7_delay_25_22;
  reg                 io_A_Valid_7_delay_26_21;
  reg                 io_A_Valid_7_delay_27_20;
  reg                 io_A_Valid_7_delay_28_19;
  reg                 io_A_Valid_7_delay_29_18;
  reg                 io_A_Valid_7_delay_30_17;
  reg                 io_A_Valid_7_delay_31_16;
  reg                 io_A_Valid_7_delay_32_15;
  reg                 io_A_Valid_7_delay_33_14;
  reg                 io_A_Valid_7_delay_34_13;
  reg                 io_A_Valid_7_delay_35_12;
  reg                 io_A_Valid_7_delay_36_11;
  reg                 io_A_Valid_7_delay_37_10;
  reg                 io_A_Valid_7_delay_38_9;
  reg                 io_A_Valid_7_delay_39_8;
  reg                 io_A_Valid_7_delay_40_7;
  reg                 io_A_Valid_7_delay_41_6;
  reg                 io_A_Valid_7_delay_42_5;
  reg                 io_A_Valid_7_delay_43_4;
  reg                 io_A_Valid_7_delay_44_3;
  reg                 io_A_Valid_7_delay_45_2;
  reg                 io_A_Valid_7_delay_46_1;
  reg                 io_A_Valid_7_delay_47;
  reg                 io_B_Valid_47_delay_1_6;
  reg                 io_B_Valid_47_delay_2_5;
  reg                 io_B_Valid_47_delay_3_4;
  reg                 io_B_Valid_47_delay_4_3;
  reg                 io_B_Valid_47_delay_5_2;
  reg                 io_B_Valid_47_delay_6_1;
  reg                 io_B_Valid_47_delay_7;
  reg                 io_A_Valid_7_delay_1_47;
  reg                 io_A_Valid_7_delay_2_46;
  reg                 io_A_Valid_7_delay_3_45;
  reg                 io_A_Valid_7_delay_4_44;
  reg                 io_A_Valid_7_delay_5_43;
  reg                 io_A_Valid_7_delay_6_42;
  reg                 io_A_Valid_7_delay_7_41;
  reg                 io_A_Valid_7_delay_8_40;
  reg                 io_A_Valid_7_delay_9_39;
  reg                 io_A_Valid_7_delay_10_38;
  reg                 io_A_Valid_7_delay_11_37;
  reg                 io_A_Valid_7_delay_12_36;
  reg                 io_A_Valid_7_delay_13_35;
  reg                 io_A_Valid_7_delay_14_34;
  reg                 io_A_Valid_7_delay_15_33;
  reg                 io_A_Valid_7_delay_16_32;
  reg                 io_A_Valid_7_delay_17_31;
  reg                 io_A_Valid_7_delay_18_30;
  reg                 io_A_Valid_7_delay_19_29;
  reg                 io_A_Valid_7_delay_20_28;
  reg                 io_A_Valid_7_delay_21_27;
  reg                 io_A_Valid_7_delay_22_26;
  reg                 io_A_Valid_7_delay_23_25;
  reg                 io_A_Valid_7_delay_24_24;
  reg                 io_A_Valid_7_delay_25_23;
  reg                 io_A_Valid_7_delay_26_22;
  reg                 io_A_Valid_7_delay_27_21;
  reg                 io_A_Valid_7_delay_28_20;
  reg                 io_A_Valid_7_delay_29_19;
  reg                 io_A_Valid_7_delay_30_18;
  reg                 io_A_Valid_7_delay_31_17;
  reg                 io_A_Valid_7_delay_32_16;
  reg                 io_A_Valid_7_delay_33_15;
  reg                 io_A_Valid_7_delay_34_14;
  reg                 io_A_Valid_7_delay_35_13;
  reg                 io_A_Valid_7_delay_36_12;
  reg                 io_A_Valid_7_delay_37_11;
  reg                 io_A_Valid_7_delay_38_10;
  reg                 io_A_Valid_7_delay_39_9;
  reg                 io_A_Valid_7_delay_40_8;
  reg                 io_A_Valid_7_delay_41_7;
  reg                 io_A_Valid_7_delay_42_6;
  reg                 io_A_Valid_7_delay_43_5;
  reg                 io_A_Valid_7_delay_44_4;
  reg                 io_A_Valid_7_delay_45_3;
  reg                 io_A_Valid_7_delay_46_2;
  reg                 io_A_Valid_7_delay_47_1;
  reg                 io_A_Valid_7_delay_48;
  reg                 io_B_Valid_48_delay_1_6;
  reg                 io_B_Valid_48_delay_2_5;
  reg                 io_B_Valid_48_delay_3_4;
  reg                 io_B_Valid_48_delay_4_3;
  reg                 io_B_Valid_48_delay_5_2;
  reg                 io_B_Valid_48_delay_6_1;
  reg                 io_B_Valid_48_delay_7;
  reg                 io_A_Valid_7_delay_1_48;
  reg                 io_A_Valid_7_delay_2_47;
  reg                 io_A_Valid_7_delay_3_46;
  reg                 io_A_Valid_7_delay_4_45;
  reg                 io_A_Valid_7_delay_5_44;
  reg                 io_A_Valid_7_delay_6_43;
  reg                 io_A_Valid_7_delay_7_42;
  reg                 io_A_Valid_7_delay_8_41;
  reg                 io_A_Valid_7_delay_9_40;
  reg                 io_A_Valid_7_delay_10_39;
  reg                 io_A_Valid_7_delay_11_38;
  reg                 io_A_Valid_7_delay_12_37;
  reg                 io_A_Valid_7_delay_13_36;
  reg                 io_A_Valid_7_delay_14_35;
  reg                 io_A_Valid_7_delay_15_34;
  reg                 io_A_Valid_7_delay_16_33;
  reg                 io_A_Valid_7_delay_17_32;
  reg                 io_A_Valid_7_delay_18_31;
  reg                 io_A_Valid_7_delay_19_30;
  reg                 io_A_Valid_7_delay_20_29;
  reg                 io_A_Valid_7_delay_21_28;
  reg                 io_A_Valid_7_delay_22_27;
  reg                 io_A_Valid_7_delay_23_26;
  reg                 io_A_Valid_7_delay_24_25;
  reg                 io_A_Valid_7_delay_25_24;
  reg                 io_A_Valid_7_delay_26_23;
  reg                 io_A_Valid_7_delay_27_22;
  reg                 io_A_Valid_7_delay_28_21;
  reg                 io_A_Valid_7_delay_29_20;
  reg                 io_A_Valid_7_delay_30_19;
  reg                 io_A_Valid_7_delay_31_18;
  reg                 io_A_Valid_7_delay_32_17;
  reg                 io_A_Valid_7_delay_33_16;
  reg                 io_A_Valid_7_delay_34_15;
  reg                 io_A_Valid_7_delay_35_14;
  reg                 io_A_Valid_7_delay_36_13;
  reg                 io_A_Valid_7_delay_37_12;
  reg                 io_A_Valid_7_delay_38_11;
  reg                 io_A_Valid_7_delay_39_10;
  reg                 io_A_Valid_7_delay_40_9;
  reg                 io_A_Valid_7_delay_41_8;
  reg                 io_A_Valid_7_delay_42_7;
  reg                 io_A_Valid_7_delay_43_6;
  reg                 io_A_Valid_7_delay_44_5;
  reg                 io_A_Valid_7_delay_45_4;
  reg                 io_A_Valid_7_delay_46_3;
  reg                 io_A_Valid_7_delay_47_2;
  reg                 io_A_Valid_7_delay_48_1;
  reg                 io_A_Valid_7_delay_49;
  reg                 io_B_Valid_49_delay_1_6;
  reg                 io_B_Valid_49_delay_2_5;
  reg                 io_B_Valid_49_delay_3_4;
  reg                 io_B_Valid_49_delay_4_3;
  reg                 io_B_Valid_49_delay_5_2;
  reg                 io_B_Valid_49_delay_6_1;
  reg                 io_B_Valid_49_delay_7;
  reg                 io_A_Valid_7_delay_1_49;
  reg                 io_A_Valid_7_delay_2_48;
  reg                 io_A_Valid_7_delay_3_47;
  reg                 io_A_Valid_7_delay_4_46;
  reg                 io_A_Valid_7_delay_5_45;
  reg                 io_A_Valid_7_delay_6_44;
  reg                 io_A_Valid_7_delay_7_43;
  reg                 io_A_Valid_7_delay_8_42;
  reg                 io_A_Valid_7_delay_9_41;
  reg                 io_A_Valid_7_delay_10_40;
  reg                 io_A_Valid_7_delay_11_39;
  reg                 io_A_Valid_7_delay_12_38;
  reg                 io_A_Valid_7_delay_13_37;
  reg                 io_A_Valid_7_delay_14_36;
  reg                 io_A_Valid_7_delay_15_35;
  reg                 io_A_Valid_7_delay_16_34;
  reg                 io_A_Valid_7_delay_17_33;
  reg                 io_A_Valid_7_delay_18_32;
  reg                 io_A_Valid_7_delay_19_31;
  reg                 io_A_Valid_7_delay_20_30;
  reg                 io_A_Valid_7_delay_21_29;
  reg                 io_A_Valid_7_delay_22_28;
  reg                 io_A_Valid_7_delay_23_27;
  reg                 io_A_Valid_7_delay_24_26;
  reg                 io_A_Valid_7_delay_25_25;
  reg                 io_A_Valid_7_delay_26_24;
  reg                 io_A_Valid_7_delay_27_23;
  reg                 io_A_Valid_7_delay_28_22;
  reg                 io_A_Valid_7_delay_29_21;
  reg                 io_A_Valid_7_delay_30_20;
  reg                 io_A_Valid_7_delay_31_19;
  reg                 io_A_Valid_7_delay_32_18;
  reg                 io_A_Valid_7_delay_33_17;
  reg                 io_A_Valid_7_delay_34_16;
  reg                 io_A_Valid_7_delay_35_15;
  reg                 io_A_Valid_7_delay_36_14;
  reg                 io_A_Valid_7_delay_37_13;
  reg                 io_A_Valid_7_delay_38_12;
  reg                 io_A_Valid_7_delay_39_11;
  reg                 io_A_Valid_7_delay_40_10;
  reg                 io_A_Valid_7_delay_41_9;
  reg                 io_A_Valid_7_delay_42_8;
  reg                 io_A_Valid_7_delay_43_7;
  reg                 io_A_Valid_7_delay_44_6;
  reg                 io_A_Valid_7_delay_45_5;
  reg                 io_A_Valid_7_delay_46_4;
  reg                 io_A_Valid_7_delay_47_3;
  reg                 io_A_Valid_7_delay_48_2;
  reg                 io_A_Valid_7_delay_49_1;
  reg                 io_A_Valid_7_delay_50;
  reg                 io_B_Valid_50_delay_1_6;
  reg                 io_B_Valid_50_delay_2_5;
  reg                 io_B_Valid_50_delay_3_4;
  reg                 io_B_Valid_50_delay_4_3;
  reg                 io_B_Valid_50_delay_5_2;
  reg                 io_B_Valid_50_delay_6_1;
  reg                 io_B_Valid_50_delay_7;
  reg                 io_A_Valid_7_delay_1_50;
  reg                 io_A_Valid_7_delay_2_49;
  reg                 io_A_Valid_7_delay_3_48;
  reg                 io_A_Valid_7_delay_4_47;
  reg                 io_A_Valid_7_delay_5_46;
  reg                 io_A_Valid_7_delay_6_45;
  reg                 io_A_Valid_7_delay_7_44;
  reg                 io_A_Valid_7_delay_8_43;
  reg                 io_A_Valid_7_delay_9_42;
  reg                 io_A_Valid_7_delay_10_41;
  reg                 io_A_Valid_7_delay_11_40;
  reg                 io_A_Valid_7_delay_12_39;
  reg                 io_A_Valid_7_delay_13_38;
  reg                 io_A_Valid_7_delay_14_37;
  reg                 io_A_Valid_7_delay_15_36;
  reg                 io_A_Valid_7_delay_16_35;
  reg                 io_A_Valid_7_delay_17_34;
  reg                 io_A_Valid_7_delay_18_33;
  reg                 io_A_Valid_7_delay_19_32;
  reg                 io_A_Valid_7_delay_20_31;
  reg                 io_A_Valid_7_delay_21_30;
  reg                 io_A_Valid_7_delay_22_29;
  reg                 io_A_Valid_7_delay_23_28;
  reg                 io_A_Valid_7_delay_24_27;
  reg                 io_A_Valid_7_delay_25_26;
  reg                 io_A_Valid_7_delay_26_25;
  reg                 io_A_Valid_7_delay_27_24;
  reg                 io_A_Valid_7_delay_28_23;
  reg                 io_A_Valid_7_delay_29_22;
  reg                 io_A_Valid_7_delay_30_21;
  reg                 io_A_Valid_7_delay_31_20;
  reg                 io_A_Valid_7_delay_32_19;
  reg                 io_A_Valid_7_delay_33_18;
  reg                 io_A_Valid_7_delay_34_17;
  reg                 io_A_Valid_7_delay_35_16;
  reg                 io_A_Valid_7_delay_36_15;
  reg                 io_A_Valid_7_delay_37_14;
  reg                 io_A_Valid_7_delay_38_13;
  reg                 io_A_Valid_7_delay_39_12;
  reg                 io_A_Valid_7_delay_40_11;
  reg                 io_A_Valid_7_delay_41_10;
  reg                 io_A_Valid_7_delay_42_9;
  reg                 io_A_Valid_7_delay_43_8;
  reg                 io_A_Valid_7_delay_44_7;
  reg                 io_A_Valid_7_delay_45_6;
  reg                 io_A_Valid_7_delay_46_5;
  reg                 io_A_Valid_7_delay_47_4;
  reg                 io_A_Valid_7_delay_48_3;
  reg                 io_A_Valid_7_delay_49_2;
  reg                 io_A_Valid_7_delay_50_1;
  reg                 io_A_Valid_7_delay_51;
  reg                 io_B_Valid_51_delay_1_6;
  reg                 io_B_Valid_51_delay_2_5;
  reg                 io_B_Valid_51_delay_3_4;
  reg                 io_B_Valid_51_delay_4_3;
  reg                 io_B_Valid_51_delay_5_2;
  reg                 io_B_Valid_51_delay_6_1;
  reg                 io_B_Valid_51_delay_7;
  reg                 io_A_Valid_7_delay_1_51;
  reg                 io_A_Valid_7_delay_2_50;
  reg                 io_A_Valid_7_delay_3_49;
  reg                 io_A_Valid_7_delay_4_48;
  reg                 io_A_Valid_7_delay_5_47;
  reg                 io_A_Valid_7_delay_6_46;
  reg                 io_A_Valid_7_delay_7_45;
  reg                 io_A_Valid_7_delay_8_44;
  reg                 io_A_Valid_7_delay_9_43;
  reg                 io_A_Valid_7_delay_10_42;
  reg                 io_A_Valid_7_delay_11_41;
  reg                 io_A_Valid_7_delay_12_40;
  reg                 io_A_Valid_7_delay_13_39;
  reg                 io_A_Valid_7_delay_14_38;
  reg                 io_A_Valid_7_delay_15_37;
  reg                 io_A_Valid_7_delay_16_36;
  reg                 io_A_Valid_7_delay_17_35;
  reg                 io_A_Valid_7_delay_18_34;
  reg                 io_A_Valid_7_delay_19_33;
  reg                 io_A_Valid_7_delay_20_32;
  reg                 io_A_Valid_7_delay_21_31;
  reg                 io_A_Valid_7_delay_22_30;
  reg                 io_A_Valid_7_delay_23_29;
  reg                 io_A_Valid_7_delay_24_28;
  reg                 io_A_Valid_7_delay_25_27;
  reg                 io_A_Valid_7_delay_26_26;
  reg                 io_A_Valid_7_delay_27_25;
  reg                 io_A_Valid_7_delay_28_24;
  reg                 io_A_Valid_7_delay_29_23;
  reg                 io_A_Valid_7_delay_30_22;
  reg                 io_A_Valid_7_delay_31_21;
  reg                 io_A_Valid_7_delay_32_20;
  reg                 io_A_Valid_7_delay_33_19;
  reg                 io_A_Valid_7_delay_34_18;
  reg                 io_A_Valid_7_delay_35_17;
  reg                 io_A_Valid_7_delay_36_16;
  reg                 io_A_Valid_7_delay_37_15;
  reg                 io_A_Valid_7_delay_38_14;
  reg                 io_A_Valid_7_delay_39_13;
  reg                 io_A_Valid_7_delay_40_12;
  reg                 io_A_Valid_7_delay_41_11;
  reg                 io_A_Valid_7_delay_42_10;
  reg                 io_A_Valid_7_delay_43_9;
  reg                 io_A_Valid_7_delay_44_8;
  reg                 io_A_Valid_7_delay_45_7;
  reg                 io_A_Valid_7_delay_46_6;
  reg                 io_A_Valid_7_delay_47_5;
  reg                 io_A_Valid_7_delay_48_4;
  reg                 io_A_Valid_7_delay_49_3;
  reg                 io_A_Valid_7_delay_50_2;
  reg                 io_A_Valid_7_delay_51_1;
  reg                 io_A_Valid_7_delay_52;
  reg                 io_B_Valid_52_delay_1_6;
  reg                 io_B_Valid_52_delay_2_5;
  reg                 io_B_Valid_52_delay_3_4;
  reg                 io_B_Valid_52_delay_4_3;
  reg                 io_B_Valid_52_delay_5_2;
  reg                 io_B_Valid_52_delay_6_1;
  reg                 io_B_Valid_52_delay_7;
  reg                 io_A_Valid_7_delay_1_52;
  reg                 io_A_Valid_7_delay_2_51;
  reg                 io_A_Valid_7_delay_3_50;
  reg                 io_A_Valid_7_delay_4_49;
  reg                 io_A_Valid_7_delay_5_48;
  reg                 io_A_Valid_7_delay_6_47;
  reg                 io_A_Valid_7_delay_7_46;
  reg                 io_A_Valid_7_delay_8_45;
  reg                 io_A_Valid_7_delay_9_44;
  reg                 io_A_Valid_7_delay_10_43;
  reg                 io_A_Valid_7_delay_11_42;
  reg                 io_A_Valid_7_delay_12_41;
  reg                 io_A_Valid_7_delay_13_40;
  reg                 io_A_Valid_7_delay_14_39;
  reg                 io_A_Valid_7_delay_15_38;
  reg                 io_A_Valid_7_delay_16_37;
  reg                 io_A_Valid_7_delay_17_36;
  reg                 io_A_Valid_7_delay_18_35;
  reg                 io_A_Valid_7_delay_19_34;
  reg                 io_A_Valid_7_delay_20_33;
  reg                 io_A_Valid_7_delay_21_32;
  reg                 io_A_Valid_7_delay_22_31;
  reg                 io_A_Valid_7_delay_23_30;
  reg                 io_A_Valid_7_delay_24_29;
  reg                 io_A_Valid_7_delay_25_28;
  reg                 io_A_Valid_7_delay_26_27;
  reg                 io_A_Valid_7_delay_27_26;
  reg                 io_A_Valid_7_delay_28_25;
  reg                 io_A_Valid_7_delay_29_24;
  reg                 io_A_Valid_7_delay_30_23;
  reg                 io_A_Valid_7_delay_31_22;
  reg                 io_A_Valid_7_delay_32_21;
  reg                 io_A_Valid_7_delay_33_20;
  reg                 io_A_Valid_7_delay_34_19;
  reg                 io_A_Valid_7_delay_35_18;
  reg                 io_A_Valid_7_delay_36_17;
  reg                 io_A_Valid_7_delay_37_16;
  reg                 io_A_Valid_7_delay_38_15;
  reg                 io_A_Valid_7_delay_39_14;
  reg                 io_A_Valid_7_delay_40_13;
  reg                 io_A_Valid_7_delay_41_12;
  reg                 io_A_Valid_7_delay_42_11;
  reg                 io_A_Valid_7_delay_43_10;
  reg                 io_A_Valid_7_delay_44_9;
  reg                 io_A_Valid_7_delay_45_8;
  reg                 io_A_Valid_7_delay_46_7;
  reg                 io_A_Valid_7_delay_47_6;
  reg                 io_A_Valid_7_delay_48_5;
  reg                 io_A_Valid_7_delay_49_4;
  reg                 io_A_Valid_7_delay_50_3;
  reg                 io_A_Valid_7_delay_51_2;
  reg                 io_A_Valid_7_delay_52_1;
  reg                 io_A_Valid_7_delay_53;
  reg                 io_B_Valid_53_delay_1_6;
  reg                 io_B_Valid_53_delay_2_5;
  reg                 io_B_Valid_53_delay_3_4;
  reg                 io_B_Valid_53_delay_4_3;
  reg                 io_B_Valid_53_delay_5_2;
  reg                 io_B_Valid_53_delay_6_1;
  reg                 io_B_Valid_53_delay_7;
  reg                 io_A_Valid_7_delay_1_53;
  reg                 io_A_Valid_7_delay_2_52;
  reg                 io_A_Valid_7_delay_3_51;
  reg                 io_A_Valid_7_delay_4_50;
  reg                 io_A_Valid_7_delay_5_49;
  reg                 io_A_Valid_7_delay_6_48;
  reg                 io_A_Valid_7_delay_7_47;
  reg                 io_A_Valid_7_delay_8_46;
  reg                 io_A_Valid_7_delay_9_45;
  reg                 io_A_Valid_7_delay_10_44;
  reg                 io_A_Valid_7_delay_11_43;
  reg                 io_A_Valid_7_delay_12_42;
  reg                 io_A_Valid_7_delay_13_41;
  reg                 io_A_Valid_7_delay_14_40;
  reg                 io_A_Valid_7_delay_15_39;
  reg                 io_A_Valid_7_delay_16_38;
  reg                 io_A_Valid_7_delay_17_37;
  reg                 io_A_Valid_7_delay_18_36;
  reg                 io_A_Valid_7_delay_19_35;
  reg                 io_A_Valid_7_delay_20_34;
  reg                 io_A_Valid_7_delay_21_33;
  reg                 io_A_Valid_7_delay_22_32;
  reg                 io_A_Valid_7_delay_23_31;
  reg                 io_A_Valid_7_delay_24_30;
  reg                 io_A_Valid_7_delay_25_29;
  reg                 io_A_Valid_7_delay_26_28;
  reg                 io_A_Valid_7_delay_27_27;
  reg                 io_A_Valid_7_delay_28_26;
  reg                 io_A_Valid_7_delay_29_25;
  reg                 io_A_Valid_7_delay_30_24;
  reg                 io_A_Valid_7_delay_31_23;
  reg                 io_A_Valid_7_delay_32_22;
  reg                 io_A_Valid_7_delay_33_21;
  reg                 io_A_Valid_7_delay_34_20;
  reg                 io_A_Valid_7_delay_35_19;
  reg                 io_A_Valid_7_delay_36_18;
  reg                 io_A_Valid_7_delay_37_17;
  reg                 io_A_Valid_7_delay_38_16;
  reg                 io_A_Valid_7_delay_39_15;
  reg                 io_A_Valid_7_delay_40_14;
  reg                 io_A_Valid_7_delay_41_13;
  reg                 io_A_Valid_7_delay_42_12;
  reg                 io_A_Valid_7_delay_43_11;
  reg                 io_A_Valid_7_delay_44_10;
  reg                 io_A_Valid_7_delay_45_9;
  reg                 io_A_Valid_7_delay_46_8;
  reg                 io_A_Valid_7_delay_47_7;
  reg                 io_A_Valid_7_delay_48_6;
  reg                 io_A_Valid_7_delay_49_5;
  reg                 io_A_Valid_7_delay_50_4;
  reg                 io_A_Valid_7_delay_51_3;
  reg                 io_A_Valid_7_delay_52_2;
  reg                 io_A_Valid_7_delay_53_1;
  reg                 io_A_Valid_7_delay_54;
  reg                 io_B_Valid_54_delay_1_6;
  reg                 io_B_Valid_54_delay_2_5;
  reg                 io_B_Valid_54_delay_3_4;
  reg                 io_B_Valid_54_delay_4_3;
  reg                 io_B_Valid_54_delay_5_2;
  reg                 io_B_Valid_54_delay_6_1;
  reg                 io_B_Valid_54_delay_7;
  reg                 io_A_Valid_7_delay_1_54;
  reg                 io_A_Valid_7_delay_2_53;
  reg                 io_A_Valid_7_delay_3_52;
  reg                 io_A_Valid_7_delay_4_51;
  reg                 io_A_Valid_7_delay_5_50;
  reg                 io_A_Valid_7_delay_6_49;
  reg                 io_A_Valid_7_delay_7_48;
  reg                 io_A_Valid_7_delay_8_47;
  reg                 io_A_Valid_7_delay_9_46;
  reg                 io_A_Valid_7_delay_10_45;
  reg                 io_A_Valid_7_delay_11_44;
  reg                 io_A_Valid_7_delay_12_43;
  reg                 io_A_Valid_7_delay_13_42;
  reg                 io_A_Valid_7_delay_14_41;
  reg                 io_A_Valid_7_delay_15_40;
  reg                 io_A_Valid_7_delay_16_39;
  reg                 io_A_Valid_7_delay_17_38;
  reg                 io_A_Valid_7_delay_18_37;
  reg                 io_A_Valid_7_delay_19_36;
  reg                 io_A_Valid_7_delay_20_35;
  reg                 io_A_Valid_7_delay_21_34;
  reg                 io_A_Valid_7_delay_22_33;
  reg                 io_A_Valid_7_delay_23_32;
  reg                 io_A_Valid_7_delay_24_31;
  reg                 io_A_Valid_7_delay_25_30;
  reg                 io_A_Valid_7_delay_26_29;
  reg                 io_A_Valid_7_delay_27_28;
  reg                 io_A_Valid_7_delay_28_27;
  reg                 io_A_Valid_7_delay_29_26;
  reg                 io_A_Valid_7_delay_30_25;
  reg                 io_A_Valid_7_delay_31_24;
  reg                 io_A_Valid_7_delay_32_23;
  reg                 io_A_Valid_7_delay_33_22;
  reg                 io_A_Valid_7_delay_34_21;
  reg                 io_A_Valid_7_delay_35_20;
  reg                 io_A_Valid_7_delay_36_19;
  reg                 io_A_Valid_7_delay_37_18;
  reg                 io_A_Valid_7_delay_38_17;
  reg                 io_A_Valid_7_delay_39_16;
  reg                 io_A_Valid_7_delay_40_15;
  reg                 io_A_Valid_7_delay_41_14;
  reg                 io_A_Valid_7_delay_42_13;
  reg                 io_A_Valid_7_delay_43_12;
  reg                 io_A_Valid_7_delay_44_11;
  reg                 io_A_Valid_7_delay_45_10;
  reg                 io_A_Valid_7_delay_46_9;
  reg                 io_A_Valid_7_delay_47_8;
  reg                 io_A_Valid_7_delay_48_7;
  reg                 io_A_Valid_7_delay_49_6;
  reg                 io_A_Valid_7_delay_50_5;
  reg                 io_A_Valid_7_delay_51_4;
  reg                 io_A_Valid_7_delay_52_3;
  reg                 io_A_Valid_7_delay_53_2;
  reg                 io_A_Valid_7_delay_54_1;
  reg                 io_A_Valid_7_delay_55;
  reg                 io_B_Valid_55_delay_1_6;
  reg                 io_B_Valid_55_delay_2_5;
  reg                 io_B_Valid_55_delay_3_4;
  reg                 io_B_Valid_55_delay_4_3;
  reg                 io_B_Valid_55_delay_5_2;
  reg                 io_B_Valid_55_delay_6_1;
  reg                 io_B_Valid_55_delay_7;
  reg                 io_A_Valid_7_delay_1_55;
  reg                 io_A_Valid_7_delay_2_54;
  reg                 io_A_Valid_7_delay_3_53;
  reg                 io_A_Valid_7_delay_4_52;
  reg                 io_A_Valid_7_delay_5_51;
  reg                 io_A_Valid_7_delay_6_50;
  reg                 io_A_Valid_7_delay_7_49;
  reg                 io_A_Valid_7_delay_8_48;
  reg                 io_A_Valid_7_delay_9_47;
  reg                 io_A_Valid_7_delay_10_46;
  reg                 io_A_Valid_7_delay_11_45;
  reg                 io_A_Valid_7_delay_12_44;
  reg                 io_A_Valid_7_delay_13_43;
  reg                 io_A_Valid_7_delay_14_42;
  reg                 io_A_Valid_7_delay_15_41;
  reg                 io_A_Valid_7_delay_16_40;
  reg                 io_A_Valid_7_delay_17_39;
  reg                 io_A_Valid_7_delay_18_38;
  reg                 io_A_Valid_7_delay_19_37;
  reg                 io_A_Valid_7_delay_20_36;
  reg                 io_A_Valid_7_delay_21_35;
  reg                 io_A_Valid_7_delay_22_34;
  reg                 io_A_Valid_7_delay_23_33;
  reg                 io_A_Valid_7_delay_24_32;
  reg                 io_A_Valid_7_delay_25_31;
  reg                 io_A_Valid_7_delay_26_30;
  reg                 io_A_Valid_7_delay_27_29;
  reg                 io_A_Valid_7_delay_28_28;
  reg                 io_A_Valid_7_delay_29_27;
  reg                 io_A_Valid_7_delay_30_26;
  reg                 io_A_Valid_7_delay_31_25;
  reg                 io_A_Valid_7_delay_32_24;
  reg                 io_A_Valid_7_delay_33_23;
  reg                 io_A_Valid_7_delay_34_22;
  reg                 io_A_Valid_7_delay_35_21;
  reg                 io_A_Valid_7_delay_36_20;
  reg                 io_A_Valid_7_delay_37_19;
  reg                 io_A_Valid_7_delay_38_18;
  reg                 io_A_Valid_7_delay_39_17;
  reg                 io_A_Valid_7_delay_40_16;
  reg                 io_A_Valid_7_delay_41_15;
  reg                 io_A_Valid_7_delay_42_14;
  reg                 io_A_Valid_7_delay_43_13;
  reg                 io_A_Valid_7_delay_44_12;
  reg                 io_A_Valid_7_delay_45_11;
  reg                 io_A_Valid_7_delay_46_10;
  reg                 io_A_Valid_7_delay_47_9;
  reg                 io_A_Valid_7_delay_48_8;
  reg                 io_A_Valid_7_delay_49_7;
  reg                 io_A_Valid_7_delay_50_6;
  reg                 io_A_Valid_7_delay_51_5;
  reg                 io_A_Valid_7_delay_52_4;
  reg                 io_A_Valid_7_delay_53_3;
  reg                 io_A_Valid_7_delay_54_2;
  reg                 io_A_Valid_7_delay_55_1;
  reg                 io_A_Valid_7_delay_56;
  reg                 io_B_Valid_56_delay_1_6;
  reg                 io_B_Valid_56_delay_2_5;
  reg                 io_B_Valid_56_delay_3_4;
  reg                 io_B_Valid_56_delay_4_3;
  reg                 io_B_Valid_56_delay_5_2;
  reg                 io_B_Valid_56_delay_6_1;
  reg                 io_B_Valid_56_delay_7;
  reg                 io_A_Valid_7_delay_1_56;
  reg                 io_A_Valid_7_delay_2_55;
  reg                 io_A_Valid_7_delay_3_54;
  reg                 io_A_Valid_7_delay_4_53;
  reg                 io_A_Valid_7_delay_5_52;
  reg                 io_A_Valid_7_delay_6_51;
  reg                 io_A_Valid_7_delay_7_50;
  reg                 io_A_Valid_7_delay_8_49;
  reg                 io_A_Valid_7_delay_9_48;
  reg                 io_A_Valid_7_delay_10_47;
  reg                 io_A_Valid_7_delay_11_46;
  reg                 io_A_Valid_7_delay_12_45;
  reg                 io_A_Valid_7_delay_13_44;
  reg                 io_A_Valid_7_delay_14_43;
  reg                 io_A_Valid_7_delay_15_42;
  reg                 io_A_Valid_7_delay_16_41;
  reg                 io_A_Valid_7_delay_17_40;
  reg                 io_A_Valid_7_delay_18_39;
  reg                 io_A_Valid_7_delay_19_38;
  reg                 io_A_Valid_7_delay_20_37;
  reg                 io_A_Valid_7_delay_21_36;
  reg                 io_A_Valid_7_delay_22_35;
  reg                 io_A_Valid_7_delay_23_34;
  reg                 io_A_Valid_7_delay_24_33;
  reg                 io_A_Valid_7_delay_25_32;
  reg                 io_A_Valid_7_delay_26_31;
  reg                 io_A_Valid_7_delay_27_30;
  reg                 io_A_Valid_7_delay_28_29;
  reg                 io_A_Valid_7_delay_29_28;
  reg                 io_A_Valid_7_delay_30_27;
  reg                 io_A_Valid_7_delay_31_26;
  reg                 io_A_Valid_7_delay_32_25;
  reg                 io_A_Valid_7_delay_33_24;
  reg                 io_A_Valid_7_delay_34_23;
  reg                 io_A_Valid_7_delay_35_22;
  reg                 io_A_Valid_7_delay_36_21;
  reg                 io_A_Valid_7_delay_37_20;
  reg                 io_A_Valid_7_delay_38_19;
  reg                 io_A_Valid_7_delay_39_18;
  reg                 io_A_Valid_7_delay_40_17;
  reg                 io_A_Valid_7_delay_41_16;
  reg                 io_A_Valid_7_delay_42_15;
  reg                 io_A_Valid_7_delay_43_14;
  reg                 io_A_Valid_7_delay_44_13;
  reg                 io_A_Valid_7_delay_45_12;
  reg                 io_A_Valid_7_delay_46_11;
  reg                 io_A_Valid_7_delay_47_10;
  reg                 io_A_Valid_7_delay_48_9;
  reg                 io_A_Valid_7_delay_49_8;
  reg                 io_A_Valid_7_delay_50_7;
  reg                 io_A_Valid_7_delay_51_6;
  reg                 io_A_Valid_7_delay_52_5;
  reg                 io_A_Valid_7_delay_53_4;
  reg                 io_A_Valid_7_delay_54_3;
  reg                 io_A_Valid_7_delay_55_2;
  reg                 io_A_Valid_7_delay_56_1;
  reg                 io_A_Valid_7_delay_57;
  reg                 io_B_Valid_57_delay_1_6;
  reg                 io_B_Valid_57_delay_2_5;
  reg                 io_B_Valid_57_delay_3_4;
  reg                 io_B_Valid_57_delay_4_3;
  reg                 io_B_Valid_57_delay_5_2;
  reg                 io_B_Valid_57_delay_6_1;
  reg                 io_B_Valid_57_delay_7;
  reg                 io_A_Valid_7_delay_1_57;
  reg                 io_A_Valid_7_delay_2_56;
  reg                 io_A_Valid_7_delay_3_55;
  reg                 io_A_Valid_7_delay_4_54;
  reg                 io_A_Valid_7_delay_5_53;
  reg                 io_A_Valid_7_delay_6_52;
  reg                 io_A_Valid_7_delay_7_51;
  reg                 io_A_Valid_7_delay_8_50;
  reg                 io_A_Valid_7_delay_9_49;
  reg                 io_A_Valid_7_delay_10_48;
  reg                 io_A_Valid_7_delay_11_47;
  reg                 io_A_Valid_7_delay_12_46;
  reg                 io_A_Valid_7_delay_13_45;
  reg                 io_A_Valid_7_delay_14_44;
  reg                 io_A_Valid_7_delay_15_43;
  reg                 io_A_Valid_7_delay_16_42;
  reg                 io_A_Valid_7_delay_17_41;
  reg                 io_A_Valid_7_delay_18_40;
  reg                 io_A_Valid_7_delay_19_39;
  reg                 io_A_Valid_7_delay_20_38;
  reg                 io_A_Valid_7_delay_21_37;
  reg                 io_A_Valid_7_delay_22_36;
  reg                 io_A_Valid_7_delay_23_35;
  reg                 io_A_Valid_7_delay_24_34;
  reg                 io_A_Valid_7_delay_25_33;
  reg                 io_A_Valid_7_delay_26_32;
  reg                 io_A_Valid_7_delay_27_31;
  reg                 io_A_Valid_7_delay_28_30;
  reg                 io_A_Valid_7_delay_29_29;
  reg                 io_A_Valid_7_delay_30_28;
  reg                 io_A_Valid_7_delay_31_27;
  reg                 io_A_Valid_7_delay_32_26;
  reg                 io_A_Valid_7_delay_33_25;
  reg                 io_A_Valid_7_delay_34_24;
  reg                 io_A_Valid_7_delay_35_23;
  reg                 io_A_Valid_7_delay_36_22;
  reg                 io_A_Valid_7_delay_37_21;
  reg                 io_A_Valid_7_delay_38_20;
  reg                 io_A_Valid_7_delay_39_19;
  reg                 io_A_Valid_7_delay_40_18;
  reg                 io_A_Valid_7_delay_41_17;
  reg                 io_A_Valid_7_delay_42_16;
  reg                 io_A_Valid_7_delay_43_15;
  reg                 io_A_Valid_7_delay_44_14;
  reg                 io_A_Valid_7_delay_45_13;
  reg                 io_A_Valid_7_delay_46_12;
  reg                 io_A_Valid_7_delay_47_11;
  reg                 io_A_Valid_7_delay_48_10;
  reg                 io_A_Valid_7_delay_49_9;
  reg                 io_A_Valid_7_delay_50_8;
  reg                 io_A_Valid_7_delay_51_7;
  reg                 io_A_Valid_7_delay_52_6;
  reg                 io_A_Valid_7_delay_53_5;
  reg                 io_A_Valid_7_delay_54_4;
  reg                 io_A_Valid_7_delay_55_3;
  reg                 io_A_Valid_7_delay_56_2;
  reg                 io_A_Valid_7_delay_57_1;
  reg                 io_A_Valid_7_delay_58;
  reg                 io_B_Valid_58_delay_1_6;
  reg                 io_B_Valid_58_delay_2_5;
  reg                 io_B_Valid_58_delay_3_4;
  reg                 io_B_Valid_58_delay_4_3;
  reg                 io_B_Valid_58_delay_5_2;
  reg                 io_B_Valid_58_delay_6_1;
  reg                 io_B_Valid_58_delay_7;
  reg                 io_A_Valid_7_delay_1_58;
  reg                 io_A_Valid_7_delay_2_57;
  reg                 io_A_Valid_7_delay_3_56;
  reg                 io_A_Valid_7_delay_4_55;
  reg                 io_A_Valid_7_delay_5_54;
  reg                 io_A_Valid_7_delay_6_53;
  reg                 io_A_Valid_7_delay_7_52;
  reg                 io_A_Valid_7_delay_8_51;
  reg                 io_A_Valid_7_delay_9_50;
  reg                 io_A_Valid_7_delay_10_49;
  reg                 io_A_Valid_7_delay_11_48;
  reg                 io_A_Valid_7_delay_12_47;
  reg                 io_A_Valid_7_delay_13_46;
  reg                 io_A_Valid_7_delay_14_45;
  reg                 io_A_Valid_7_delay_15_44;
  reg                 io_A_Valid_7_delay_16_43;
  reg                 io_A_Valid_7_delay_17_42;
  reg                 io_A_Valid_7_delay_18_41;
  reg                 io_A_Valid_7_delay_19_40;
  reg                 io_A_Valid_7_delay_20_39;
  reg                 io_A_Valid_7_delay_21_38;
  reg                 io_A_Valid_7_delay_22_37;
  reg                 io_A_Valid_7_delay_23_36;
  reg                 io_A_Valid_7_delay_24_35;
  reg                 io_A_Valid_7_delay_25_34;
  reg                 io_A_Valid_7_delay_26_33;
  reg                 io_A_Valid_7_delay_27_32;
  reg                 io_A_Valid_7_delay_28_31;
  reg                 io_A_Valid_7_delay_29_30;
  reg                 io_A_Valid_7_delay_30_29;
  reg                 io_A_Valid_7_delay_31_28;
  reg                 io_A_Valid_7_delay_32_27;
  reg                 io_A_Valid_7_delay_33_26;
  reg                 io_A_Valid_7_delay_34_25;
  reg                 io_A_Valid_7_delay_35_24;
  reg                 io_A_Valid_7_delay_36_23;
  reg                 io_A_Valid_7_delay_37_22;
  reg                 io_A_Valid_7_delay_38_21;
  reg                 io_A_Valid_7_delay_39_20;
  reg                 io_A_Valid_7_delay_40_19;
  reg                 io_A_Valid_7_delay_41_18;
  reg                 io_A_Valid_7_delay_42_17;
  reg                 io_A_Valid_7_delay_43_16;
  reg                 io_A_Valid_7_delay_44_15;
  reg                 io_A_Valid_7_delay_45_14;
  reg                 io_A_Valid_7_delay_46_13;
  reg                 io_A_Valid_7_delay_47_12;
  reg                 io_A_Valid_7_delay_48_11;
  reg                 io_A_Valid_7_delay_49_10;
  reg                 io_A_Valid_7_delay_50_9;
  reg                 io_A_Valid_7_delay_51_8;
  reg                 io_A_Valid_7_delay_52_7;
  reg                 io_A_Valid_7_delay_53_6;
  reg                 io_A_Valid_7_delay_54_5;
  reg                 io_A_Valid_7_delay_55_4;
  reg                 io_A_Valid_7_delay_56_3;
  reg                 io_A_Valid_7_delay_57_2;
  reg                 io_A_Valid_7_delay_58_1;
  reg                 io_A_Valid_7_delay_59;
  reg                 io_B_Valid_59_delay_1_6;
  reg                 io_B_Valid_59_delay_2_5;
  reg                 io_B_Valid_59_delay_3_4;
  reg                 io_B_Valid_59_delay_4_3;
  reg                 io_B_Valid_59_delay_5_2;
  reg                 io_B_Valid_59_delay_6_1;
  reg                 io_B_Valid_59_delay_7;
  reg                 io_A_Valid_7_delay_1_59;
  reg                 io_A_Valid_7_delay_2_58;
  reg                 io_A_Valid_7_delay_3_57;
  reg                 io_A_Valid_7_delay_4_56;
  reg                 io_A_Valid_7_delay_5_55;
  reg                 io_A_Valid_7_delay_6_54;
  reg                 io_A_Valid_7_delay_7_53;
  reg                 io_A_Valid_7_delay_8_52;
  reg                 io_A_Valid_7_delay_9_51;
  reg                 io_A_Valid_7_delay_10_50;
  reg                 io_A_Valid_7_delay_11_49;
  reg                 io_A_Valid_7_delay_12_48;
  reg                 io_A_Valid_7_delay_13_47;
  reg                 io_A_Valid_7_delay_14_46;
  reg                 io_A_Valid_7_delay_15_45;
  reg                 io_A_Valid_7_delay_16_44;
  reg                 io_A_Valid_7_delay_17_43;
  reg                 io_A_Valid_7_delay_18_42;
  reg                 io_A_Valid_7_delay_19_41;
  reg                 io_A_Valid_7_delay_20_40;
  reg                 io_A_Valid_7_delay_21_39;
  reg                 io_A_Valid_7_delay_22_38;
  reg                 io_A_Valid_7_delay_23_37;
  reg                 io_A_Valid_7_delay_24_36;
  reg                 io_A_Valid_7_delay_25_35;
  reg                 io_A_Valid_7_delay_26_34;
  reg                 io_A_Valid_7_delay_27_33;
  reg                 io_A_Valid_7_delay_28_32;
  reg                 io_A_Valid_7_delay_29_31;
  reg                 io_A_Valid_7_delay_30_30;
  reg                 io_A_Valid_7_delay_31_29;
  reg                 io_A_Valid_7_delay_32_28;
  reg                 io_A_Valid_7_delay_33_27;
  reg                 io_A_Valid_7_delay_34_26;
  reg                 io_A_Valid_7_delay_35_25;
  reg                 io_A_Valid_7_delay_36_24;
  reg                 io_A_Valid_7_delay_37_23;
  reg                 io_A_Valid_7_delay_38_22;
  reg                 io_A_Valid_7_delay_39_21;
  reg                 io_A_Valid_7_delay_40_20;
  reg                 io_A_Valid_7_delay_41_19;
  reg                 io_A_Valid_7_delay_42_18;
  reg                 io_A_Valid_7_delay_43_17;
  reg                 io_A_Valid_7_delay_44_16;
  reg                 io_A_Valid_7_delay_45_15;
  reg                 io_A_Valid_7_delay_46_14;
  reg                 io_A_Valid_7_delay_47_13;
  reg                 io_A_Valid_7_delay_48_12;
  reg                 io_A_Valid_7_delay_49_11;
  reg                 io_A_Valid_7_delay_50_10;
  reg                 io_A_Valid_7_delay_51_9;
  reg                 io_A_Valid_7_delay_52_8;
  reg                 io_A_Valid_7_delay_53_7;
  reg                 io_A_Valid_7_delay_54_6;
  reg                 io_A_Valid_7_delay_55_5;
  reg                 io_A_Valid_7_delay_56_4;
  reg                 io_A_Valid_7_delay_57_3;
  reg                 io_A_Valid_7_delay_58_2;
  reg                 io_A_Valid_7_delay_59_1;
  reg                 io_A_Valid_7_delay_60;
  reg                 io_B_Valid_60_delay_1_6;
  reg                 io_B_Valid_60_delay_2_5;
  reg                 io_B_Valid_60_delay_3_4;
  reg                 io_B_Valid_60_delay_4_3;
  reg                 io_B_Valid_60_delay_5_2;
  reg                 io_B_Valid_60_delay_6_1;
  reg                 io_B_Valid_60_delay_7;
  reg                 io_A_Valid_7_delay_1_60;
  reg                 io_A_Valid_7_delay_2_59;
  reg                 io_A_Valid_7_delay_3_58;
  reg                 io_A_Valid_7_delay_4_57;
  reg                 io_A_Valid_7_delay_5_56;
  reg                 io_A_Valid_7_delay_6_55;
  reg                 io_A_Valid_7_delay_7_54;
  reg                 io_A_Valid_7_delay_8_53;
  reg                 io_A_Valid_7_delay_9_52;
  reg                 io_A_Valid_7_delay_10_51;
  reg                 io_A_Valid_7_delay_11_50;
  reg                 io_A_Valid_7_delay_12_49;
  reg                 io_A_Valid_7_delay_13_48;
  reg                 io_A_Valid_7_delay_14_47;
  reg                 io_A_Valid_7_delay_15_46;
  reg                 io_A_Valid_7_delay_16_45;
  reg                 io_A_Valid_7_delay_17_44;
  reg                 io_A_Valid_7_delay_18_43;
  reg                 io_A_Valid_7_delay_19_42;
  reg                 io_A_Valid_7_delay_20_41;
  reg                 io_A_Valid_7_delay_21_40;
  reg                 io_A_Valid_7_delay_22_39;
  reg                 io_A_Valid_7_delay_23_38;
  reg                 io_A_Valid_7_delay_24_37;
  reg                 io_A_Valid_7_delay_25_36;
  reg                 io_A_Valid_7_delay_26_35;
  reg                 io_A_Valid_7_delay_27_34;
  reg                 io_A_Valid_7_delay_28_33;
  reg                 io_A_Valid_7_delay_29_32;
  reg                 io_A_Valid_7_delay_30_31;
  reg                 io_A_Valid_7_delay_31_30;
  reg                 io_A_Valid_7_delay_32_29;
  reg                 io_A_Valid_7_delay_33_28;
  reg                 io_A_Valid_7_delay_34_27;
  reg                 io_A_Valid_7_delay_35_26;
  reg                 io_A_Valid_7_delay_36_25;
  reg                 io_A_Valid_7_delay_37_24;
  reg                 io_A_Valid_7_delay_38_23;
  reg                 io_A_Valid_7_delay_39_22;
  reg                 io_A_Valid_7_delay_40_21;
  reg                 io_A_Valid_7_delay_41_20;
  reg                 io_A_Valid_7_delay_42_19;
  reg                 io_A_Valid_7_delay_43_18;
  reg                 io_A_Valid_7_delay_44_17;
  reg                 io_A_Valid_7_delay_45_16;
  reg                 io_A_Valid_7_delay_46_15;
  reg                 io_A_Valid_7_delay_47_14;
  reg                 io_A_Valid_7_delay_48_13;
  reg                 io_A_Valid_7_delay_49_12;
  reg                 io_A_Valid_7_delay_50_11;
  reg                 io_A_Valid_7_delay_51_10;
  reg                 io_A_Valid_7_delay_52_9;
  reg                 io_A_Valid_7_delay_53_8;
  reg                 io_A_Valid_7_delay_54_7;
  reg                 io_A_Valid_7_delay_55_6;
  reg                 io_A_Valid_7_delay_56_5;
  reg                 io_A_Valid_7_delay_57_4;
  reg                 io_A_Valid_7_delay_58_3;
  reg                 io_A_Valid_7_delay_59_2;
  reg                 io_A_Valid_7_delay_60_1;
  reg                 io_A_Valid_7_delay_61;
  reg                 io_B_Valid_61_delay_1_6;
  reg                 io_B_Valid_61_delay_2_5;
  reg                 io_B_Valid_61_delay_3_4;
  reg                 io_B_Valid_61_delay_4_3;
  reg                 io_B_Valid_61_delay_5_2;
  reg                 io_B_Valid_61_delay_6_1;
  reg                 io_B_Valid_61_delay_7;
  reg                 io_A_Valid_7_delay_1_61;
  reg                 io_A_Valid_7_delay_2_60;
  reg                 io_A_Valid_7_delay_3_59;
  reg                 io_A_Valid_7_delay_4_58;
  reg                 io_A_Valid_7_delay_5_57;
  reg                 io_A_Valid_7_delay_6_56;
  reg                 io_A_Valid_7_delay_7_55;
  reg                 io_A_Valid_7_delay_8_54;
  reg                 io_A_Valid_7_delay_9_53;
  reg                 io_A_Valid_7_delay_10_52;
  reg                 io_A_Valid_7_delay_11_51;
  reg                 io_A_Valid_7_delay_12_50;
  reg                 io_A_Valid_7_delay_13_49;
  reg                 io_A_Valid_7_delay_14_48;
  reg                 io_A_Valid_7_delay_15_47;
  reg                 io_A_Valid_7_delay_16_46;
  reg                 io_A_Valid_7_delay_17_45;
  reg                 io_A_Valid_7_delay_18_44;
  reg                 io_A_Valid_7_delay_19_43;
  reg                 io_A_Valid_7_delay_20_42;
  reg                 io_A_Valid_7_delay_21_41;
  reg                 io_A_Valid_7_delay_22_40;
  reg                 io_A_Valid_7_delay_23_39;
  reg                 io_A_Valid_7_delay_24_38;
  reg                 io_A_Valid_7_delay_25_37;
  reg                 io_A_Valid_7_delay_26_36;
  reg                 io_A_Valid_7_delay_27_35;
  reg                 io_A_Valid_7_delay_28_34;
  reg                 io_A_Valid_7_delay_29_33;
  reg                 io_A_Valid_7_delay_30_32;
  reg                 io_A_Valid_7_delay_31_31;
  reg                 io_A_Valid_7_delay_32_30;
  reg                 io_A_Valid_7_delay_33_29;
  reg                 io_A_Valid_7_delay_34_28;
  reg                 io_A_Valid_7_delay_35_27;
  reg                 io_A_Valid_7_delay_36_26;
  reg                 io_A_Valid_7_delay_37_25;
  reg                 io_A_Valid_7_delay_38_24;
  reg                 io_A_Valid_7_delay_39_23;
  reg                 io_A_Valid_7_delay_40_22;
  reg                 io_A_Valid_7_delay_41_21;
  reg                 io_A_Valid_7_delay_42_20;
  reg                 io_A_Valid_7_delay_43_19;
  reg                 io_A_Valid_7_delay_44_18;
  reg                 io_A_Valid_7_delay_45_17;
  reg                 io_A_Valid_7_delay_46_16;
  reg                 io_A_Valid_7_delay_47_15;
  reg                 io_A_Valid_7_delay_48_14;
  reg                 io_A_Valid_7_delay_49_13;
  reg                 io_A_Valid_7_delay_50_12;
  reg                 io_A_Valid_7_delay_51_11;
  reg                 io_A_Valid_7_delay_52_10;
  reg                 io_A_Valid_7_delay_53_9;
  reg                 io_A_Valid_7_delay_54_8;
  reg                 io_A_Valid_7_delay_55_7;
  reg                 io_A_Valid_7_delay_56_6;
  reg                 io_A_Valid_7_delay_57_5;
  reg                 io_A_Valid_7_delay_58_4;
  reg                 io_A_Valid_7_delay_59_3;
  reg                 io_A_Valid_7_delay_60_2;
  reg                 io_A_Valid_7_delay_61_1;
  reg                 io_A_Valid_7_delay_62;
  reg                 io_B_Valid_62_delay_1_6;
  reg                 io_B_Valid_62_delay_2_5;
  reg                 io_B_Valid_62_delay_3_4;
  reg                 io_B_Valid_62_delay_4_3;
  reg                 io_B_Valid_62_delay_5_2;
  reg                 io_B_Valid_62_delay_6_1;
  reg                 io_B_Valid_62_delay_7;
  reg                 io_A_Valid_7_delay_1_62;
  reg                 io_A_Valid_7_delay_2_61;
  reg                 io_A_Valid_7_delay_3_60;
  reg                 io_A_Valid_7_delay_4_59;
  reg                 io_A_Valid_7_delay_5_58;
  reg                 io_A_Valid_7_delay_6_57;
  reg                 io_A_Valid_7_delay_7_56;
  reg                 io_A_Valid_7_delay_8_55;
  reg                 io_A_Valid_7_delay_9_54;
  reg                 io_A_Valid_7_delay_10_53;
  reg                 io_A_Valid_7_delay_11_52;
  reg                 io_A_Valid_7_delay_12_51;
  reg                 io_A_Valid_7_delay_13_50;
  reg                 io_A_Valid_7_delay_14_49;
  reg                 io_A_Valid_7_delay_15_48;
  reg                 io_A_Valid_7_delay_16_47;
  reg                 io_A_Valid_7_delay_17_46;
  reg                 io_A_Valid_7_delay_18_45;
  reg                 io_A_Valid_7_delay_19_44;
  reg                 io_A_Valid_7_delay_20_43;
  reg                 io_A_Valid_7_delay_21_42;
  reg                 io_A_Valid_7_delay_22_41;
  reg                 io_A_Valid_7_delay_23_40;
  reg                 io_A_Valid_7_delay_24_39;
  reg                 io_A_Valid_7_delay_25_38;
  reg                 io_A_Valid_7_delay_26_37;
  reg                 io_A_Valid_7_delay_27_36;
  reg                 io_A_Valid_7_delay_28_35;
  reg                 io_A_Valid_7_delay_29_34;
  reg                 io_A_Valid_7_delay_30_33;
  reg                 io_A_Valid_7_delay_31_32;
  reg                 io_A_Valid_7_delay_32_31;
  reg                 io_A_Valid_7_delay_33_30;
  reg                 io_A_Valid_7_delay_34_29;
  reg                 io_A_Valid_7_delay_35_28;
  reg                 io_A_Valid_7_delay_36_27;
  reg                 io_A_Valid_7_delay_37_26;
  reg                 io_A_Valid_7_delay_38_25;
  reg                 io_A_Valid_7_delay_39_24;
  reg                 io_A_Valid_7_delay_40_23;
  reg                 io_A_Valid_7_delay_41_22;
  reg                 io_A_Valid_7_delay_42_21;
  reg                 io_A_Valid_7_delay_43_20;
  reg                 io_A_Valid_7_delay_44_19;
  reg                 io_A_Valid_7_delay_45_18;
  reg                 io_A_Valid_7_delay_46_17;
  reg                 io_A_Valid_7_delay_47_16;
  reg                 io_A_Valid_7_delay_48_15;
  reg                 io_A_Valid_7_delay_49_14;
  reg                 io_A_Valid_7_delay_50_13;
  reg                 io_A_Valid_7_delay_51_12;
  reg                 io_A_Valid_7_delay_52_11;
  reg                 io_A_Valid_7_delay_53_10;
  reg                 io_A_Valid_7_delay_54_9;
  reg                 io_A_Valid_7_delay_55_8;
  reg                 io_A_Valid_7_delay_56_7;
  reg                 io_A_Valid_7_delay_57_6;
  reg                 io_A_Valid_7_delay_58_5;
  reg                 io_A_Valid_7_delay_59_4;
  reg                 io_A_Valid_7_delay_60_3;
  reg                 io_A_Valid_7_delay_61_2;
  reg                 io_A_Valid_7_delay_62_1;
  reg                 io_A_Valid_7_delay_63;
  reg                 io_B_Valid_63_delay_1_6;
  reg                 io_B_Valid_63_delay_2_5;
  reg                 io_B_Valid_63_delay_3_4;
  reg                 io_B_Valid_63_delay_4_3;
  reg                 io_B_Valid_63_delay_5_2;
  reg                 io_B_Valid_63_delay_6_1;
  reg                 io_B_Valid_63_delay_7;

  PE PE00 (
    .activate  (io_MatrixA_0[7:0]             ), //i
    .weight    (io_MatrixB_0[7:0]             ), //i
    .valid     (PE00_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE00_acount[7:0]              ), //o
    .bcount    (PE00_bcount[7:0]              ), //o
    .PE_OUT    (PE00_PE_OUT[31:0]             ), //o
    .finish    (PE00_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE01 (
    .activate  (PE00_acount[7:0]              ), //i
    .weight    (io_MatrixB_1[7:0]             ), //i
    .valid     (PE01_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE01_acount[7:0]              ), //o
    .bcount    (PE01_bcount[7:0]              ), //o
    .PE_OUT    (PE01_PE_OUT[31:0]             ), //o
    .finish    (PE01_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE02 (
    .activate  (PE01_acount[7:0]              ), //i
    .weight    (io_MatrixB_2[7:0]             ), //i
    .valid     (PE02_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE02_acount[7:0]              ), //o
    .bcount    (PE02_bcount[7:0]              ), //o
    .PE_OUT    (PE02_PE_OUT[31:0]             ), //o
    .finish    (PE02_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE03 (
    .activate  (PE02_acount[7:0]              ), //i
    .weight    (io_MatrixB_3[7:0]             ), //i
    .valid     (PE03_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE03_acount[7:0]              ), //o
    .bcount    (PE03_bcount[7:0]              ), //o
    .PE_OUT    (PE03_PE_OUT[31:0]             ), //o
    .finish    (PE03_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE04 (
    .activate  (PE03_acount[7:0]              ), //i
    .weight    (io_MatrixB_4[7:0]             ), //i
    .valid     (PE04_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE04_acount[7:0]              ), //o
    .bcount    (PE04_bcount[7:0]              ), //o
    .PE_OUT    (PE04_PE_OUT[31:0]             ), //o
    .finish    (PE04_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE05 (
    .activate  (PE04_acount[7:0]              ), //i
    .weight    (io_MatrixB_5[7:0]             ), //i
    .valid     (PE05_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE05_acount[7:0]              ), //o
    .bcount    (PE05_bcount[7:0]              ), //o
    .PE_OUT    (PE05_PE_OUT[31:0]             ), //o
    .finish    (PE05_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE06 (
    .activate  (PE05_acount[7:0]              ), //i
    .weight    (io_MatrixB_6[7:0]             ), //i
    .valid     (PE06_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE06_acount[7:0]              ), //o
    .bcount    (PE06_bcount[7:0]              ), //o
    .PE_OUT    (PE06_PE_OUT[31:0]             ), //o
    .finish    (PE06_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE07 (
    .activate  (PE06_acount[7:0]              ), //i
    .weight    (io_MatrixB_7[7:0]             ), //i
    .valid     (PE07_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE07_acount[7:0]              ), //o
    .bcount    (PE07_bcount[7:0]              ), //o
    .PE_OUT    (PE07_PE_OUT[31:0]             ), //o
    .finish    (PE07_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE08 (
    .activate  (PE07_acount[7:0]              ), //i
    .weight    (io_MatrixB_8[7:0]             ), //i
    .valid     (PE08_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE08_acount[7:0]              ), //o
    .bcount    (PE08_bcount[7:0]              ), //o
    .PE_OUT    (PE08_PE_OUT[31:0]             ), //o
    .finish    (PE08_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE09 (
    .activate  (PE08_acount[7:0]              ), //i
    .weight    (io_MatrixB_9[7:0]             ), //i
    .valid     (PE09_valid                    ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE09_acount[7:0]              ), //o
    .bcount    (PE09_bcount[7:0]              ), //o
    .PE_OUT    (PE09_PE_OUT[31:0]             ), //o
    .finish    (PE09_finish                   ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE010 (
    .activate  (PE09_acount[7:0]              ), //i
    .weight    (io_MatrixB_10[7:0]            ), //i
    .valid     (PE010_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE010_acount[7:0]             ), //o
    .bcount    (PE010_bcount[7:0]             ), //o
    .PE_OUT    (PE010_PE_OUT[31:0]            ), //o
    .finish    (PE010_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE011 (
    .activate  (PE010_acount[7:0]             ), //i
    .weight    (io_MatrixB_11[7:0]            ), //i
    .valid     (PE011_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE011_acount[7:0]             ), //o
    .bcount    (PE011_bcount[7:0]             ), //o
    .PE_OUT    (PE011_PE_OUT[31:0]            ), //o
    .finish    (PE011_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE012 (
    .activate  (PE011_acount[7:0]             ), //i
    .weight    (io_MatrixB_12[7:0]            ), //i
    .valid     (PE012_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE012_acount[7:0]             ), //o
    .bcount    (PE012_bcount[7:0]             ), //o
    .PE_OUT    (PE012_PE_OUT[31:0]            ), //o
    .finish    (PE012_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE013 (
    .activate  (PE012_acount[7:0]             ), //i
    .weight    (io_MatrixB_13[7:0]            ), //i
    .valid     (PE013_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE013_acount[7:0]             ), //o
    .bcount    (PE013_bcount[7:0]             ), //o
    .PE_OUT    (PE013_PE_OUT[31:0]            ), //o
    .finish    (PE013_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE014 (
    .activate  (PE013_acount[7:0]             ), //i
    .weight    (io_MatrixB_14[7:0]            ), //i
    .valid     (PE014_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE014_acount[7:0]             ), //o
    .bcount    (PE014_bcount[7:0]             ), //o
    .PE_OUT    (PE014_PE_OUT[31:0]            ), //o
    .finish    (PE014_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE015 (
    .activate  (PE014_acount[7:0]             ), //i
    .weight    (io_MatrixB_15[7:0]            ), //i
    .valid     (PE015_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE015_acount[7:0]             ), //o
    .bcount    (PE015_bcount[7:0]             ), //o
    .PE_OUT    (PE015_PE_OUT[31:0]            ), //o
    .finish    (PE015_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE016 (
    .activate  (PE015_acount[7:0]             ), //i
    .weight    (io_MatrixB_16[7:0]            ), //i
    .valid     (PE016_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE016_acount[7:0]             ), //o
    .bcount    (PE016_bcount[7:0]             ), //o
    .PE_OUT    (PE016_PE_OUT[31:0]            ), //o
    .finish    (PE016_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE017 (
    .activate  (PE016_acount[7:0]             ), //i
    .weight    (io_MatrixB_17[7:0]            ), //i
    .valid     (PE017_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE017_acount[7:0]             ), //o
    .bcount    (PE017_bcount[7:0]             ), //o
    .PE_OUT    (PE017_PE_OUT[31:0]            ), //o
    .finish    (PE017_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE018 (
    .activate  (PE017_acount[7:0]             ), //i
    .weight    (io_MatrixB_18[7:0]            ), //i
    .valid     (PE018_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE018_acount[7:0]             ), //o
    .bcount    (PE018_bcount[7:0]             ), //o
    .PE_OUT    (PE018_PE_OUT[31:0]            ), //o
    .finish    (PE018_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE019 (
    .activate  (PE018_acount[7:0]             ), //i
    .weight    (io_MatrixB_19[7:0]            ), //i
    .valid     (PE019_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE019_acount[7:0]             ), //o
    .bcount    (PE019_bcount[7:0]             ), //o
    .PE_OUT    (PE019_PE_OUT[31:0]            ), //o
    .finish    (PE019_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE020 (
    .activate  (PE019_acount[7:0]             ), //i
    .weight    (io_MatrixB_20[7:0]            ), //i
    .valid     (PE020_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE020_acount[7:0]             ), //o
    .bcount    (PE020_bcount[7:0]             ), //o
    .PE_OUT    (PE020_PE_OUT[31:0]            ), //o
    .finish    (PE020_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE021 (
    .activate  (PE020_acount[7:0]             ), //i
    .weight    (io_MatrixB_21[7:0]            ), //i
    .valid     (PE021_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE021_acount[7:0]             ), //o
    .bcount    (PE021_bcount[7:0]             ), //o
    .PE_OUT    (PE021_PE_OUT[31:0]            ), //o
    .finish    (PE021_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE022 (
    .activate  (PE021_acount[7:0]             ), //i
    .weight    (io_MatrixB_22[7:0]            ), //i
    .valid     (PE022_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE022_acount[7:0]             ), //o
    .bcount    (PE022_bcount[7:0]             ), //o
    .PE_OUT    (PE022_PE_OUT[31:0]            ), //o
    .finish    (PE022_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE023 (
    .activate  (PE022_acount[7:0]             ), //i
    .weight    (io_MatrixB_23[7:0]            ), //i
    .valid     (PE023_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE023_acount[7:0]             ), //o
    .bcount    (PE023_bcount[7:0]             ), //o
    .PE_OUT    (PE023_PE_OUT[31:0]            ), //o
    .finish    (PE023_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE024 (
    .activate  (PE023_acount[7:0]             ), //i
    .weight    (io_MatrixB_24[7:0]            ), //i
    .valid     (PE024_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE024_acount[7:0]             ), //o
    .bcount    (PE024_bcount[7:0]             ), //o
    .PE_OUT    (PE024_PE_OUT[31:0]            ), //o
    .finish    (PE024_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE025 (
    .activate  (PE024_acount[7:0]             ), //i
    .weight    (io_MatrixB_25[7:0]            ), //i
    .valid     (PE025_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE025_acount[7:0]             ), //o
    .bcount    (PE025_bcount[7:0]             ), //o
    .PE_OUT    (PE025_PE_OUT[31:0]            ), //o
    .finish    (PE025_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE026 (
    .activate  (PE025_acount[7:0]             ), //i
    .weight    (io_MatrixB_26[7:0]            ), //i
    .valid     (PE026_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE026_acount[7:0]             ), //o
    .bcount    (PE026_bcount[7:0]             ), //o
    .PE_OUT    (PE026_PE_OUT[31:0]            ), //o
    .finish    (PE026_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE027 (
    .activate  (PE026_acount[7:0]             ), //i
    .weight    (io_MatrixB_27[7:0]            ), //i
    .valid     (PE027_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE027_acount[7:0]             ), //o
    .bcount    (PE027_bcount[7:0]             ), //o
    .PE_OUT    (PE027_PE_OUT[31:0]            ), //o
    .finish    (PE027_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE028 (
    .activate  (PE027_acount[7:0]             ), //i
    .weight    (io_MatrixB_28[7:0]            ), //i
    .valid     (PE028_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE028_acount[7:0]             ), //o
    .bcount    (PE028_bcount[7:0]             ), //o
    .PE_OUT    (PE028_PE_OUT[31:0]            ), //o
    .finish    (PE028_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE029 (
    .activate  (PE028_acount[7:0]             ), //i
    .weight    (io_MatrixB_29[7:0]            ), //i
    .valid     (PE029_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE029_acount[7:0]             ), //o
    .bcount    (PE029_bcount[7:0]             ), //o
    .PE_OUT    (PE029_PE_OUT[31:0]            ), //o
    .finish    (PE029_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE030 (
    .activate  (PE029_acount[7:0]             ), //i
    .weight    (io_MatrixB_30[7:0]            ), //i
    .valid     (PE030_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE030_acount[7:0]             ), //o
    .bcount    (PE030_bcount[7:0]             ), //o
    .PE_OUT    (PE030_PE_OUT[31:0]            ), //o
    .finish    (PE030_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE031 (
    .activate  (PE030_acount[7:0]             ), //i
    .weight    (io_MatrixB_31[7:0]            ), //i
    .valid     (PE031_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE031_acount[7:0]             ), //o
    .bcount    (PE031_bcount[7:0]             ), //o
    .PE_OUT    (PE031_PE_OUT[31:0]            ), //o
    .finish    (PE031_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE032 (
    .activate  (PE031_acount[7:0]             ), //i
    .weight    (io_MatrixB_32[7:0]            ), //i
    .valid     (PE032_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE032_acount[7:0]             ), //o
    .bcount    (PE032_bcount[7:0]             ), //o
    .PE_OUT    (PE032_PE_OUT[31:0]            ), //o
    .finish    (PE032_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE033 (
    .activate  (PE032_acount[7:0]             ), //i
    .weight    (io_MatrixB_33[7:0]            ), //i
    .valid     (PE033_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE033_acount[7:0]             ), //o
    .bcount    (PE033_bcount[7:0]             ), //o
    .PE_OUT    (PE033_PE_OUT[31:0]            ), //o
    .finish    (PE033_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE034 (
    .activate  (PE033_acount[7:0]             ), //i
    .weight    (io_MatrixB_34[7:0]            ), //i
    .valid     (PE034_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE034_acount[7:0]             ), //o
    .bcount    (PE034_bcount[7:0]             ), //o
    .PE_OUT    (PE034_PE_OUT[31:0]            ), //o
    .finish    (PE034_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE035 (
    .activate  (PE034_acount[7:0]             ), //i
    .weight    (io_MatrixB_35[7:0]            ), //i
    .valid     (PE035_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE035_acount[7:0]             ), //o
    .bcount    (PE035_bcount[7:0]             ), //o
    .PE_OUT    (PE035_PE_OUT[31:0]            ), //o
    .finish    (PE035_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE036 (
    .activate  (PE035_acount[7:0]             ), //i
    .weight    (io_MatrixB_36[7:0]            ), //i
    .valid     (PE036_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE036_acount[7:0]             ), //o
    .bcount    (PE036_bcount[7:0]             ), //o
    .PE_OUT    (PE036_PE_OUT[31:0]            ), //o
    .finish    (PE036_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE037 (
    .activate  (PE036_acount[7:0]             ), //i
    .weight    (io_MatrixB_37[7:0]            ), //i
    .valid     (PE037_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE037_acount[7:0]             ), //o
    .bcount    (PE037_bcount[7:0]             ), //o
    .PE_OUT    (PE037_PE_OUT[31:0]            ), //o
    .finish    (PE037_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE038 (
    .activate  (PE037_acount[7:0]             ), //i
    .weight    (io_MatrixB_38[7:0]            ), //i
    .valid     (PE038_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE038_acount[7:0]             ), //o
    .bcount    (PE038_bcount[7:0]             ), //o
    .PE_OUT    (PE038_PE_OUT[31:0]            ), //o
    .finish    (PE038_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE039 (
    .activate  (PE038_acount[7:0]             ), //i
    .weight    (io_MatrixB_39[7:0]            ), //i
    .valid     (PE039_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE039_acount[7:0]             ), //o
    .bcount    (PE039_bcount[7:0]             ), //o
    .PE_OUT    (PE039_PE_OUT[31:0]            ), //o
    .finish    (PE039_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE040 (
    .activate  (PE039_acount[7:0]             ), //i
    .weight    (io_MatrixB_40[7:0]            ), //i
    .valid     (PE040_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE040_acount[7:0]             ), //o
    .bcount    (PE040_bcount[7:0]             ), //o
    .PE_OUT    (PE040_PE_OUT[31:0]            ), //o
    .finish    (PE040_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE041 (
    .activate  (PE040_acount[7:0]             ), //i
    .weight    (io_MatrixB_41[7:0]            ), //i
    .valid     (PE041_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE041_acount[7:0]             ), //o
    .bcount    (PE041_bcount[7:0]             ), //o
    .PE_OUT    (PE041_PE_OUT[31:0]            ), //o
    .finish    (PE041_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE042 (
    .activate  (PE041_acount[7:0]             ), //i
    .weight    (io_MatrixB_42[7:0]            ), //i
    .valid     (PE042_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE042_acount[7:0]             ), //o
    .bcount    (PE042_bcount[7:0]             ), //o
    .PE_OUT    (PE042_PE_OUT[31:0]            ), //o
    .finish    (PE042_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE043 (
    .activate  (PE042_acount[7:0]             ), //i
    .weight    (io_MatrixB_43[7:0]            ), //i
    .valid     (PE043_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE043_acount[7:0]             ), //o
    .bcount    (PE043_bcount[7:0]             ), //o
    .PE_OUT    (PE043_PE_OUT[31:0]            ), //o
    .finish    (PE043_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE044 (
    .activate  (PE043_acount[7:0]             ), //i
    .weight    (io_MatrixB_44[7:0]            ), //i
    .valid     (PE044_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE044_acount[7:0]             ), //o
    .bcount    (PE044_bcount[7:0]             ), //o
    .PE_OUT    (PE044_PE_OUT[31:0]            ), //o
    .finish    (PE044_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE045 (
    .activate  (PE044_acount[7:0]             ), //i
    .weight    (io_MatrixB_45[7:0]            ), //i
    .valid     (PE045_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE045_acount[7:0]             ), //o
    .bcount    (PE045_bcount[7:0]             ), //o
    .PE_OUT    (PE045_PE_OUT[31:0]            ), //o
    .finish    (PE045_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE046 (
    .activate  (PE045_acount[7:0]             ), //i
    .weight    (io_MatrixB_46[7:0]            ), //i
    .valid     (PE046_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE046_acount[7:0]             ), //o
    .bcount    (PE046_bcount[7:0]             ), //o
    .PE_OUT    (PE046_PE_OUT[31:0]            ), //o
    .finish    (PE046_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE047 (
    .activate  (PE046_acount[7:0]             ), //i
    .weight    (io_MatrixB_47[7:0]            ), //i
    .valid     (PE047_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE047_acount[7:0]             ), //o
    .bcount    (PE047_bcount[7:0]             ), //o
    .PE_OUT    (PE047_PE_OUT[31:0]            ), //o
    .finish    (PE047_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE048 (
    .activate  (PE047_acount[7:0]             ), //i
    .weight    (io_MatrixB_48[7:0]            ), //i
    .valid     (PE048_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE048_acount[7:0]             ), //o
    .bcount    (PE048_bcount[7:0]             ), //o
    .PE_OUT    (PE048_PE_OUT[31:0]            ), //o
    .finish    (PE048_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE049 (
    .activate  (PE048_acount[7:0]             ), //i
    .weight    (io_MatrixB_49[7:0]            ), //i
    .valid     (PE049_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE049_acount[7:0]             ), //o
    .bcount    (PE049_bcount[7:0]             ), //o
    .PE_OUT    (PE049_PE_OUT[31:0]            ), //o
    .finish    (PE049_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE050 (
    .activate  (PE049_acount[7:0]             ), //i
    .weight    (io_MatrixB_50[7:0]            ), //i
    .valid     (PE050_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE050_acount[7:0]             ), //o
    .bcount    (PE050_bcount[7:0]             ), //o
    .PE_OUT    (PE050_PE_OUT[31:0]            ), //o
    .finish    (PE050_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE051 (
    .activate  (PE050_acount[7:0]             ), //i
    .weight    (io_MatrixB_51[7:0]            ), //i
    .valid     (PE051_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE051_acount[7:0]             ), //o
    .bcount    (PE051_bcount[7:0]             ), //o
    .PE_OUT    (PE051_PE_OUT[31:0]            ), //o
    .finish    (PE051_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE052 (
    .activate  (PE051_acount[7:0]             ), //i
    .weight    (io_MatrixB_52[7:0]            ), //i
    .valid     (PE052_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE052_acount[7:0]             ), //o
    .bcount    (PE052_bcount[7:0]             ), //o
    .PE_OUT    (PE052_PE_OUT[31:0]            ), //o
    .finish    (PE052_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE053 (
    .activate  (PE052_acount[7:0]             ), //i
    .weight    (io_MatrixB_53[7:0]            ), //i
    .valid     (PE053_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE053_acount[7:0]             ), //o
    .bcount    (PE053_bcount[7:0]             ), //o
    .PE_OUT    (PE053_PE_OUT[31:0]            ), //o
    .finish    (PE053_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE054 (
    .activate  (PE053_acount[7:0]             ), //i
    .weight    (io_MatrixB_54[7:0]            ), //i
    .valid     (PE054_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE054_acount[7:0]             ), //o
    .bcount    (PE054_bcount[7:0]             ), //o
    .PE_OUT    (PE054_PE_OUT[31:0]            ), //o
    .finish    (PE054_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE055 (
    .activate  (PE054_acount[7:0]             ), //i
    .weight    (io_MatrixB_55[7:0]            ), //i
    .valid     (PE055_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE055_acount[7:0]             ), //o
    .bcount    (PE055_bcount[7:0]             ), //o
    .PE_OUT    (PE055_PE_OUT[31:0]            ), //o
    .finish    (PE055_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE056 (
    .activate  (PE055_acount[7:0]             ), //i
    .weight    (io_MatrixB_56[7:0]            ), //i
    .valid     (PE056_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE056_acount[7:0]             ), //o
    .bcount    (PE056_bcount[7:0]             ), //o
    .PE_OUT    (PE056_PE_OUT[31:0]            ), //o
    .finish    (PE056_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE057 (
    .activate  (PE056_acount[7:0]             ), //i
    .weight    (io_MatrixB_57[7:0]            ), //i
    .valid     (PE057_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE057_acount[7:0]             ), //o
    .bcount    (PE057_bcount[7:0]             ), //o
    .PE_OUT    (PE057_PE_OUT[31:0]            ), //o
    .finish    (PE057_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE058 (
    .activate  (PE057_acount[7:0]             ), //i
    .weight    (io_MatrixB_58[7:0]            ), //i
    .valid     (PE058_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE058_acount[7:0]             ), //o
    .bcount    (PE058_bcount[7:0]             ), //o
    .PE_OUT    (PE058_PE_OUT[31:0]            ), //o
    .finish    (PE058_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE059 (
    .activate  (PE058_acount[7:0]             ), //i
    .weight    (io_MatrixB_59[7:0]            ), //i
    .valid     (PE059_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE059_acount[7:0]             ), //o
    .bcount    (PE059_bcount[7:0]             ), //o
    .PE_OUT    (PE059_PE_OUT[31:0]            ), //o
    .finish    (PE059_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE060 (
    .activate  (PE059_acount[7:0]             ), //i
    .weight    (io_MatrixB_60[7:0]            ), //i
    .valid     (PE060_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE060_acount[7:0]             ), //o
    .bcount    (PE060_bcount[7:0]             ), //o
    .PE_OUT    (PE060_PE_OUT[31:0]            ), //o
    .finish    (PE060_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE061 (
    .activate  (PE060_acount[7:0]             ), //i
    .weight    (io_MatrixB_61[7:0]            ), //i
    .valid     (PE061_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE061_acount[7:0]             ), //o
    .bcount    (PE061_bcount[7:0]             ), //o
    .PE_OUT    (PE061_PE_OUT[31:0]            ), //o
    .finish    (PE061_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE062 (
    .activate  (PE061_acount[7:0]             ), //i
    .weight    (io_MatrixB_62[7:0]            ), //i
    .valid     (PE062_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE062_acount[7:0]             ), //o
    .bcount    (PE062_bcount[7:0]             ), //o
    .PE_OUT    (PE062_PE_OUT[31:0]            ), //o
    .finish    (PE062_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE063 (
    .activate  (PE062_acount[7:0]             ), //i
    .weight    (io_MatrixB_63[7:0]            ), //i
    .valid     (PE063_valid                   ), //i
    .signCount (io_signCount_regNextWhen[15:0]), //i
    .acount    (PE063_acount[7:0]             ), //o
    .bcount    (PE063_bcount[7:0]             ), //o
    .PE_OUT    (PE063_PE_OUT[31:0]            ), //o
    .finish    (PE063_finish                  ), //o
    .clk       (clk                           ), //i
    .reset     (reset                         )  //i
  );
  PE PE10 (
    .activate  (io_MatrixA_1[7:0]               ), //i
    .weight    (PE00_bcount[7:0]                ), //i
    .valid     (PE10_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE10_acount[7:0]                ), //o
    .bcount    (PE10_bcount[7:0]                ), //o
    .PE_OUT    (PE10_PE_OUT[31:0]               ), //o
    .finish    (PE10_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE11 (
    .activate  (PE10_acount[7:0]                ), //i
    .weight    (PE01_bcount[7:0]                ), //i
    .valid     (PE11_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE11_acount[7:0]                ), //o
    .bcount    (PE11_bcount[7:0]                ), //o
    .PE_OUT    (PE11_PE_OUT[31:0]               ), //o
    .finish    (PE11_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE12 (
    .activate  (PE11_acount[7:0]                ), //i
    .weight    (PE02_bcount[7:0]                ), //i
    .valid     (PE12_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE12_acount[7:0]                ), //o
    .bcount    (PE12_bcount[7:0]                ), //o
    .PE_OUT    (PE12_PE_OUT[31:0]               ), //o
    .finish    (PE12_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE13 (
    .activate  (PE12_acount[7:0]                ), //i
    .weight    (PE03_bcount[7:0]                ), //i
    .valid     (PE13_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE13_acount[7:0]                ), //o
    .bcount    (PE13_bcount[7:0]                ), //o
    .PE_OUT    (PE13_PE_OUT[31:0]               ), //o
    .finish    (PE13_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE14 (
    .activate  (PE13_acount[7:0]                ), //i
    .weight    (PE04_bcount[7:0]                ), //i
    .valid     (PE14_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE14_acount[7:0]                ), //o
    .bcount    (PE14_bcount[7:0]                ), //o
    .PE_OUT    (PE14_PE_OUT[31:0]               ), //o
    .finish    (PE14_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE15 (
    .activate  (PE14_acount[7:0]                ), //i
    .weight    (PE05_bcount[7:0]                ), //i
    .valid     (PE15_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE15_acount[7:0]                ), //o
    .bcount    (PE15_bcount[7:0]                ), //o
    .PE_OUT    (PE15_PE_OUT[31:0]               ), //o
    .finish    (PE15_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE16 (
    .activate  (PE15_acount[7:0]                ), //i
    .weight    (PE06_bcount[7:0]                ), //i
    .valid     (PE16_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE16_acount[7:0]                ), //o
    .bcount    (PE16_bcount[7:0]                ), //o
    .PE_OUT    (PE16_PE_OUT[31:0]               ), //o
    .finish    (PE16_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE17 (
    .activate  (PE16_acount[7:0]                ), //i
    .weight    (PE07_bcount[7:0]                ), //i
    .valid     (PE17_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE17_acount[7:0]                ), //o
    .bcount    (PE17_bcount[7:0]                ), //o
    .PE_OUT    (PE17_PE_OUT[31:0]               ), //o
    .finish    (PE17_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE18 (
    .activate  (PE17_acount[7:0]                ), //i
    .weight    (PE08_bcount[7:0]                ), //i
    .valid     (PE18_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE18_acount[7:0]                ), //o
    .bcount    (PE18_bcount[7:0]                ), //o
    .PE_OUT    (PE18_PE_OUT[31:0]               ), //o
    .finish    (PE18_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE19 (
    .activate  (PE18_acount[7:0]                ), //i
    .weight    (PE09_bcount[7:0]                ), //i
    .valid     (PE19_valid                      ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE19_acount[7:0]                ), //o
    .bcount    (PE19_bcount[7:0]                ), //o
    .PE_OUT    (PE19_PE_OUT[31:0]               ), //o
    .finish    (PE19_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE110 (
    .activate  (PE19_acount[7:0]                ), //i
    .weight    (PE010_bcount[7:0]               ), //i
    .valid     (PE110_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE110_acount[7:0]               ), //o
    .bcount    (PE110_bcount[7:0]               ), //o
    .PE_OUT    (PE110_PE_OUT[31:0]              ), //o
    .finish    (PE110_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE111 (
    .activate  (PE110_acount[7:0]               ), //i
    .weight    (PE011_bcount[7:0]               ), //i
    .valid     (PE111_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE111_acount[7:0]               ), //o
    .bcount    (PE111_bcount[7:0]               ), //o
    .PE_OUT    (PE111_PE_OUT[31:0]              ), //o
    .finish    (PE111_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE112 (
    .activate  (PE111_acount[7:0]               ), //i
    .weight    (PE012_bcount[7:0]               ), //i
    .valid     (PE112_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE112_acount[7:0]               ), //o
    .bcount    (PE112_bcount[7:0]               ), //o
    .PE_OUT    (PE112_PE_OUT[31:0]              ), //o
    .finish    (PE112_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE113 (
    .activate  (PE112_acount[7:0]               ), //i
    .weight    (PE013_bcount[7:0]               ), //i
    .valid     (PE113_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE113_acount[7:0]               ), //o
    .bcount    (PE113_bcount[7:0]               ), //o
    .PE_OUT    (PE113_PE_OUT[31:0]              ), //o
    .finish    (PE113_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE114 (
    .activate  (PE113_acount[7:0]               ), //i
    .weight    (PE014_bcount[7:0]               ), //i
    .valid     (PE114_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE114_acount[7:0]               ), //o
    .bcount    (PE114_bcount[7:0]               ), //o
    .PE_OUT    (PE114_PE_OUT[31:0]              ), //o
    .finish    (PE114_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE115 (
    .activate  (PE114_acount[7:0]               ), //i
    .weight    (PE015_bcount[7:0]               ), //i
    .valid     (PE115_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE115_acount[7:0]               ), //o
    .bcount    (PE115_bcount[7:0]               ), //o
    .PE_OUT    (PE115_PE_OUT[31:0]              ), //o
    .finish    (PE115_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE116 (
    .activate  (PE115_acount[7:0]               ), //i
    .weight    (PE016_bcount[7:0]               ), //i
    .valid     (PE116_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE116_acount[7:0]               ), //o
    .bcount    (PE116_bcount[7:0]               ), //o
    .PE_OUT    (PE116_PE_OUT[31:0]              ), //o
    .finish    (PE116_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE117 (
    .activate  (PE116_acount[7:0]               ), //i
    .weight    (PE017_bcount[7:0]               ), //i
    .valid     (PE117_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE117_acount[7:0]               ), //o
    .bcount    (PE117_bcount[7:0]               ), //o
    .PE_OUT    (PE117_PE_OUT[31:0]              ), //o
    .finish    (PE117_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE118 (
    .activate  (PE117_acount[7:0]               ), //i
    .weight    (PE018_bcount[7:0]               ), //i
    .valid     (PE118_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE118_acount[7:0]               ), //o
    .bcount    (PE118_bcount[7:0]               ), //o
    .PE_OUT    (PE118_PE_OUT[31:0]              ), //o
    .finish    (PE118_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE119 (
    .activate  (PE118_acount[7:0]               ), //i
    .weight    (PE019_bcount[7:0]               ), //i
    .valid     (PE119_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE119_acount[7:0]               ), //o
    .bcount    (PE119_bcount[7:0]               ), //o
    .PE_OUT    (PE119_PE_OUT[31:0]              ), //o
    .finish    (PE119_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE120 (
    .activate  (PE119_acount[7:0]               ), //i
    .weight    (PE020_bcount[7:0]               ), //i
    .valid     (PE120_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE120_acount[7:0]               ), //o
    .bcount    (PE120_bcount[7:0]               ), //o
    .PE_OUT    (PE120_PE_OUT[31:0]              ), //o
    .finish    (PE120_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE121 (
    .activate  (PE120_acount[7:0]               ), //i
    .weight    (PE021_bcount[7:0]               ), //i
    .valid     (PE121_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE121_acount[7:0]               ), //o
    .bcount    (PE121_bcount[7:0]               ), //o
    .PE_OUT    (PE121_PE_OUT[31:0]              ), //o
    .finish    (PE121_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE122 (
    .activate  (PE121_acount[7:0]               ), //i
    .weight    (PE022_bcount[7:0]               ), //i
    .valid     (PE122_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE122_acount[7:0]               ), //o
    .bcount    (PE122_bcount[7:0]               ), //o
    .PE_OUT    (PE122_PE_OUT[31:0]              ), //o
    .finish    (PE122_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE123 (
    .activate  (PE122_acount[7:0]               ), //i
    .weight    (PE023_bcount[7:0]               ), //i
    .valid     (PE123_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE123_acount[7:0]               ), //o
    .bcount    (PE123_bcount[7:0]               ), //o
    .PE_OUT    (PE123_PE_OUT[31:0]              ), //o
    .finish    (PE123_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE124 (
    .activate  (PE123_acount[7:0]               ), //i
    .weight    (PE024_bcount[7:0]               ), //i
    .valid     (PE124_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE124_acount[7:0]               ), //o
    .bcount    (PE124_bcount[7:0]               ), //o
    .PE_OUT    (PE124_PE_OUT[31:0]              ), //o
    .finish    (PE124_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE125 (
    .activate  (PE124_acount[7:0]               ), //i
    .weight    (PE025_bcount[7:0]               ), //i
    .valid     (PE125_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE125_acount[7:0]               ), //o
    .bcount    (PE125_bcount[7:0]               ), //o
    .PE_OUT    (PE125_PE_OUT[31:0]              ), //o
    .finish    (PE125_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE126 (
    .activate  (PE125_acount[7:0]               ), //i
    .weight    (PE026_bcount[7:0]               ), //i
    .valid     (PE126_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE126_acount[7:0]               ), //o
    .bcount    (PE126_bcount[7:0]               ), //o
    .PE_OUT    (PE126_PE_OUT[31:0]              ), //o
    .finish    (PE126_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE127 (
    .activate  (PE126_acount[7:0]               ), //i
    .weight    (PE027_bcount[7:0]               ), //i
    .valid     (PE127_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE127_acount[7:0]               ), //o
    .bcount    (PE127_bcount[7:0]               ), //o
    .PE_OUT    (PE127_PE_OUT[31:0]              ), //o
    .finish    (PE127_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE128 (
    .activate  (PE127_acount[7:0]               ), //i
    .weight    (PE028_bcount[7:0]               ), //i
    .valid     (PE128_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE128_acount[7:0]               ), //o
    .bcount    (PE128_bcount[7:0]               ), //o
    .PE_OUT    (PE128_PE_OUT[31:0]              ), //o
    .finish    (PE128_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE129 (
    .activate  (PE128_acount[7:0]               ), //i
    .weight    (PE029_bcount[7:0]               ), //i
    .valid     (PE129_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE129_acount[7:0]               ), //o
    .bcount    (PE129_bcount[7:0]               ), //o
    .PE_OUT    (PE129_PE_OUT[31:0]              ), //o
    .finish    (PE129_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE130 (
    .activate  (PE129_acount[7:0]               ), //i
    .weight    (PE030_bcount[7:0]               ), //i
    .valid     (PE130_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE130_acount[7:0]               ), //o
    .bcount    (PE130_bcount[7:0]               ), //o
    .PE_OUT    (PE130_PE_OUT[31:0]              ), //o
    .finish    (PE130_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE131 (
    .activate  (PE130_acount[7:0]               ), //i
    .weight    (PE031_bcount[7:0]               ), //i
    .valid     (PE131_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE131_acount[7:0]               ), //o
    .bcount    (PE131_bcount[7:0]               ), //o
    .PE_OUT    (PE131_PE_OUT[31:0]              ), //o
    .finish    (PE131_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE132 (
    .activate  (PE131_acount[7:0]               ), //i
    .weight    (PE032_bcount[7:0]               ), //i
    .valid     (PE132_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE132_acount[7:0]               ), //o
    .bcount    (PE132_bcount[7:0]               ), //o
    .PE_OUT    (PE132_PE_OUT[31:0]              ), //o
    .finish    (PE132_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE133 (
    .activate  (PE132_acount[7:0]               ), //i
    .weight    (PE033_bcount[7:0]               ), //i
    .valid     (PE133_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE133_acount[7:0]               ), //o
    .bcount    (PE133_bcount[7:0]               ), //o
    .PE_OUT    (PE133_PE_OUT[31:0]              ), //o
    .finish    (PE133_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE134 (
    .activate  (PE133_acount[7:0]               ), //i
    .weight    (PE034_bcount[7:0]               ), //i
    .valid     (PE134_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE134_acount[7:0]               ), //o
    .bcount    (PE134_bcount[7:0]               ), //o
    .PE_OUT    (PE134_PE_OUT[31:0]              ), //o
    .finish    (PE134_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE135 (
    .activate  (PE134_acount[7:0]               ), //i
    .weight    (PE035_bcount[7:0]               ), //i
    .valid     (PE135_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE135_acount[7:0]               ), //o
    .bcount    (PE135_bcount[7:0]               ), //o
    .PE_OUT    (PE135_PE_OUT[31:0]              ), //o
    .finish    (PE135_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE136 (
    .activate  (PE135_acount[7:0]               ), //i
    .weight    (PE036_bcount[7:0]               ), //i
    .valid     (PE136_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE136_acount[7:0]               ), //o
    .bcount    (PE136_bcount[7:0]               ), //o
    .PE_OUT    (PE136_PE_OUT[31:0]              ), //o
    .finish    (PE136_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE137 (
    .activate  (PE136_acount[7:0]               ), //i
    .weight    (PE037_bcount[7:0]               ), //i
    .valid     (PE137_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE137_acount[7:0]               ), //o
    .bcount    (PE137_bcount[7:0]               ), //o
    .PE_OUT    (PE137_PE_OUT[31:0]              ), //o
    .finish    (PE137_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE138 (
    .activate  (PE137_acount[7:0]               ), //i
    .weight    (PE038_bcount[7:0]               ), //i
    .valid     (PE138_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE138_acount[7:0]               ), //o
    .bcount    (PE138_bcount[7:0]               ), //o
    .PE_OUT    (PE138_PE_OUT[31:0]              ), //o
    .finish    (PE138_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE139 (
    .activate  (PE138_acount[7:0]               ), //i
    .weight    (PE039_bcount[7:0]               ), //i
    .valid     (PE139_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE139_acount[7:0]               ), //o
    .bcount    (PE139_bcount[7:0]               ), //o
    .PE_OUT    (PE139_PE_OUT[31:0]              ), //o
    .finish    (PE139_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE140 (
    .activate  (PE139_acount[7:0]               ), //i
    .weight    (PE040_bcount[7:0]               ), //i
    .valid     (PE140_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE140_acount[7:0]               ), //o
    .bcount    (PE140_bcount[7:0]               ), //o
    .PE_OUT    (PE140_PE_OUT[31:0]              ), //o
    .finish    (PE140_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE141 (
    .activate  (PE140_acount[7:0]               ), //i
    .weight    (PE041_bcount[7:0]               ), //i
    .valid     (PE141_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE141_acount[7:0]               ), //o
    .bcount    (PE141_bcount[7:0]               ), //o
    .PE_OUT    (PE141_PE_OUT[31:0]              ), //o
    .finish    (PE141_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE142 (
    .activate  (PE141_acount[7:0]               ), //i
    .weight    (PE042_bcount[7:0]               ), //i
    .valid     (PE142_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE142_acount[7:0]               ), //o
    .bcount    (PE142_bcount[7:0]               ), //o
    .PE_OUT    (PE142_PE_OUT[31:0]              ), //o
    .finish    (PE142_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE143 (
    .activate  (PE142_acount[7:0]               ), //i
    .weight    (PE043_bcount[7:0]               ), //i
    .valid     (PE143_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE143_acount[7:0]               ), //o
    .bcount    (PE143_bcount[7:0]               ), //o
    .PE_OUT    (PE143_PE_OUT[31:0]              ), //o
    .finish    (PE143_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE144 (
    .activate  (PE143_acount[7:0]               ), //i
    .weight    (PE044_bcount[7:0]               ), //i
    .valid     (PE144_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE144_acount[7:0]               ), //o
    .bcount    (PE144_bcount[7:0]               ), //o
    .PE_OUT    (PE144_PE_OUT[31:0]              ), //o
    .finish    (PE144_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE145 (
    .activate  (PE144_acount[7:0]               ), //i
    .weight    (PE045_bcount[7:0]               ), //i
    .valid     (PE145_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE145_acount[7:0]               ), //o
    .bcount    (PE145_bcount[7:0]               ), //o
    .PE_OUT    (PE145_PE_OUT[31:0]              ), //o
    .finish    (PE145_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE146 (
    .activate  (PE145_acount[7:0]               ), //i
    .weight    (PE046_bcount[7:0]               ), //i
    .valid     (PE146_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE146_acount[7:0]               ), //o
    .bcount    (PE146_bcount[7:0]               ), //o
    .PE_OUT    (PE146_PE_OUT[31:0]              ), //o
    .finish    (PE146_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE147 (
    .activate  (PE146_acount[7:0]               ), //i
    .weight    (PE047_bcount[7:0]               ), //i
    .valid     (PE147_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE147_acount[7:0]               ), //o
    .bcount    (PE147_bcount[7:0]               ), //o
    .PE_OUT    (PE147_PE_OUT[31:0]              ), //o
    .finish    (PE147_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE148 (
    .activate  (PE147_acount[7:0]               ), //i
    .weight    (PE048_bcount[7:0]               ), //i
    .valid     (PE148_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE148_acount[7:0]               ), //o
    .bcount    (PE148_bcount[7:0]               ), //o
    .PE_OUT    (PE148_PE_OUT[31:0]              ), //o
    .finish    (PE148_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE149 (
    .activate  (PE148_acount[7:0]               ), //i
    .weight    (PE049_bcount[7:0]               ), //i
    .valid     (PE149_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE149_acount[7:0]               ), //o
    .bcount    (PE149_bcount[7:0]               ), //o
    .PE_OUT    (PE149_PE_OUT[31:0]              ), //o
    .finish    (PE149_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE150 (
    .activate  (PE149_acount[7:0]               ), //i
    .weight    (PE050_bcount[7:0]               ), //i
    .valid     (PE150_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE150_acount[7:0]               ), //o
    .bcount    (PE150_bcount[7:0]               ), //o
    .PE_OUT    (PE150_PE_OUT[31:0]              ), //o
    .finish    (PE150_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE151 (
    .activate  (PE150_acount[7:0]               ), //i
    .weight    (PE051_bcount[7:0]               ), //i
    .valid     (PE151_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE151_acount[7:0]               ), //o
    .bcount    (PE151_bcount[7:0]               ), //o
    .PE_OUT    (PE151_PE_OUT[31:0]              ), //o
    .finish    (PE151_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE152 (
    .activate  (PE151_acount[7:0]               ), //i
    .weight    (PE052_bcount[7:0]               ), //i
    .valid     (PE152_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE152_acount[7:0]               ), //o
    .bcount    (PE152_bcount[7:0]               ), //o
    .PE_OUT    (PE152_PE_OUT[31:0]              ), //o
    .finish    (PE152_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE153 (
    .activate  (PE152_acount[7:0]               ), //i
    .weight    (PE053_bcount[7:0]               ), //i
    .valid     (PE153_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE153_acount[7:0]               ), //o
    .bcount    (PE153_bcount[7:0]               ), //o
    .PE_OUT    (PE153_PE_OUT[31:0]              ), //o
    .finish    (PE153_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE154 (
    .activate  (PE153_acount[7:0]               ), //i
    .weight    (PE054_bcount[7:0]               ), //i
    .valid     (PE154_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE154_acount[7:0]               ), //o
    .bcount    (PE154_bcount[7:0]               ), //o
    .PE_OUT    (PE154_PE_OUT[31:0]              ), //o
    .finish    (PE154_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE155 (
    .activate  (PE154_acount[7:0]               ), //i
    .weight    (PE055_bcount[7:0]               ), //i
    .valid     (PE155_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE155_acount[7:0]               ), //o
    .bcount    (PE155_bcount[7:0]               ), //o
    .PE_OUT    (PE155_PE_OUT[31:0]              ), //o
    .finish    (PE155_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE156 (
    .activate  (PE155_acount[7:0]               ), //i
    .weight    (PE056_bcount[7:0]               ), //i
    .valid     (PE156_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE156_acount[7:0]               ), //o
    .bcount    (PE156_bcount[7:0]               ), //o
    .PE_OUT    (PE156_PE_OUT[31:0]              ), //o
    .finish    (PE156_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE157 (
    .activate  (PE156_acount[7:0]               ), //i
    .weight    (PE057_bcount[7:0]               ), //i
    .valid     (PE157_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE157_acount[7:0]               ), //o
    .bcount    (PE157_bcount[7:0]               ), //o
    .PE_OUT    (PE157_PE_OUT[31:0]              ), //o
    .finish    (PE157_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE158 (
    .activate  (PE157_acount[7:0]               ), //i
    .weight    (PE058_bcount[7:0]               ), //i
    .valid     (PE158_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE158_acount[7:0]               ), //o
    .bcount    (PE158_bcount[7:0]               ), //o
    .PE_OUT    (PE158_PE_OUT[31:0]              ), //o
    .finish    (PE158_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE159 (
    .activate  (PE158_acount[7:0]               ), //i
    .weight    (PE059_bcount[7:0]               ), //i
    .valid     (PE159_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE159_acount[7:0]               ), //o
    .bcount    (PE159_bcount[7:0]               ), //o
    .PE_OUT    (PE159_PE_OUT[31:0]              ), //o
    .finish    (PE159_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE160 (
    .activate  (PE159_acount[7:0]               ), //i
    .weight    (PE060_bcount[7:0]               ), //i
    .valid     (PE160_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE160_acount[7:0]               ), //o
    .bcount    (PE160_bcount[7:0]               ), //o
    .PE_OUT    (PE160_PE_OUT[31:0]              ), //o
    .finish    (PE160_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE161 (
    .activate  (PE160_acount[7:0]               ), //i
    .weight    (PE061_bcount[7:0]               ), //i
    .valid     (PE161_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE161_acount[7:0]               ), //o
    .bcount    (PE161_bcount[7:0]               ), //o
    .PE_OUT    (PE161_PE_OUT[31:0]              ), //o
    .finish    (PE161_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE162 (
    .activate  (PE161_acount[7:0]               ), //i
    .weight    (PE062_bcount[7:0]               ), //i
    .valid     (PE162_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE162_acount[7:0]               ), //o
    .bcount    (PE162_bcount[7:0]               ), //o
    .PE_OUT    (PE162_PE_OUT[31:0]              ), //o
    .finish    (PE162_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE163 (
    .activate  (PE162_acount[7:0]               ), //i
    .weight    (PE063_bcount[7:0]               ), //i
    .valid     (PE163_valid                     ), //i
    .signCount (io_signCount_regNextWhen_1[15:0]), //i
    .acount    (PE163_acount[7:0]               ), //o
    .bcount    (PE163_bcount[7:0]               ), //o
    .PE_OUT    (PE163_PE_OUT[31:0]              ), //o
    .finish    (PE163_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE20 (
    .activate  (io_MatrixA_2[7:0]               ), //i
    .weight    (PE10_bcount[7:0]                ), //i
    .valid     (PE20_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE20_acount[7:0]                ), //o
    .bcount    (PE20_bcount[7:0]                ), //o
    .PE_OUT    (PE20_PE_OUT[31:0]               ), //o
    .finish    (PE20_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE21 (
    .activate  (PE20_acount[7:0]                ), //i
    .weight    (PE11_bcount[7:0]                ), //i
    .valid     (PE21_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE21_acount[7:0]                ), //o
    .bcount    (PE21_bcount[7:0]                ), //o
    .PE_OUT    (PE21_PE_OUT[31:0]               ), //o
    .finish    (PE21_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE22 (
    .activate  (PE21_acount[7:0]                ), //i
    .weight    (PE12_bcount[7:0]                ), //i
    .valid     (PE22_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE22_acount[7:0]                ), //o
    .bcount    (PE22_bcount[7:0]                ), //o
    .PE_OUT    (PE22_PE_OUT[31:0]               ), //o
    .finish    (PE22_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE23 (
    .activate  (PE22_acount[7:0]                ), //i
    .weight    (PE13_bcount[7:0]                ), //i
    .valid     (PE23_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE23_acount[7:0]                ), //o
    .bcount    (PE23_bcount[7:0]                ), //o
    .PE_OUT    (PE23_PE_OUT[31:0]               ), //o
    .finish    (PE23_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE24 (
    .activate  (PE23_acount[7:0]                ), //i
    .weight    (PE14_bcount[7:0]                ), //i
    .valid     (PE24_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE24_acount[7:0]                ), //o
    .bcount    (PE24_bcount[7:0]                ), //o
    .PE_OUT    (PE24_PE_OUT[31:0]               ), //o
    .finish    (PE24_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE25 (
    .activate  (PE24_acount[7:0]                ), //i
    .weight    (PE15_bcount[7:0]                ), //i
    .valid     (PE25_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE25_acount[7:0]                ), //o
    .bcount    (PE25_bcount[7:0]                ), //o
    .PE_OUT    (PE25_PE_OUT[31:0]               ), //o
    .finish    (PE25_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE26 (
    .activate  (PE25_acount[7:0]                ), //i
    .weight    (PE16_bcount[7:0]                ), //i
    .valid     (PE26_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE26_acount[7:0]                ), //o
    .bcount    (PE26_bcount[7:0]                ), //o
    .PE_OUT    (PE26_PE_OUT[31:0]               ), //o
    .finish    (PE26_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE27 (
    .activate  (PE26_acount[7:0]                ), //i
    .weight    (PE17_bcount[7:0]                ), //i
    .valid     (PE27_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE27_acount[7:0]                ), //o
    .bcount    (PE27_bcount[7:0]                ), //o
    .PE_OUT    (PE27_PE_OUT[31:0]               ), //o
    .finish    (PE27_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE28 (
    .activate  (PE27_acount[7:0]                ), //i
    .weight    (PE18_bcount[7:0]                ), //i
    .valid     (PE28_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE28_acount[7:0]                ), //o
    .bcount    (PE28_bcount[7:0]                ), //o
    .PE_OUT    (PE28_PE_OUT[31:0]               ), //o
    .finish    (PE28_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE29 (
    .activate  (PE28_acount[7:0]                ), //i
    .weight    (PE19_bcount[7:0]                ), //i
    .valid     (PE29_valid                      ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE29_acount[7:0]                ), //o
    .bcount    (PE29_bcount[7:0]                ), //o
    .PE_OUT    (PE29_PE_OUT[31:0]               ), //o
    .finish    (PE29_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE210 (
    .activate  (PE29_acount[7:0]                ), //i
    .weight    (PE110_bcount[7:0]               ), //i
    .valid     (PE210_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE210_acount[7:0]               ), //o
    .bcount    (PE210_bcount[7:0]               ), //o
    .PE_OUT    (PE210_PE_OUT[31:0]              ), //o
    .finish    (PE210_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE211 (
    .activate  (PE210_acount[7:0]               ), //i
    .weight    (PE111_bcount[7:0]               ), //i
    .valid     (PE211_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE211_acount[7:0]               ), //o
    .bcount    (PE211_bcount[7:0]               ), //o
    .PE_OUT    (PE211_PE_OUT[31:0]              ), //o
    .finish    (PE211_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE212 (
    .activate  (PE211_acount[7:0]               ), //i
    .weight    (PE112_bcount[7:0]               ), //i
    .valid     (PE212_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE212_acount[7:0]               ), //o
    .bcount    (PE212_bcount[7:0]               ), //o
    .PE_OUT    (PE212_PE_OUT[31:0]              ), //o
    .finish    (PE212_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE213 (
    .activate  (PE212_acount[7:0]               ), //i
    .weight    (PE113_bcount[7:0]               ), //i
    .valid     (PE213_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE213_acount[7:0]               ), //o
    .bcount    (PE213_bcount[7:0]               ), //o
    .PE_OUT    (PE213_PE_OUT[31:0]              ), //o
    .finish    (PE213_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE214 (
    .activate  (PE213_acount[7:0]               ), //i
    .weight    (PE114_bcount[7:0]               ), //i
    .valid     (PE214_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE214_acount[7:0]               ), //o
    .bcount    (PE214_bcount[7:0]               ), //o
    .PE_OUT    (PE214_PE_OUT[31:0]              ), //o
    .finish    (PE214_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE215 (
    .activate  (PE214_acount[7:0]               ), //i
    .weight    (PE115_bcount[7:0]               ), //i
    .valid     (PE215_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE215_acount[7:0]               ), //o
    .bcount    (PE215_bcount[7:0]               ), //o
    .PE_OUT    (PE215_PE_OUT[31:0]              ), //o
    .finish    (PE215_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE216 (
    .activate  (PE215_acount[7:0]               ), //i
    .weight    (PE116_bcount[7:0]               ), //i
    .valid     (PE216_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE216_acount[7:0]               ), //o
    .bcount    (PE216_bcount[7:0]               ), //o
    .PE_OUT    (PE216_PE_OUT[31:0]              ), //o
    .finish    (PE216_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE217 (
    .activate  (PE216_acount[7:0]               ), //i
    .weight    (PE117_bcount[7:0]               ), //i
    .valid     (PE217_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE217_acount[7:0]               ), //o
    .bcount    (PE217_bcount[7:0]               ), //o
    .PE_OUT    (PE217_PE_OUT[31:0]              ), //o
    .finish    (PE217_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE218 (
    .activate  (PE217_acount[7:0]               ), //i
    .weight    (PE118_bcount[7:0]               ), //i
    .valid     (PE218_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE218_acount[7:0]               ), //o
    .bcount    (PE218_bcount[7:0]               ), //o
    .PE_OUT    (PE218_PE_OUT[31:0]              ), //o
    .finish    (PE218_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE219 (
    .activate  (PE218_acount[7:0]               ), //i
    .weight    (PE119_bcount[7:0]               ), //i
    .valid     (PE219_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE219_acount[7:0]               ), //o
    .bcount    (PE219_bcount[7:0]               ), //o
    .PE_OUT    (PE219_PE_OUT[31:0]              ), //o
    .finish    (PE219_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE220 (
    .activate  (PE219_acount[7:0]               ), //i
    .weight    (PE120_bcount[7:0]               ), //i
    .valid     (PE220_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE220_acount[7:0]               ), //o
    .bcount    (PE220_bcount[7:0]               ), //o
    .PE_OUT    (PE220_PE_OUT[31:0]              ), //o
    .finish    (PE220_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE221 (
    .activate  (PE220_acount[7:0]               ), //i
    .weight    (PE121_bcount[7:0]               ), //i
    .valid     (PE221_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE221_acount[7:0]               ), //o
    .bcount    (PE221_bcount[7:0]               ), //o
    .PE_OUT    (PE221_PE_OUT[31:0]              ), //o
    .finish    (PE221_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE222 (
    .activate  (PE221_acount[7:0]               ), //i
    .weight    (PE122_bcount[7:0]               ), //i
    .valid     (PE222_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE222_acount[7:0]               ), //o
    .bcount    (PE222_bcount[7:0]               ), //o
    .PE_OUT    (PE222_PE_OUT[31:0]              ), //o
    .finish    (PE222_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE223 (
    .activate  (PE222_acount[7:0]               ), //i
    .weight    (PE123_bcount[7:0]               ), //i
    .valid     (PE223_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE223_acount[7:0]               ), //o
    .bcount    (PE223_bcount[7:0]               ), //o
    .PE_OUT    (PE223_PE_OUT[31:0]              ), //o
    .finish    (PE223_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE224 (
    .activate  (PE223_acount[7:0]               ), //i
    .weight    (PE124_bcount[7:0]               ), //i
    .valid     (PE224_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE224_acount[7:0]               ), //o
    .bcount    (PE224_bcount[7:0]               ), //o
    .PE_OUT    (PE224_PE_OUT[31:0]              ), //o
    .finish    (PE224_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE225 (
    .activate  (PE224_acount[7:0]               ), //i
    .weight    (PE125_bcount[7:0]               ), //i
    .valid     (PE225_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE225_acount[7:0]               ), //o
    .bcount    (PE225_bcount[7:0]               ), //o
    .PE_OUT    (PE225_PE_OUT[31:0]              ), //o
    .finish    (PE225_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE226 (
    .activate  (PE225_acount[7:0]               ), //i
    .weight    (PE126_bcount[7:0]               ), //i
    .valid     (PE226_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE226_acount[7:0]               ), //o
    .bcount    (PE226_bcount[7:0]               ), //o
    .PE_OUT    (PE226_PE_OUT[31:0]              ), //o
    .finish    (PE226_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE227 (
    .activate  (PE226_acount[7:0]               ), //i
    .weight    (PE127_bcount[7:0]               ), //i
    .valid     (PE227_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE227_acount[7:0]               ), //o
    .bcount    (PE227_bcount[7:0]               ), //o
    .PE_OUT    (PE227_PE_OUT[31:0]              ), //o
    .finish    (PE227_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE228 (
    .activate  (PE227_acount[7:0]               ), //i
    .weight    (PE128_bcount[7:0]               ), //i
    .valid     (PE228_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE228_acount[7:0]               ), //o
    .bcount    (PE228_bcount[7:0]               ), //o
    .PE_OUT    (PE228_PE_OUT[31:0]              ), //o
    .finish    (PE228_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE229 (
    .activate  (PE228_acount[7:0]               ), //i
    .weight    (PE129_bcount[7:0]               ), //i
    .valid     (PE229_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE229_acount[7:0]               ), //o
    .bcount    (PE229_bcount[7:0]               ), //o
    .PE_OUT    (PE229_PE_OUT[31:0]              ), //o
    .finish    (PE229_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE230 (
    .activate  (PE229_acount[7:0]               ), //i
    .weight    (PE130_bcount[7:0]               ), //i
    .valid     (PE230_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE230_acount[7:0]               ), //o
    .bcount    (PE230_bcount[7:0]               ), //o
    .PE_OUT    (PE230_PE_OUT[31:0]              ), //o
    .finish    (PE230_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE231 (
    .activate  (PE230_acount[7:0]               ), //i
    .weight    (PE131_bcount[7:0]               ), //i
    .valid     (PE231_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE231_acount[7:0]               ), //o
    .bcount    (PE231_bcount[7:0]               ), //o
    .PE_OUT    (PE231_PE_OUT[31:0]              ), //o
    .finish    (PE231_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE232 (
    .activate  (PE231_acount[7:0]               ), //i
    .weight    (PE132_bcount[7:0]               ), //i
    .valid     (PE232_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE232_acount[7:0]               ), //o
    .bcount    (PE232_bcount[7:0]               ), //o
    .PE_OUT    (PE232_PE_OUT[31:0]              ), //o
    .finish    (PE232_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE233 (
    .activate  (PE232_acount[7:0]               ), //i
    .weight    (PE133_bcount[7:0]               ), //i
    .valid     (PE233_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE233_acount[7:0]               ), //o
    .bcount    (PE233_bcount[7:0]               ), //o
    .PE_OUT    (PE233_PE_OUT[31:0]              ), //o
    .finish    (PE233_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE234 (
    .activate  (PE233_acount[7:0]               ), //i
    .weight    (PE134_bcount[7:0]               ), //i
    .valid     (PE234_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE234_acount[7:0]               ), //o
    .bcount    (PE234_bcount[7:0]               ), //o
    .PE_OUT    (PE234_PE_OUT[31:0]              ), //o
    .finish    (PE234_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE235 (
    .activate  (PE234_acount[7:0]               ), //i
    .weight    (PE135_bcount[7:0]               ), //i
    .valid     (PE235_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE235_acount[7:0]               ), //o
    .bcount    (PE235_bcount[7:0]               ), //o
    .PE_OUT    (PE235_PE_OUT[31:0]              ), //o
    .finish    (PE235_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE236 (
    .activate  (PE235_acount[7:0]               ), //i
    .weight    (PE136_bcount[7:0]               ), //i
    .valid     (PE236_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE236_acount[7:0]               ), //o
    .bcount    (PE236_bcount[7:0]               ), //o
    .PE_OUT    (PE236_PE_OUT[31:0]              ), //o
    .finish    (PE236_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE237 (
    .activate  (PE236_acount[7:0]               ), //i
    .weight    (PE137_bcount[7:0]               ), //i
    .valid     (PE237_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE237_acount[7:0]               ), //o
    .bcount    (PE237_bcount[7:0]               ), //o
    .PE_OUT    (PE237_PE_OUT[31:0]              ), //o
    .finish    (PE237_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE238 (
    .activate  (PE237_acount[7:0]               ), //i
    .weight    (PE138_bcount[7:0]               ), //i
    .valid     (PE238_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE238_acount[7:0]               ), //o
    .bcount    (PE238_bcount[7:0]               ), //o
    .PE_OUT    (PE238_PE_OUT[31:0]              ), //o
    .finish    (PE238_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE239 (
    .activate  (PE238_acount[7:0]               ), //i
    .weight    (PE139_bcount[7:0]               ), //i
    .valid     (PE239_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE239_acount[7:0]               ), //o
    .bcount    (PE239_bcount[7:0]               ), //o
    .PE_OUT    (PE239_PE_OUT[31:0]              ), //o
    .finish    (PE239_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE240 (
    .activate  (PE239_acount[7:0]               ), //i
    .weight    (PE140_bcount[7:0]               ), //i
    .valid     (PE240_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE240_acount[7:0]               ), //o
    .bcount    (PE240_bcount[7:0]               ), //o
    .PE_OUT    (PE240_PE_OUT[31:0]              ), //o
    .finish    (PE240_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE241 (
    .activate  (PE240_acount[7:0]               ), //i
    .weight    (PE141_bcount[7:0]               ), //i
    .valid     (PE241_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE241_acount[7:0]               ), //o
    .bcount    (PE241_bcount[7:0]               ), //o
    .PE_OUT    (PE241_PE_OUT[31:0]              ), //o
    .finish    (PE241_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE242 (
    .activate  (PE241_acount[7:0]               ), //i
    .weight    (PE142_bcount[7:0]               ), //i
    .valid     (PE242_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE242_acount[7:0]               ), //o
    .bcount    (PE242_bcount[7:0]               ), //o
    .PE_OUT    (PE242_PE_OUT[31:0]              ), //o
    .finish    (PE242_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE243 (
    .activate  (PE242_acount[7:0]               ), //i
    .weight    (PE143_bcount[7:0]               ), //i
    .valid     (PE243_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE243_acount[7:0]               ), //o
    .bcount    (PE243_bcount[7:0]               ), //o
    .PE_OUT    (PE243_PE_OUT[31:0]              ), //o
    .finish    (PE243_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE244 (
    .activate  (PE243_acount[7:0]               ), //i
    .weight    (PE144_bcount[7:0]               ), //i
    .valid     (PE244_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE244_acount[7:0]               ), //o
    .bcount    (PE244_bcount[7:0]               ), //o
    .PE_OUT    (PE244_PE_OUT[31:0]              ), //o
    .finish    (PE244_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE245 (
    .activate  (PE244_acount[7:0]               ), //i
    .weight    (PE145_bcount[7:0]               ), //i
    .valid     (PE245_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE245_acount[7:0]               ), //o
    .bcount    (PE245_bcount[7:0]               ), //o
    .PE_OUT    (PE245_PE_OUT[31:0]              ), //o
    .finish    (PE245_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE246 (
    .activate  (PE245_acount[7:0]               ), //i
    .weight    (PE146_bcount[7:0]               ), //i
    .valid     (PE246_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE246_acount[7:0]               ), //o
    .bcount    (PE246_bcount[7:0]               ), //o
    .PE_OUT    (PE246_PE_OUT[31:0]              ), //o
    .finish    (PE246_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE247 (
    .activate  (PE246_acount[7:0]               ), //i
    .weight    (PE147_bcount[7:0]               ), //i
    .valid     (PE247_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE247_acount[7:0]               ), //o
    .bcount    (PE247_bcount[7:0]               ), //o
    .PE_OUT    (PE247_PE_OUT[31:0]              ), //o
    .finish    (PE247_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE248 (
    .activate  (PE247_acount[7:0]               ), //i
    .weight    (PE148_bcount[7:0]               ), //i
    .valid     (PE248_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE248_acount[7:0]               ), //o
    .bcount    (PE248_bcount[7:0]               ), //o
    .PE_OUT    (PE248_PE_OUT[31:0]              ), //o
    .finish    (PE248_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE249 (
    .activate  (PE248_acount[7:0]               ), //i
    .weight    (PE149_bcount[7:0]               ), //i
    .valid     (PE249_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE249_acount[7:0]               ), //o
    .bcount    (PE249_bcount[7:0]               ), //o
    .PE_OUT    (PE249_PE_OUT[31:0]              ), //o
    .finish    (PE249_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE250 (
    .activate  (PE249_acount[7:0]               ), //i
    .weight    (PE150_bcount[7:0]               ), //i
    .valid     (PE250_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE250_acount[7:0]               ), //o
    .bcount    (PE250_bcount[7:0]               ), //o
    .PE_OUT    (PE250_PE_OUT[31:0]              ), //o
    .finish    (PE250_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE251 (
    .activate  (PE250_acount[7:0]               ), //i
    .weight    (PE151_bcount[7:0]               ), //i
    .valid     (PE251_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE251_acount[7:0]               ), //o
    .bcount    (PE251_bcount[7:0]               ), //o
    .PE_OUT    (PE251_PE_OUT[31:0]              ), //o
    .finish    (PE251_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE252 (
    .activate  (PE251_acount[7:0]               ), //i
    .weight    (PE152_bcount[7:0]               ), //i
    .valid     (PE252_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE252_acount[7:0]               ), //o
    .bcount    (PE252_bcount[7:0]               ), //o
    .PE_OUT    (PE252_PE_OUT[31:0]              ), //o
    .finish    (PE252_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE253 (
    .activate  (PE252_acount[7:0]               ), //i
    .weight    (PE153_bcount[7:0]               ), //i
    .valid     (PE253_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE253_acount[7:0]               ), //o
    .bcount    (PE253_bcount[7:0]               ), //o
    .PE_OUT    (PE253_PE_OUT[31:0]              ), //o
    .finish    (PE253_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE254 (
    .activate  (PE253_acount[7:0]               ), //i
    .weight    (PE154_bcount[7:0]               ), //i
    .valid     (PE254_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE254_acount[7:0]               ), //o
    .bcount    (PE254_bcount[7:0]               ), //o
    .PE_OUT    (PE254_PE_OUT[31:0]              ), //o
    .finish    (PE254_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE255 (
    .activate  (PE254_acount[7:0]               ), //i
    .weight    (PE155_bcount[7:0]               ), //i
    .valid     (PE255_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE255_acount[7:0]               ), //o
    .bcount    (PE255_bcount[7:0]               ), //o
    .PE_OUT    (PE255_PE_OUT[31:0]              ), //o
    .finish    (PE255_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE256 (
    .activate  (PE255_acount[7:0]               ), //i
    .weight    (PE156_bcount[7:0]               ), //i
    .valid     (PE256_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE256_acount[7:0]               ), //o
    .bcount    (PE256_bcount[7:0]               ), //o
    .PE_OUT    (PE256_PE_OUT[31:0]              ), //o
    .finish    (PE256_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE257 (
    .activate  (PE256_acount[7:0]               ), //i
    .weight    (PE157_bcount[7:0]               ), //i
    .valid     (PE257_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE257_acount[7:0]               ), //o
    .bcount    (PE257_bcount[7:0]               ), //o
    .PE_OUT    (PE257_PE_OUT[31:0]              ), //o
    .finish    (PE257_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE258 (
    .activate  (PE257_acount[7:0]               ), //i
    .weight    (PE158_bcount[7:0]               ), //i
    .valid     (PE258_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE258_acount[7:0]               ), //o
    .bcount    (PE258_bcount[7:0]               ), //o
    .PE_OUT    (PE258_PE_OUT[31:0]              ), //o
    .finish    (PE258_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE259 (
    .activate  (PE258_acount[7:0]               ), //i
    .weight    (PE159_bcount[7:0]               ), //i
    .valid     (PE259_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE259_acount[7:0]               ), //o
    .bcount    (PE259_bcount[7:0]               ), //o
    .PE_OUT    (PE259_PE_OUT[31:0]              ), //o
    .finish    (PE259_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE260 (
    .activate  (PE259_acount[7:0]               ), //i
    .weight    (PE160_bcount[7:0]               ), //i
    .valid     (PE260_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE260_acount[7:0]               ), //o
    .bcount    (PE260_bcount[7:0]               ), //o
    .PE_OUT    (PE260_PE_OUT[31:0]              ), //o
    .finish    (PE260_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE261 (
    .activate  (PE260_acount[7:0]               ), //i
    .weight    (PE161_bcount[7:0]               ), //i
    .valid     (PE261_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE261_acount[7:0]               ), //o
    .bcount    (PE261_bcount[7:0]               ), //o
    .PE_OUT    (PE261_PE_OUT[31:0]              ), //o
    .finish    (PE261_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE262 (
    .activate  (PE261_acount[7:0]               ), //i
    .weight    (PE162_bcount[7:0]               ), //i
    .valid     (PE262_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE262_acount[7:0]               ), //o
    .bcount    (PE262_bcount[7:0]               ), //o
    .PE_OUT    (PE262_PE_OUT[31:0]              ), //o
    .finish    (PE262_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE263 (
    .activate  (PE262_acount[7:0]               ), //i
    .weight    (PE163_bcount[7:0]               ), //i
    .valid     (PE263_valid                     ), //i
    .signCount (io_signCount_regNextWhen_2[15:0]), //i
    .acount    (PE263_acount[7:0]               ), //o
    .bcount    (PE263_bcount[7:0]               ), //o
    .PE_OUT    (PE263_PE_OUT[31:0]              ), //o
    .finish    (PE263_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE30 (
    .activate  (io_MatrixA_3[7:0]               ), //i
    .weight    (PE20_bcount[7:0]                ), //i
    .valid     (PE30_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE30_acount[7:0]                ), //o
    .bcount    (PE30_bcount[7:0]                ), //o
    .PE_OUT    (PE30_PE_OUT[31:0]               ), //o
    .finish    (PE30_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE31 (
    .activate  (PE30_acount[7:0]                ), //i
    .weight    (PE21_bcount[7:0]                ), //i
    .valid     (PE31_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE31_acount[7:0]                ), //o
    .bcount    (PE31_bcount[7:0]                ), //o
    .PE_OUT    (PE31_PE_OUT[31:0]               ), //o
    .finish    (PE31_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE32 (
    .activate  (PE31_acount[7:0]                ), //i
    .weight    (PE22_bcount[7:0]                ), //i
    .valid     (PE32_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE32_acount[7:0]                ), //o
    .bcount    (PE32_bcount[7:0]                ), //o
    .PE_OUT    (PE32_PE_OUT[31:0]               ), //o
    .finish    (PE32_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE33 (
    .activate  (PE32_acount[7:0]                ), //i
    .weight    (PE23_bcount[7:0]                ), //i
    .valid     (PE33_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE33_acount[7:0]                ), //o
    .bcount    (PE33_bcount[7:0]                ), //o
    .PE_OUT    (PE33_PE_OUT[31:0]               ), //o
    .finish    (PE33_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE34 (
    .activate  (PE33_acount[7:0]                ), //i
    .weight    (PE24_bcount[7:0]                ), //i
    .valid     (PE34_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE34_acount[7:0]                ), //o
    .bcount    (PE34_bcount[7:0]                ), //o
    .PE_OUT    (PE34_PE_OUT[31:0]               ), //o
    .finish    (PE34_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE35 (
    .activate  (PE34_acount[7:0]                ), //i
    .weight    (PE25_bcount[7:0]                ), //i
    .valid     (PE35_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE35_acount[7:0]                ), //o
    .bcount    (PE35_bcount[7:0]                ), //o
    .PE_OUT    (PE35_PE_OUT[31:0]               ), //o
    .finish    (PE35_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE36 (
    .activate  (PE35_acount[7:0]                ), //i
    .weight    (PE26_bcount[7:0]                ), //i
    .valid     (PE36_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE36_acount[7:0]                ), //o
    .bcount    (PE36_bcount[7:0]                ), //o
    .PE_OUT    (PE36_PE_OUT[31:0]               ), //o
    .finish    (PE36_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE37 (
    .activate  (PE36_acount[7:0]                ), //i
    .weight    (PE27_bcount[7:0]                ), //i
    .valid     (PE37_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE37_acount[7:0]                ), //o
    .bcount    (PE37_bcount[7:0]                ), //o
    .PE_OUT    (PE37_PE_OUT[31:0]               ), //o
    .finish    (PE37_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE38 (
    .activate  (PE37_acount[7:0]                ), //i
    .weight    (PE28_bcount[7:0]                ), //i
    .valid     (PE38_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE38_acount[7:0]                ), //o
    .bcount    (PE38_bcount[7:0]                ), //o
    .PE_OUT    (PE38_PE_OUT[31:0]               ), //o
    .finish    (PE38_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE39 (
    .activate  (PE38_acount[7:0]                ), //i
    .weight    (PE29_bcount[7:0]                ), //i
    .valid     (PE39_valid                      ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE39_acount[7:0]                ), //o
    .bcount    (PE39_bcount[7:0]                ), //o
    .PE_OUT    (PE39_PE_OUT[31:0]               ), //o
    .finish    (PE39_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE310 (
    .activate  (PE39_acount[7:0]                ), //i
    .weight    (PE210_bcount[7:0]               ), //i
    .valid     (PE310_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE310_acount[7:0]               ), //o
    .bcount    (PE310_bcount[7:0]               ), //o
    .PE_OUT    (PE310_PE_OUT[31:0]              ), //o
    .finish    (PE310_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE311 (
    .activate  (PE310_acount[7:0]               ), //i
    .weight    (PE211_bcount[7:0]               ), //i
    .valid     (PE311_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE311_acount[7:0]               ), //o
    .bcount    (PE311_bcount[7:0]               ), //o
    .PE_OUT    (PE311_PE_OUT[31:0]              ), //o
    .finish    (PE311_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE312 (
    .activate  (PE311_acount[7:0]               ), //i
    .weight    (PE212_bcount[7:0]               ), //i
    .valid     (PE312_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE312_acount[7:0]               ), //o
    .bcount    (PE312_bcount[7:0]               ), //o
    .PE_OUT    (PE312_PE_OUT[31:0]              ), //o
    .finish    (PE312_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE313 (
    .activate  (PE312_acount[7:0]               ), //i
    .weight    (PE213_bcount[7:0]               ), //i
    .valid     (PE313_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE313_acount[7:0]               ), //o
    .bcount    (PE313_bcount[7:0]               ), //o
    .PE_OUT    (PE313_PE_OUT[31:0]              ), //o
    .finish    (PE313_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE314 (
    .activate  (PE313_acount[7:0]               ), //i
    .weight    (PE214_bcount[7:0]               ), //i
    .valid     (PE314_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE314_acount[7:0]               ), //o
    .bcount    (PE314_bcount[7:0]               ), //o
    .PE_OUT    (PE314_PE_OUT[31:0]              ), //o
    .finish    (PE314_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE315 (
    .activate  (PE314_acount[7:0]               ), //i
    .weight    (PE215_bcount[7:0]               ), //i
    .valid     (PE315_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE315_acount[7:0]               ), //o
    .bcount    (PE315_bcount[7:0]               ), //o
    .PE_OUT    (PE315_PE_OUT[31:0]              ), //o
    .finish    (PE315_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE316 (
    .activate  (PE315_acount[7:0]               ), //i
    .weight    (PE216_bcount[7:0]               ), //i
    .valid     (PE316_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE316_acount[7:0]               ), //o
    .bcount    (PE316_bcount[7:0]               ), //o
    .PE_OUT    (PE316_PE_OUT[31:0]              ), //o
    .finish    (PE316_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE317 (
    .activate  (PE316_acount[7:0]               ), //i
    .weight    (PE217_bcount[7:0]               ), //i
    .valid     (PE317_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE317_acount[7:0]               ), //o
    .bcount    (PE317_bcount[7:0]               ), //o
    .PE_OUT    (PE317_PE_OUT[31:0]              ), //o
    .finish    (PE317_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE318 (
    .activate  (PE317_acount[7:0]               ), //i
    .weight    (PE218_bcount[7:0]               ), //i
    .valid     (PE318_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE318_acount[7:0]               ), //o
    .bcount    (PE318_bcount[7:0]               ), //o
    .PE_OUT    (PE318_PE_OUT[31:0]              ), //o
    .finish    (PE318_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE319 (
    .activate  (PE318_acount[7:0]               ), //i
    .weight    (PE219_bcount[7:0]               ), //i
    .valid     (PE319_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE319_acount[7:0]               ), //o
    .bcount    (PE319_bcount[7:0]               ), //o
    .PE_OUT    (PE319_PE_OUT[31:0]              ), //o
    .finish    (PE319_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE320 (
    .activate  (PE319_acount[7:0]               ), //i
    .weight    (PE220_bcount[7:0]               ), //i
    .valid     (PE320_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE320_acount[7:0]               ), //o
    .bcount    (PE320_bcount[7:0]               ), //o
    .PE_OUT    (PE320_PE_OUT[31:0]              ), //o
    .finish    (PE320_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE321 (
    .activate  (PE320_acount[7:0]               ), //i
    .weight    (PE221_bcount[7:0]               ), //i
    .valid     (PE321_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE321_acount[7:0]               ), //o
    .bcount    (PE321_bcount[7:0]               ), //o
    .PE_OUT    (PE321_PE_OUT[31:0]              ), //o
    .finish    (PE321_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE322 (
    .activate  (PE321_acount[7:0]               ), //i
    .weight    (PE222_bcount[7:0]               ), //i
    .valid     (PE322_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE322_acount[7:0]               ), //o
    .bcount    (PE322_bcount[7:0]               ), //o
    .PE_OUT    (PE322_PE_OUT[31:0]              ), //o
    .finish    (PE322_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE323 (
    .activate  (PE322_acount[7:0]               ), //i
    .weight    (PE223_bcount[7:0]               ), //i
    .valid     (PE323_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE323_acount[7:0]               ), //o
    .bcount    (PE323_bcount[7:0]               ), //o
    .PE_OUT    (PE323_PE_OUT[31:0]              ), //o
    .finish    (PE323_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE324 (
    .activate  (PE323_acount[7:0]               ), //i
    .weight    (PE224_bcount[7:0]               ), //i
    .valid     (PE324_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE324_acount[7:0]               ), //o
    .bcount    (PE324_bcount[7:0]               ), //o
    .PE_OUT    (PE324_PE_OUT[31:0]              ), //o
    .finish    (PE324_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE325 (
    .activate  (PE324_acount[7:0]               ), //i
    .weight    (PE225_bcount[7:0]               ), //i
    .valid     (PE325_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE325_acount[7:0]               ), //o
    .bcount    (PE325_bcount[7:0]               ), //o
    .PE_OUT    (PE325_PE_OUT[31:0]              ), //o
    .finish    (PE325_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE326 (
    .activate  (PE325_acount[7:0]               ), //i
    .weight    (PE226_bcount[7:0]               ), //i
    .valid     (PE326_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE326_acount[7:0]               ), //o
    .bcount    (PE326_bcount[7:0]               ), //o
    .PE_OUT    (PE326_PE_OUT[31:0]              ), //o
    .finish    (PE326_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE327 (
    .activate  (PE326_acount[7:0]               ), //i
    .weight    (PE227_bcount[7:0]               ), //i
    .valid     (PE327_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE327_acount[7:0]               ), //o
    .bcount    (PE327_bcount[7:0]               ), //o
    .PE_OUT    (PE327_PE_OUT[31:0]              ), //o
    .finish    (PE327_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE328 (
    .activate  (PE327_acount[7:0]               ), //i
    .weight    (PE228_bcount[7:0]               ), //i
    .valid     (PE328_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE328_acount[7:0]               ), //o
    .bcount    (PE328_bcount[7:0]               ), //o
    .PE_OUT    (PE328_PE_OUT[31:0]              ), //o
    .finish    (PE328_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE329 (
    .activate  (PE328_acount[7:0]               ), //i
    .weight    (PE229_bcount[7:0]               ), //i
    .valid     (PE329_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE329_acount[7:0]               ), //o
    .bcount    (PE329_bcount[7:0]               ), //o
    .PE_OUT    (PE329_PE_OUT[31:0]              ), //o
    .finish    (PE329_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE330 (
    .activate  (PE329_acount[7:0]               ), //i
    .weight    (PE230_bcount[7:0]               ), //i
    .valid     (PE330_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE330_acount[7:0]               ), //o
    .bcount    (PE330_bcount[7:0]               ), //o
    .PE_OUT    (PE330_PE_OUT[31:0]              ), //o
    .finish    (PE330_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE331 (
    .activate  (PE330_acount[7:0]               ), //i
    .weight    (PE231_bcount[7:0]               ), //i
    .valid     (PE331_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE331_acount[7:0]               ), //o
    .bcount    (PE331_bcount[7:0]               ), //o
    .PE_OUT    (PE331_PE_OUT[31:0]              ), //o
    .finish    (PE331_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE332 (
    .activate  (PE331_acount[7:0]               ), //i
    .weight    (PE232_bcount[7:0]               ), //i
    .valid     (PE332_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE332_acount[7:0]               ), //o
    .bcount    (PE332_bcount[7:0]               ), //o
    .PE_OUT    (PE332_PE_OUT[31:0]              ), //o
    .finish    (PE332_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE333 (
    .activate  (PE332_acount[7:0]               ), //i
    .weight    (PE233_bcount[7:0]               ), //i
    .valid     (PE333_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE333_acount[7:0]               ), //o
    .bcount    (PE333_bcount[7:0]               ), //o
    .PE_OUT    (PE333_PE_OUT[31:0]              ), //o
    .finish    (PE333_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE334 (
    .activate  (PE333_acount[7:0]               ), //i
    .weight    (PE234_bcount[7:0]               ), //i
    .valid     (PE334_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE334_acount[7:0]               ), //o
    .bcount    (PE334_bcount[7:0]               ), //o
    .PE_OUT    (PE334_PE_OUT[31:0]              ), //o
    .finish    (PE334_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE335 (
    .activate  (PE334_acount[7:0]               ), //i
    .weight    (PE235_bcount[7:0]               ), //i
    .valid     (PE335_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE335_acount[7:0]               ), //o
    .bcount    (PE335_bcount[7:0]               ), //o
    .PE_OUT    (PE335_PE_OUT[31:0]              ), //o
    .finish    (PE335_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE336 (
    .activate  (PE335_acount[7:0]               ), //i
    .weight    (PE236_bcount[7:0]               ), //i
    .valid     (PE336_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE336_acount[7:0]               ), //o
    .bcount    (PE336_bcount[7:0]               ), //o
    .PE_OUT    (PE336_PE_OUT[31:0]              ), //o
    .finish    (PE336_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE337 (
    .activate  (PE336_acount[7:0]               ), //i
    .weight    (PE237_bcount[7:0]               ), //i
    .valid     (PE337_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE337_acount[7:0]               ), //o
    .bcount    (PE337_bcount[7:0]               ), //o
    .PE_OUT    (PE337_PE_OUT[31:0]              ), //o
    .finish    (PE337_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE338 (
    .activate  (PE337_acount[7:0]               ), //i
    .weight    (PE238_bcount[7:0]               ), //i
    .valid     (PE338_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE338_acount[7:0]               ), //o
    .bcount    (PE338_bcount[7:0]               ), //o
    .PE_OUT    (PE338_PE_OUT[31:0]              ), //o
    .finish    (PE338_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE339 (
    .activate  (PE338_acount[7:0]               ), //i
    .weight    (PE239_bcount[7:0]               ), //i
    .valid     (PE339_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE339_acount[7:0]               ), //o
    .bcount    (PE339_bcount[7:0]               ), //o
    .PE_OUT    (PE339_PE_OUT[31:0]              ), //o
    .finish    (PE339_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE340 (
    .activate  (PE339_acount[7:0]               ), //i
    .weight    (PE240_bcount[7:0]               ), //i
    .valid     (PE340_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE340_acount[7:0]               ), //o
    .bcount    (PE340_bcount[7:0]               ), //o
    .PE_OUT    (PE340_PE_OUT[31:0]              ), //o
    .finish    (PE340_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE341 (
    .activate  (PE340_acount[7:0]               ), //i
    .weight    (PE241_bcount[7:0]               ), //i
    .valid     (PE341_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE341_acount[7:0]               ), //o
    .bcount    (PE341_bcount[7:0]               ), //o
    .PE_OUT    (PE341_PE_OUT[31:0]              ), //o
    .finish    (PE341_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE342 (
    .activate  (PE341_acount[7:0]               ), //i
    .weight    (PE242_bcount[7:0]               ), //i
    .valid     (PE342_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE342_acount[7:0]               ), //o
    .bcount    (PE342_bcount[7:0]               ), //o
    .PE_OUT    (PE342_PE_OUT[31:0]              ), //o
    .finish    (PE342_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE343 (
    .activate  (PE342_acount[7:0]               ), //i
    .weight    (PE243_bcount[7:0]               ), //i
    .valid     (PE343_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE343_acount[7:0]               ), //o
    .bcount    (PE343_bcount[7:0]               ), //o
    .PE_OUT    (PE343_PE_OUT[31:0]              ), //o
    .finish    (PE343_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE344 (
    .activate  (PE343_acount[7:0]               ), //i
    .weight    (PE244_bcount[7:0]               ), //i
    .valid     (PE344_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE344_acount[7:0]               ), //o
    .bcount    (PE344_bcount[7:0]               ), //o
    .PE_OUT    (PE344_PE_OUT[31:0]              ), //o
    .finish    (PE344_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE345 (
    .activate  (PE344_acount[7:0]               ), //i
    .weight    (PE245_bcount[7:0]               ), //i
    .valid     (PE345_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE345_acount[7:0]               ), //o
    .bcount    (PE345_bcount[7:0]               ), //o
    .PE_OUT    (PE345_PE_OUT[31:0]              ), //o
    .finish    (PE345_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE346 (
    .activate  (PE345_acount[7:0]               ), //i
    .weight    (PE246_bcount[7:0]               ), //i
    .valid     (PE346_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE346_acount[7:0]               ), //o
    .bcount    (PE346_bcount[7:0]               ), //o
    .PE_OUT    (PE346_PE_OUT[31:0]              ), //o
    .finish    (PE346_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE347 (
    .activate  (PE346_acount[7:0]               ), //i
    .weight    (PE247_bcount[7:0]               ), //i
    .valid     (PE347_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE347_acount[7:0]               ), //o
    .bcount    (PE347_bcount[7:0]               ), //o
    .PE_OUT    (PE347_PE_OUT[31:0]              ), //o
    .finish    (PE347_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE348 (
    .activate  (PE347_acount[7:0]               ), //i
    .weight    (PE248_bcount[7:0]               ), //i
    .valid     (PE348_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE348_acount[7:0]               ), //o
    .bcount    (PE348_bcount[7:0]               ), //o
    .PE_OUT    (PE348_PE_OUT[31:0]              ), //o
    .finish    (PE348_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE349 (
    .activate  (PE348_acount[7:0]               ), //i
    .weight    (PE249_bcount[7:0]               ), //i
    .valid     (PE349_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE349_acount[7:0]               ), //o
    .bcount    (PE349_bcount[7:0]               ), //o
    .PE_OUT    (PE349_PE_OUT[31:0]              ), //o
    .finish    (PE349_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE350 (
    .activate  (PE349_acount[7:0]               ), //i
    .weight    (PE250_bcount[7:0]               ), //i
    .valid     (PE350_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE350_acount[7:0]               ), //o
    .bcount    (PE350_bcount[7:0]               ), //o
    .PE_OUT    (PE350_PE_OUT[31:0]              ), //o
    .finish    (PE350_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE351 (
    .activate  (PE350_acount[7:0]               ), //i
    .weight    (PE251_bcount[7:0]               ), //i
    .valid     (PE351_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE351_acount[7:0]               ), //o
    .bcount    (PE351_bcount[7:0]               ), //o
    .PE_OUT    (PE351_PE_OUT[31:0]              ), //o
    .finish    (PE351_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE352 (
    .activate  (PE351_acount[7:0]               ), //i
    .weight    (PE252_bcount[7:0]               ), //i
    .valid     (PE352_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE352_acount[7:0]               ), //o
    .bcount    (PE352_bcount[7:0]               ), //o
    .PE_OUT    (PE352_PE_OUT[31:0]              ), //o
    .finish    (PE352_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE353 (
    .activate  (PE352_acount[7:0]               ), //i
    .weight    (PE253_bcount[7:0]               ), //i
    .valid     (PE353_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE353_acount[7:0]               ), //o
    .bcount    (PE353_bcount[7:0]               ), //o
    .PE_OUT    (PE353_PE_OUT[31:0]              ), //o
    .finish    (PE353_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE354 (
    .activate  (PE353_acount[7:0]               ), //i
    .weight    (PE254_bcount[7:0]               ), //i
    .valid     (PE354_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE354_acount[7:0]               ), //o
    .bcount    (PE354_bcount[7:0]               ), //o
    .PE_OUT    (PE354_PE_OUT[31:0]              ), //o
    .finish    (PE354_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE355 (
    .activate  (PE354_acount[7:0]               ), //i
    .weight    (PE255_bcount[7:0]               ), //i
    .valid     (PE355_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE355_acount[7:0]               ), //o
    .bcount    (PE355_bcount[7:0]               ), //o
    .PE_OUT    (PE355_PE_OUT[31:0]              ), //o
    .finish    (PE355_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE356 (
    .activate  (PE355_acount[7:0]               ), //i
    .weight    (PE256_bcount[7:0]               ), //i
    .valid     (PE356_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE356_acount[7:0]               ), //o
    .bcount    (PE356_bcount[7:0]               ), //o
    .PE_OUT    (PE356_PE_OUT[31:0]              ), //o
    .finish    (PE356_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE357 (
    .activate  (PE356_acount[7:0]               ), //i
    .weight    (PE257_bcount[7:0]               ), //i
    .valid     (PE357_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE357_acount[7:0]               ), //o
    .bcount    (PE357_bcount[7:0]               ), //o
    .PE_OUT    (PE357_PE_OUT[31:0]              ), //o
    .finish    (PE357_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE358 (
    .activate  (PE357_acount[7:0]               ), //i
    .weight    (PE258_bcount[7:0]               ), //i
    .valid     (PE358_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE358_acount[7:0]               ), //o
    .bcount    (PE358_bcount[7:0]               ), //o
    .PE_OUT    (PE358_PE_OUT[31:0]              ), //o
    .finish    (PE358_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE359 (
    .activate  (PE358_acount[7:0]               ), //i
    .weight    (PE259_bcount[7:0]               ), //i
    .valid     (PE359_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE359_acount[7:0]               ), //o
    .bcount    (PE359_bcount[7:0]               ), //o
    .PE_OUT    (PE359_PE_OUT[31:0]              ), //o
    .finish    (PE359_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE360 (
    .activate  (PE359_acount[7:0]               ), //i
    .weight    (PE260_bcount[7:0]               ), //i
    .valid     (PE360_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE360_acount[7:0]               ), //o
    .bcount    (PE360_bcount[7:0]               ), //o
    .PE_OUT    (PE360_PE_OUT[31:0]              ), //o
    .finish    (PE360_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE361 (
    .activate  (PE360_acount[7:0]               ), //i
    .weight    (PE261_bcount[7:0]               ), //i
    .valid     (PE361_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE361_acount[7:0]               ), //o
    .bcount    (PE361_bcount[7:0]               ), //o
    .PE_OUT    (PE361_PE_OUT[31:0]              ), //o
    .finish    (PE361_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE362 (
    .activate  (PE361_acount[7:0]               ), //i
    .weight    (PE262_bcount[7:0]               ), //i
    .valid     (PE362_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE362_acount[7:0]               ), //o
    .bcount    (PE362_bcount[7:0]               ), //o
    .PE_OUT    (PE362_PE_OUT[31:0]              ), //o
    .finish    (PE362_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE363 (
    .activate  (PE362_acount[7:0]               ), //i
    .weight    (PE263_bcount[7:0]               ), //i
    .valid     (PE363_valid                     ), //i
    .signCount (io_signCount_regNextWhen_3[15:0]), //i
    .acount    (PE363_acount[7:0]               ), //o
    .bcount    (PE363_bcount[7:0]               ), //o
    .PE_OUT    (PE363_PE_OUT[31:0]              ), //o
    .finish    (PE363_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE40 (
    .activate  (io_MatrixA_4[7:0]               ), //i
    .weight    (PE30_bcount[7:0]                ), //i
    .valid     (PE40_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE40_acount[7:0]                ), //o
    .bcount    (PE40_bcount[7:0]                ), //o
    .PE_OUT    (PE40_PE_OUT[31:0]               ), //o
    .finish    (PE40_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE41 (
    .activate  (PE40_acount[7:0]                ), //i
    .weight    (PE31_bcount[7:0]                ), //i
    .valid     (PE41_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE41_acount[7:0]                ), //o
    .bcount    (PE41_bcount[7:0]                ), //o
    .PE_OUT    (PE41_PE_OUT[31:0]               ), //o
    .finish    (PE41_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE42 (
    .activate  (PE41_acount[7:0]                ), //i
    .weight    (PE32_bcount[7:0]                ), //i
    .valid     (PE42_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE42_acount[7:0]                ), //o
    .bcount    (PE42_bcount[7:0]                ), //o
    .PE_OUT    (PE42_PE_OUT[31:0]               ), //o
    .finish    (PE42_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE43 (
    .activate  (PE42_acount[7:0]                ), //i
    .weight    (PE33_bcount[7:0]                ), //i
    .valid     (PE43_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE43_acount[7:0]                ), //o
    .bcount    (PE43_bcount[7:0]                ), //o
    .PE_OUT    (PE43_PE_OUT[31:0]               ), //o
    .finish    (PE43_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE44 (
    .activate  (PE43_acount[7:0]                ), //i
    .weight    (PE34_bcount[7:0]                ), //i
    .valid     (PE44_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE44_acount[7:0]                ), //o
    .bcount    (PE44_bcount[7:0]                ), //o
    .PE_OUT    (PE44_PE_OUT[31:0]               ), //o
    .finish    (PE44_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE45 (
    .activate  (PE44_acount[7:0]                ), //i
    .weight    (PE35_bcount[7:0]                ), //i
    .valid     (PE45_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE45_acount[7:0]                ), //o
    .bcount    (PE45_bcount[7:0]                ), //o
    .PE_OUT    (PE45_PE_OUT[31:0]               ), //o
    .finish    (PE45_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE46 (
    .activate  (PE45_acount[7:0]                ), //i
    .weight    (PE36_bcount[7:0]                ), //i
    .valid     (PE46_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE46_acount[7:0]                ), //o
    .bcount    (PE46_bcount[7:0]                ), //o
    .PE_OUT    (PE46_PE_OUT[31:0]               ), //o
    .finish    (PE46_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE47 (
    .activate  (PE46_acount[7:0]                ), //i
    .weight    (PE37_bcount[7:0]                ), //i
    .valid     (PE47_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE47_acount[7:0]                ), //o
    .bcount    (PE47_bcount[7:0]                ), //o
    .PE_OUT    (PE47_PE_OUT[31:0]               ), //o
    .finish    (PE47_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE48 (
    .activate  (PE47_acount[7:0]                ), //i
    .weight    (PE38_bcount[7:0]                ), //i
    .valid     (PE48_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE48_acount[7:0]                ), //o
    .bcount    (PE48_bcount[7:0]                ), //o
    .PE_OUT    (PE48_PE_OUT[31:0]               ), //o
    .finish    (PE48_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE49 (
    .activate  (PE48_acount[7:0]                ), //i
    .weight    (PE39_bcount[7:0]                ), //i
    .valid     (PE49_valid                      ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE49_acount[7:0]                ), //o
    .bcount    (PE49_bcount[7:0]                ), //o
    .PE_OUT    (PE49_PE_OUT[31:0]               ), //o
    .finish    (PE49_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE410 (
    .activate  (PE49_acount[7:0]                ), //i
    .weight    (PE310_bcount[7:0]               ), //i
    .valid     (PE410_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE410_acount[7:0]               ), //o
    .bcount    (PE410_bcount[7:0]               ), //o
    .PE_OUT    (PE410_PE_OUT[31:0]              ), //o
    .finish    (PE410_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE411 (
    .activate  (PE410_acount[7:0]               ), //i
    .weight    (PE311_bcount[7:0]               ), //i
    .valid     (PE411_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE411_acount[7:0]               ), //o
    .bcount    (PE411_bcount[7:0]               ), //o
    .PE_OUT    (PE411_PE_OUT[31:0]              ), //o
    .finish    (PE411_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE412 (
    .activate  (PE411_acount[7:0]               ), //i
    .weight    (PE312_bcount[7:0]               ), //i
    .valid     (PE412_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE412_acount[7:0]               ), //o
    .bcount    (PE412_bcount[7:0]               ), //o
    .PE_OUT    (PE412_PE_OUT[31:0]              ), //o
    .finish    (PE412_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE413 (
    .activate  (PE412_acount[7:0]               ), //i
    .weight    (PE313_bcount[7:0]               ), //i
    .valid     (PE413_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE413_acount[7:0]               ), //o
    .bcount    (PE413_bcount[7:0]               ), //o
    .PE_OUT    (PE413_PE_OUT[31:0]              ), //o
    .finish    (PE413_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE414 (
    .activate  (PE413_acount[7:0]               ), //i
    .weight    (PE314_bcount[7:0]               ), //i
    .valid     (PE414_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE414_acount[7:0]               ), //o
    .bcount    (PE414_bcount[7:0]               ), //o
    .PE_OUT    (PE414_PE_OUT[31:0]              ), //o
    .finish    (PE414_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE415 (
    .activate  (PE414_acount[7:0]               ), //i
    .weight    (PE315_bcount[7:0]               ), //i
    .valid     (PE415_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE415_acount[7:0]               ), //o
    .bcount    (PE415_bcount[7:0]               ), //o
    .PE_OUT    (PE415_PE_OUT[31:0]              ), //o
    .finish    (PE415_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE416 (
    .activate  (PE415_acount[7:0]               ), //i
    .weight    (PE316_bcount[7:0]               ), //i
    .valid     (PE416_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE416_acount[7:0]               ), //o
    .bcount    (PE416_bcount[7:0]               ), //o
    .PE_OUT    (PE416_PE_OUT[31:0]              ), //o
    .finish    (PE416_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE417 (
    .activate  (PE416_acount[7:0]               ), //i
    .weight    (PE317_bcount[7:0]               ), //i
    .valid     (PE417_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE417_acount[7:0]               ), //o
    .bcount    (PE417_bcount[7:0]               ), //o
    .PE_OUT    (PE417_PE_OUT[31:0]              ), //o
    .finish    (PE417_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE418 (
    .activate  (PE417_acount[7:0]               ), //i
    .weight    (PE318_bcount[7:0]               ), //i
    .valid     (PE418_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE418_acount[7:0]               ), //o
    .bcount    (PE418_bcount[7:0]               ), //o
    .PE_OUT    (PE418_PE_OUT[31:0]              ), //o
    .finish    (PE418_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE419 (
    .activate  (PE418_acount[7:0]               ), //i
    .weight    (PE319_bcount[7:0]               ), //i
    .valid     (PE419_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE419_acount[7:0]               ), //o
    .bcount    (PE419_bcount[7:0]               ), //o
    .PE_OUT    (PE419_PE_OUT[31:0]              ), //o
    .finish    (PE419_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE420 (
    .activate  (PE419_acount[7:0]               ), //i
    .weight    (PE320_bcount[7:0]               ), //i
    .valid     (PE420_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE420_acount[7:0]               ), //o
    .bcount    (PE420_bcount[7:0]               ), //o
    .PE_OUT    (PE420_PE_OUT[31:0]              ), //o
    .finish    (PE420_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE421 (
    .activate  (PE420_acount[7:0]               ), //i
    .weight    (PE321_bcount[7:0]               ), //i
    .valid     (PE421_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE421_acount[7:0]               ), //o
    .bcount    (PE421_bcount[7:0]               ), //o
    .PE_OUT    (PE421_PE_OUT[31:0]              ), //o
    .finish    (PE421_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE422 (
    .activate  (PE421_acount[7:0]               ), //i
    .weight    (PE322_bcount[7:0]               ), //i
    .valid     (PE422_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE422_acount[7:0]               ), //o
    .bcount    (PE422_bcount[7:0]               ), //o
    .PE_OUT    (PE422_PE_OUT[31:0]              ), //o
    .finish    (PE422_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE423 (
    .activate  (PE422_acount[7:0]               ), //i
    .weight    (PE323_bcount[7:0]               ), //i
    .valid     (PE423_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE423_acount[7:0]               ), //o
    .bcount    (PE423_bcount[7:0]               ), //o
    .PE_OUT    (PE423_PE_OUT[31:0]              ), //o
    .finish    (PE423_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE424 (
    .activate  (PE423_acount[7:0]               ), //i
    .weight    (PE324_bcount[7:0]               ), //i
    .valid     (PE424_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE424_acount[7:0]               ), //o
    .bcount    (PE424_bcount[7:0]               ), //o
    .PE_OUT    (PE424_PE_OUT[31:0]              ), //o
    .finish    (PE424_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE425 (
    .activate  (PE424_acount[7:0]               ), //i
    .weight    (PE325_bcount[7:0]               ), //i
    .valid     (PE425_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE425_acount[7:0]               ), //o
    .bcount    (PE425_bcount[7:0]               ), //o
    .PE_OUT    (PE425_PE_OUT[31:0]              ), //o
    .finish    (PE425_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE426 (
    .activate  (PE425_acount[7:0]               ), //i
    .weight    (PE326_bcount[7:0]               ), //i
    .valid     (PE426_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE426_acount[7:0]               ), //o
    .bcount    (PE426_bcount[7:0]               ), //o
    .PE_OUT    (PE426_PE_OUT[31:0]              ), //o
    .finish    (PE426_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE427 (
    .activate  (PE426_acount[7:0]               ), //i
    .weight    (PE327_bcount[7:0]               ), //i
    .valid     (PE427_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE427_acount[7:0]               ), //o
    .bcount    (PE427_bcount[7:0]               ), //o
    .PE_OUT    (PE427_PE_OUT[31:0]              ), //o
    .finish    (PE427_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE428 (
    .activate  (PE427_acount[7:0]               ), //i
    .weight    (PE328_bcount[7:0]               ), //i
    .valid     (PE428_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE428_acount[7:0]               ), //o
    .bcount    (PE428_bcount[7:0]               ), //o
    .PE_OUT    (PE428_PE_OUT[31:0]              ), //o
    .finish    (PE428_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE429 (
    .activate  (PE428_acount[7:0]               ), //i
    .weight    (PE329_bcount[7:0]               ), //i
    .valid     (PE429_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE429_acount[7:0]               ), //o
    .bcount    (PE429_bcount[7:0]               ), //o
    .PE_OUT    (PE429_PE_OUT[31:0]              ), //o
    .finish    (PE429_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE430 (
    .activate  (PE429_acount[7:0]               ), //i
    .weight    (PE330_bcount[7:0]               ), //i
    .valid     (PE430_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE430_acount[7:0]               ), //o
    .bcount    (PE430_bcount[7:0]               ), //o
    .PE_OUT    (PE430_PE_OUT[31:0]              ), //o
    .finish    (PE430_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE431 (
    .activate  (PE430_acount[7:0]               ), //i
    .weight    (PE331_bcount[7:0]               ), //i
    .valid     (PE431_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE431_acount[7:0]               ), //o
    .bcount    (PE431_bcount[7:0]               ), //o
    .PE_OUT    (PE431_PE_OUT[31:0]              ), //o
    .finish    (PE431_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE432 (
    .activate  (PE431_acount[7:0]               ), //i
    .weight    (PE332_bcount[7:0]               ), //i
    .valid     (PE432_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE432_acount[7:0]               ), //o
    .bcount    (PE432_bcount[7:0]               ), //o
    .PE_OUT    (PE432_PE_OUT[31:0]              ), //o
    .finish    (PE432_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE433 (
    .activate  (PE432_acount[7:0]               ), //i
    .weight    (PE333_bcount[7:0]               ), //i
    .valid     (PE433_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE433_acount[7:0]               ), //o
    .bcount    (PE433_bcount[7:0]               ), //o
    .PE_OUT    (PE433_PE_OUT[31:0]              ), //o
    .finish    (PE433_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE434 (
    .activate  (PE433_acount[7:0]               ), //i
    .weight    (PE334_bcount[7:0]               ), //i
    .valid     (PE434_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE434_acount[7:0]               ), //o
    .bcount    (PE434_bcount[7:0]               ), //o
    .PE_OUT    (PE434_PE_OUT[31:0]              ), //o
    .finish    (PE434_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE435 (
    .activate  (PE434_acount[7:0]               ), //i
    .weight    (PE335_bcount[7:0]               ), //i
    .valid     (PE435_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE435_acount[7:0]               ), //o
    .bcount    (PE435_bcount[7:0]               ), //o
    .PE_OUT    (PE435_PE_OUT[31:0]              ), //o
    .finish    (PE435_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE436 (
    .activate  (PE435_acount[7:0]               ), //i
    .weight    (PE336_bcount[7:0]               ), //i
    .valid     (PE436_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE436_acount[7:0]               ), //o
    .bcount    (PE436_bcount[7:0]               ), //o
    .PE_OUT    (PE436_PE_OUT[31:0]              ), //o
    .finish    (PE436_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE437 (
    .activate  (PE436_acount[7:0]               ), //i
    .weight    (PE337_bcount[7:0]               ), //i
    .valid     (PE437_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE437_acount[7:0]               ), //o
    .bcount    (PE437_bcount[7:0]               ), //o
    .PE_OUT    (PE437_PE_OUT[31:0]              ), //o
    .finish    (PE437_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE438 (
    .activate  (PE437_acount[7:0]               ), //i
    .weight    (PE338_bcount[7:0]               ), //i
    .valid     (PE438_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE438_acount[7:0]               ), //o
    .bcount    (PE438_bcount[7:0]               ), //o
    .PE_OUT    (PE438_PE_OUT[31:0]              ), //o
    .finish    (PE438_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE439 (
    .activate  (PE438_acount[7:0]               ), //i
    .weight    (PE339_bcount[7:0]               ), //i
    .valid     (PE439_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE439_acount[7:0]               ), //o
    .bcount    (PE439_bcount[7:0]               ), //o
    .PE_OUT    (PE439_PE_OUT[31:0]              ), //o
    .finish    (PE439_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE440 (
    .activate  (PE439_acount[7:0]               ), //i
    .weight    (PE340_bcount[7:0]               ), //i
    .valid     (PE440_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE440_acount[7:0]               ), //o
    .bcount    (PE440_bcount[7:0]               ), //o
    .PE_OUT    (PE440_PE_OUT[31:0]              ), //o
    .finish    (PE440_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE441 (
    .activate  (PE440_acount[7:0]               ), //i
    .weight    (PE341_bcount[7:0]               ), //i
    .valid     (PE441_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE441_acount[7:0]               ), //o
    .bcount    (PE441_bcount[7:0]               ), //o
    .PE_OUT    (PE441_PE_OUT[31:0]              ), //o
    .finish    (PE441_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE442 (
    .activate  (PE441_acount[7:0]               ), //i
    .weight    (PE342_bcount[7:0]               ), //i
    .valid     (PE442_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE442_acount[7:0]               ), //o
    .bcount    (PE442_bcount[7:0]               ), //o
    .PE_OUT    (PE442_PE_OUT[31:0]              ), //o
    .finish    (PE442_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE443 (
    .activate  (PE442_acount[7:0]               ), //i
    .weight    (PE343_bcount[7:0]               ), //i
    .valid     (PE443_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE443_acount[7:0]               ), //o
    .bcount    (PE443_bcount[7:0]               ), //o
    .PE_OUT    (PE443_PE_OUT[31:0]              ), //o
    .finish    (PE443_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE444 (
    .activate  (PE443_acount[7:0]               ), //i
    .weight    (PE344_bcount[7:0]               ), //i
    .valid     (PE444_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE444_acount[7:0]               ), //o
    .bcount    (PE444_bcount[7:0]               ), //o
    .PE_OUT    (PE444_PE_OUT[31:0]              ), //o
    .finish    (PE444_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE445 (
    .activate  (PE444_acount[7:0]               ), //i
    .weight    (PE345_bcount[7:0]               ), //i
    .valid     (PE445_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE445_acount[7:0]               ), //o
    .bcount    (PE445_bcount[7:0]               ), //o
    .PE_OUT    (PE445_PE_OUT[31:0]              ), //o
    .finish    (PE445_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE446 (
    .activate  (PE445_acount[7:0]               ), //i
    .weight    (PE346_bcount[7:0]               ), //i
    .valid     (PE446_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE446_acount[7:0]               ), //o
    .bcount    (PE446_bcount[7:0]               ), //o
    .PE_OUT    (PE446_PE_OUT[31:0]              ), //o
    .finish    (PE446_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE447 (
    .activate  (PE446_acount[7:0]               ), //i
    .weight    (PE347_bcount[7:0]               ), //i
    .valid     (PE447_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE447_acount[7:0]               ), //o
    .bcount    (PE447_bcount[7:0]               ), //o
    .PE_OUT    (PE447_PE_OUT[31:0]              ), //o
    .finish    (PE447_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE448 (
    .activate  (PE447_acount[7:0]               ), //i
    .weight    (PE348_bcount[7:0]               ), //i
    .valid     (PE448_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE448_acount[7:0]               ), //o
    .bcount    (PE448_bcount[7:0]               ), //o
    .PE_OUT    (PE448_PE_OUT[31:0]              ), //o
    .finish    (PE448_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE449 (
    .activate  (PE448_acount[7:0]               ), //i
    .weight    (PE349_bcount[7:0]               ), //i
    .valid     (PE449_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE449_acount[7:0]               ), //o
    .bcount    (PE449_bcount[7:0]               ), //o
    .PE_OUT    (PE449_PE_OUT[31:0]              ), //o
    .finish    (PE449_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE450 (
    .activate  (PE449_acount[7:0]               ), //i
    .weight    (PE350_bcount[7:0]               ), //i
    .valid     (PE450_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE450_acount[7:0]               ), //o
    .bcount    (PE450_bcount[7:0]               ), //o
    .PE_OUT    (PE450_PE_OUT[31:0]              ), //o
    .finish    (PE450_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE451 (
    .activate  (PE450_acount[7:0]               ), //i
    .weight    (PE351_bcount[7:0]               ), //i
    .valid     (PE451_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE451_acount[7:0]               ), //o
    .bcount    (PE451_bcount[7:0]               ), //o
    .PE_OUT    (PE451_PE_OUT[31:0]              ), //o
    .finish    (PE451_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE452 (
    .activate  (PE451_acount[7:0]               ), //i
    .weight    (PE352_bcount[7:0]               ), //i
    .valid     (PE452_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE452_acount[7:0]               ), //o
    .bcount    (PE452_bcount[7:0]               ), //o
    .PE_OUT    (PE452_PE_OUT[31:0]              ), //o
    .finish    (PE452_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE453 (
    .activate  (PE452_acount[7:0]               ), //i
    .weight    (PE353_bcount[7:0]               ), //i
    .valid     (PE453_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE453_acount[7:0]               ), //o
    .bcount    (PE453_bcount[7:0]               ), //o
    .PE_OUT    (PE453_PE_OUT[31:0]              ), //o
    .finish    (PE453_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE454 (
    .activate  (PE453_acount[7:0]               ), //i
    .weight    (PE354_bcount[7:0]               ), //i
    .valid     (PE454_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE454_acount[7:0]               ), //o
    .bcount    (PE454_bcount[7:0]               ), //o
    .PE_OUT    (PE454_PE_OUT[31:0]              ), //o
    .finish    (PE454_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE455 (
    .activate  (PE454_acount[7:0]               ), //i
    .weight    (PE355_bcount[7:0]               ), //i
    .valid     (PE455_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE455_acount[7:0]               ), //o
    .bcount    (PE455_bcount[7:0]               ), //o
    .PE_OUT    (PE455_PE_OUT[31:0]              ), //o
    .finish    (PE455_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE456 (
    .activate  (PE455_acount[7:0]               ), //i
    .weight    (PE356_bcount[7:0]               ), //i
    .valid     (PE456_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE456_acount[7:0]               ), //o
    .bcount    (PE456_bcount[7:0]               ), //o
    .PE_OUT    (PE456_PE_OUT[31:0]              ), //o
    .finish    (PE456_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE457 (
    .activate  (PE456_acount[7:0]               ), //i
    .weight    (PE357_bcount[7:0]               ), //i
    .valid     (PE457_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE457_acount[7:0]               ), //o
    .bcount    (PE457_bcount[7:0]               ), //o
    .PE_OUT    (PE457_PE_OUT[31:0]              ), //o
    .finish    (PE457_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE458 (
    .activate  (PE457_acount[7:0]               ), //i
    .weight    (PE358_bcount[7:0]               ), //i
    .valid     (PE458_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE458_acount[7:0]               ), //o
    .bcount    (PE458_bcount[7:0]               ), //o
    .PE_OUT    (PE458_PE_OUT[31:0]              ), //o
    .finish    (PE458_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE459 (
    .activate  (PE458_acount[7:0]               ), //i
    .weight    (PE359_bcount[7:0]               ), //i
    .valid     (PE459_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE459_acount[7:0]               ), //o
    .bcount    (PE459_bcount[7:0]               ), //o
    .PE_OUT    (PE459_PE_OUT[31:0]              ), //o
    .finish    (PE459_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE460 (
    .activate  (PE459_acount[7:0]               ), //i
    .weight    (PE360_bcount[7:0]               ), //i
    .valid     (PE460_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE460_acount[7:0]               ), //o
    .bcount    (PE460_bcount[7:0]               ), //o
    .PE_OUT    (PE460_PE_OUT[31:0]              ), //o
    .finish    (PE460_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE461 (
    .activate  (PE460_acount[7:0]               ), //i
    .weight    (PE361_bcount[7:0]               ), //i
    .valid     (PE461_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE461_acount[7:0]               ), //o
    .bcount    (PE461_bcount[7:0]               ), //o
    .PE_OUT    (PE461_PE_OUT[31:0]              ), //o
    .finish    (PE461_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE462 (
    .activate  (PE461_acount[7:0]               ), //i
    .weight    (PE362_bcount[7:0]               ), //i
    .valid     (PE462_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE462_acount[7:0]               ), //o
    .bcount    (PE462_bcount[7:0]               ), //o
    .PE_OUT    (PE462_PE_OUT[31:0]              ), //o
    .finish    (PE462_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE463 (
    .activate  (PE462_acount[7:0]               ), //i
    .weight    (PE363_bcount[7:0]               ), //i
    .valid     (PE463_valid                     ), //i
    .signCount (io_signCount_regNextWhen_4[15:0]), //i
    .acount    (PE463_acount[7:0]               ), //o
    .bcount    (PE463_bcount[7:0]               ), //o
    .PE_OUT    (PE463_PE_OUT[31:0]              ), //o
    .finish    (PE463_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE50 (
    .activate  (io_MatrixA_5[7:0]               ), //i
    .weight    (PE40_bcount[7:0]                ), //i
    .valid     (PE50_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE50_acount[7:0]                ), //o
    .bcount    (PE50_bcount[7:0]                ), //o
    .PE_OUT    (PE50_PE_OUT[31:0]               ), //o
    .finish    (PE50_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE51 (
    .activate  (PE50_acount[7:0]                ), //i
    .weight    (PE41_bcount[7:0]                ), //i
    .valid     (PE51_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE51_acount[7:0]                ), //o
    .bcount    (PE51_bcount[7:0]                ), //o
    .PE_OUT    (PE51_PE_OUT[31:0]               ), //o
    .finish    (PE51_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE52 (
    .activate  (PE51_acount[7:0]                ), //i
    .weight    (PE42_bcount[7:0]                ), //i
    .valid     (PE52_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE52_acount[7:0]                ), //o
    .bcount    (PE52_bcount[7:0]                ), //o
    .PE_OUT    (PE52_PE_OUT[31:0]               ), //o
    .finish    (PE52_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE53 (
    .activate  (PE52_acount[7:0]                ), //i
    .weight    (PE43_bcount[7:0]                ), //i
    .valid     (PE53_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE53_acount[7:0]                ), //o
    .bcount    (PE53_bcount[7:0]                ), //o
    .PE_OUT    (PE53_PE_OUT[31:0]               ), //o
    .finish    (PE53_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE54 (
    .activate  (PE53_acount[7:0]                ), //i
    .weight    (PE44_bcount[7:0]                ), //i
    .valid     (PE54_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE54_acount[7:0]                ), //o
    .bcount    (PE54_bcount[7:0]                ), //o
    .PE_OUT    (PE54_PE_OUT[31:0]               ), //o
    .finish    (PE54_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE55 (
    .activate  (PE54_acount[7:0]                ), //i
    .weight    (PE45_bcount[7:0]                ), //i
    .valid     (PE55_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE55_acount[7:0]                ), //o
    .bcount    (PE55_bcount[7:0]                ), //o
    .PE_OUT    (PE55_PE_OUT[31:0]               ), //o
    .finish    (PE55_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE56 (
    .activate  (PE55_acount[7:0]                ), //i
    .weight    (PE46_bcount[7:0]                ), //i
    .valid     (PE56_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE56_acount[7:0]                ), //o
    .bcount    (PE56_bcount[7:0]                ), //o
    .PE_OUT    (PE56_PE_OUT[31:0]               ), //o
    .finish    (PE56_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE57 (
    .activate  (PE56_acount[7:0]                ), //i
    .weight    (PE47_bcount[7:0]                ), //i
    .valid     (PE57_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE57_acount[7:0]                ), //o
    .bcount    (PE57_bcount[7:0]                ), //o
    .PE_OUT    (PE57_PE_OUT[31:0]               ), //o
    .finish    (PE57_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE58 (
    .activate  (PE57_acount[7:0]                ), //i
    .weight    (PE48_bcount[7:0]                ), //i
    .valid     (PE58_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE58_acount[7:0]                ), //o
    .bcount    (PE58_bcount[7:0]                ), //o
    .PE_OUT    (PE58_PE_OUT[31:0]               ), //o
    .finish    (PE58_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE59 (
    .activate  (PE58_acount[7:0]                ), //i
    .weight    (PE49_bcount[7:0]                ), //i
    .valid     (PE59_valid                      ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE59_acount[7:0]                ), //o
    .bcount    (PE59_bcount[7:0]                ), //o
    .PE_OUT    (PE59_PE_OUT[31:0]               ), //o
    .finish    (PE59_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE510 (
    .activate  (PE59_acount[7:0]                ), //i
    .weight    (PE410_bcount[7:0]               ), //i
    .valid     (PE510_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE510_acount[7:0]               ), //o
    .bcount    (PE510_bcount[7:0]               ), //o
    .PE_OUT    (PE510_PE_OUT[31:0]              ), //o
    .finish    (PE510_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE511 (
    .activate  (PE510_acount[7:0]               ), //i
    .weight    (PE411_bcount[7:0]               ), //i
    .valid     (PE511_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE511_acount[7:0]               ), //o
    .bcount    (PE511_bcount[7:0]               ), //o
    .PE_OUT    (PE511_PE_OUT[31:0]              ), //o
    .finish    (PE511_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE512 (
    .activate  (PE511_acount[7:0]               ), //i
    .weight    (PE412_bcount[7:0]               ), //i
    .valid     (PE512_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE512_acount[7:0]               ), //o
    .bcount    (PE512_bcount[7:0]               ), //o
    .PE_OUT    (PE512_PE_OUT[31:0]              ), //o
    .finish    (PE512_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE513 (
    .activate  (PE512_acount[7:0]               ), //i
    .weight    (PE413_bcount[7:0]               ), //i
    .valid     (PE513_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE513_acount[7:0]               ), //o
    .bcount    (PE513_bcount[7:0]               ), //o
    .PE_OUT    (PE513_PE_OUT[31:0]              ), //o
    .finish    (PE513_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE514 (
    .activate  (PE513_acount[7:0]               ), //i
    .weight    (PE414_bcount[7:0]               ), //i
    .valid     (PE514_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE514_acount[7:0]               ), //o
    .bcount    (PE514_bcount[7:0]               ), //o
    .PE_OUT    (PE514_PE_OUT[31:0]              ), //o
    .finish    (PE514_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE515 (
    .activate  (PE514_acount[7:0]               ), //i
    .weight    (PE415_bcount[7:0]               ), //i
    .valid     (PE515_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE515_acount[7:0]               ), //o
    .bcount    (PE515_bcount[7:0]               ), //o
    .PE_OUT    (PE515_PE_OUT[31:0]              ), //o
    .finish    (PE515_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE516 (
    .activate  (PE515_acount[7:0]               ), //i
    .weight    (PE416_bcount[7:0]               ), //i
    .valid     (PE516_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE516_acount[7:0]               ), //o
    .bcount    (PE516_bcount[7:0]               ), //o
    .PE_OUT    (PE516_PE_OUT[31:0]              ), //o
    .finish    (PE516_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE517 (
    .activate  (PE516_acount[7:0]               ), //i
    .weight    (PE417_bcount[7:0]               ), //i
    .valid     (PE517_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE517_acount[7:0]               ), //o
    .bcount    (PE517_bcount[7:0]               ), //o
    .PE_OUT    (PE517_PE_OUT[31:0]              ), //o
    .finish    (PE517_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE518 (
    .activate  (PE517_acount[7:0]               ), //i
    .weight    (PE418_bcount[7:0]               ), //i
    .valid     (PE518_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE518_acount[7:0]               ), //o
    .bcount    (PE518_bcount[7:0]               ), //o
    .PE_OUT    (PE518_PE_OUT[31:0]              ), //o
    .finish    (PE518_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE519 (
    .activate  (PE518_acount[7:0]               ), //i
    .weight    (PE419_bcount[7:0]               ), //i
    .valid     (PE519_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE519_acount[7:0]               ), //o
    .bcount    (PE519_bcount[7:0]               ), //o
    .PE_OUT    (PE519_PE_OUT[31:0]              ), //o
    .finish    (PE519_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE520 (
    .activate  (PE519_acount[7:0]               ), //i
    .weight    (PE420_bcount[7:0]               ), //i
    .valid     (PE520_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE520_acount[7:0]               ), //o
    .bcount    (PE520_bcount[7:0]               ), //o
    .PE_OUT    (PE520_PE_OUT[31:0]              ), //o
    .finish    (PE520_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE521 (
    .activate  (PE520_acount[7:0]               ), //i
    .weight    (PE421_bcount[7:0]               ), //i
    .valid     (PE521_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE521_acount[7:0]               ), //o
    .bcount    (PE521_bcount[7:0]               ), //o
    .PE_OUT    (PE521_PE_OUT[31:0]              ), //o
    .finish    (PE521_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE522 (
    .activate  (PE521_acount[7:0]               ), //i
    .weight    (PE422_bcount[7:0]               ), //i
    .valid     (PE522_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE522_acount[7:0]               ), //o
    .bcount    (PE522_bcount[7:0]               ), //o
    .PE_OUT    (PE522_PE_OUT[31:0]              ), //o
    .finish    (PE522_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE523 (
    .activate  (PE522_acount[7:0]               ), //i
    .weight    (PE423_bcount[7:0]               ), //i
    .valid     (PE523_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE523_acount[7:0]               ), //o
    .bcount    (PE523_bcount[7:0]               ), //o
    .PE_OUT    (PE523_PE_OUT[31:0]              ), //o
    .finish    (PE523_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE524 (
    .activate  (PE523_acount[7:0]               ), //i
    .weight    (PE424_bcount[7:0]               ), //i
    .valid     (PE524_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE524_acount[7:0]               ), //o
    .bcount    (PE524_bcount[7:0]               ), //o
    .PE_OUT    (PE524_PE_OUT[31:0]              ), //o
    .finish    (PE524_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE525 (
    .activate  (PE524_acount[7:0]               ), //i
    .weight    (PE425_bcount[7:0]               ), //i
    .valid     (PE525_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE525_acount[7:0]               ), //o
    .bcount    (PE525_bcount[7:0]               ), //o
    .PE_OUT    (PE525_PE_OUT[31:0]              ), //o
    .finish    (PE525_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE526 (
    .activate  (PE525_acount[7:0]               ), //i
    .weight    (PE426_bcount[7:0]               ), //i
    .valid     (PE526_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE526_acount[7:0]               ), //o
    .bcount    (PE526_bcount[7:0]               ), //o
    .PE_OUT    (PE526_PE_OUT[31:0]              ), //o
    .finish    (PE526_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE527 (
    .activate  (PE526_acount[7:0]               ), //i
    .weight    (PE427_bcount[7:0]               ), //i
    .valid     (PE527_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE527_acount[7:0]               ), //o
    .bcount    (PE527_bcount[7:0]               ), //o
    .PE_OUT    (PE527_PE_OUT[31:0]              ), //o
    .finish    (PE527_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE528 (
    .activate  (PE527_acount[7:0]               ), //i
    .weight    (PE428_bcount[7:0]               ), //i
    .valid     (PE528_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE528_acount[7:0]               ), //o
    .bcount    (PE528_bcount[7:0]               ), //o
    .PE_OUT    (PE528_PE_OUT[31:0]              ), //o
    .finish    (PE528_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE529 (
    .activate  (PE528_acount[7:0]               ), //i
    .weight    (PE429_bcount[7:0]               ), //i
    .valid     (PE529_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE529_acount[7:0]               ), //o
    .bcount    (PE529_bcount[7:0]               ), //o
    .PE_OUT    (PE529_PE_OUT[31:0]              ), //o
    .finish    (PE529_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE530 (
    .activate  (PE529_acount[7:0]               ), //i
    .weight    (PE430_bcount[7:0]               ), //i
    .valid     (PE530_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE530_acount[7:0]               ), //o
    .bcount    (PE530_bcount[7:0]               ), //o
    .PE_OUT    (PE530_PE_OUT[31:0]              ), //o
    .finish    (PE530_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE531 (
    .activate  (PE530_acount[7:0]               ), //i
    .weight    (PE431_bcount[7:0]               ), //i
    .valid     (PE531_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE531_acount[7:0]               ), //o
    .bcount    (PE531_bcount[7:0]               ), //o
    .PE_OUT    (PE531_PE_OUT[31:0]              ), //o
    .finish    (PE531_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE532 (
    .activate  (PE531_acount[7:0]               ), //i
    .weight    (PE432_bcount[7:0]               ), //i
    .valid     (PE532_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE532_acount[7:0]               ), //o
    .bcount    (PE532_bcount[7:0]               ), //o
    .PE_OUT    (PE532_PE_OUT[31:0]              ), //o
    .finish    (PE532_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE533 (
    .activate  (PE532_acount[7:0]               ), //i
    .weight    (PE433_bcount[7:0]               ), //i
    .valid     (PE533_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE533_acount[7:0]               ), //o
    .bcount    (PE533_bcount[7:0]               ), //o
    .PE_OUT    (PE533_PE_OUT[31:0]              ), //o
    .finish    (PE533_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE534 (
    .activate  (PE533_acount[7:0]               ), //i
    .weight    (PE434_bcount[7:0]               ), //i
    .valid     (PE534_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE534_acount[7:0]               ), //o
    .bcount    (PE534_bcount[7:0]               ), //o
    .PE_OUT    (PE534_PE_OUT[31:0]              ), //o
    .finish    (PE534_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE535 (
    .activate  (PE534_acount[7:0]               ), //i
    .weight    (PE435_bcount[7:0]               ), //i
    .valid     (PE535_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE535_acount[7:0]               ), //o
    .bcount    (PE535_bcount[7:0]               ), //o
    .PE_OUT    (PE535_PE_OUT[31:0]              ), //o
    .finish    (PE535_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE536 (
    .activate  (PE535_acount[7:0]               ), //i
    .weight    (PE436_bcount[7:0]               ), //i
    .valid     (PE536_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE536_acount[7:0]               ), //o
    .bcount    (PE536_bcount[7:0]               ), //o
    .PE_OUT    (PE536_PE_OUT[31:0]              ), //o
    .finish    (PE536_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE537 (
    .activate  (PE536_acount[7:0]               ), //i
    .weight    (PE437_bcount[7:0]               ), //i
    .valid     (PE537_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE537_acount[7:0]               ), //o
    .bcount    (PE537_bcount[7:0]               ), //o
    .PE_OUT    (PE537_PE_OUT[31:0]              ), //o
    .finish    (PE537_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE538 (
    .activate  (PE537_acount[7:0]               ), //i
    .weight    (PE438_bcount[7:0]               ), //i
    .valid     (PE538_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE538_acount[7:0]               ), //o
    .bcount    (PE538_bcount[7:0]               ), //o
    .PE_OUT    (PE538_PE_OUT[31:0]              ), //o
    .finish    (PE538_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE539 (
    .activate  (PE538_acount[7:0]               ), //i
    .weight    (PE439_bcount[7:0]               ), //i
    .valid     (PE539_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE539_acount[7:0]               ), //o
    .bcount    (PE539_bcount[7:0]               ), //o
    .PE_OUT    (PE539_PE_OUT[31:0]              ), //o
    .finish    (PE539_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE540 (
    .activate  (PE539_acount[7:0]               ), //i
    .weight    (PE440_bcount[7:0]               ), //i
    .valid     (PE540_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE540_acount[7:0]               ), //o
    .bcount    (PE540_bcount[7:0]               ), //o
    .PE_OUT    (PE540_PE_OUT[31:0]              ), //o
    .finish    (PE540_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE541 (
    .activate  (PE540_acount[7:0]               ), //i
    .weight    (PE441_bcount[7:0]               ), //i
    .valid     (PE541_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE541_acount[7:0]               ), //o
    .bcount    (PE541_bcount[7:0]               ), //o
    .PE_OUT    (PE541_PE_OUT[31:0]              ), //o
    .finish    (PE541_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE542 (
    .activate  (PE541_acount[7:0]               ), //i
    .weight    (PE442_bcount[7:0]               ), //i
    .valid     (PE542_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE542_acount[7:0]               ), //o
    .bcount    (PE542_bcount[7:0]               ), //o
    .PE_OUT    (PE542_PE_OUT[31:0]              ), //o
    .finish    (PE542_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE543 (
    .activate  (PE542_acount[7:0]               ), //i
    .weight    (PE443_bcount[7:0]               ), //i
    .valid     (PE543_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE543_acount[7:0]               ), //o
    .bcount    (PE543_bcount[7:0]               ), //o
    .PE_OUT    (PE543_PE_OUT[31:0]              ), //o
    .finish    (PE543_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE544 (
    .activate  (PE543_acount[7:0]               ), //i
    .weight    (PE444_bcount[7:0]               ), //i
    .valid     (PE544_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE544_acount[7:0]               ), //o
    .bcount    (PE544_bcount[7:0]               ), //o
    .PE_OUT    (PE544_PE_OUT[31:0]              ), //o
    .finish    (PE544_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE545 (
    .activate  (PE544_acount[7:0]               ), //i
    .weight    (PE445_bcount[7:0]               ), //i
    .valid     (PE545_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE545_acount[7:0]               ), //o
    .bcount    (PE545_bcount[7:0]               ), //o
    .PE_OUT    (PE545_PE_OUT[31:0]              ), //o
    .finish    (PE545_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE546 (
    .activate  (PE545_acount[7:0]               ), //i
    .weight    (PE446_bcount[7:0]               ), //i
    .valid     (PE546_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE546_acount[7:0]               ), //o
    .bcount    (PE546_bcount[7:0]               ), //o
    .PE_OUT    (PE546_PE_OUT[31:0]              ), //o
    .finish    (PE546_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE547 (
    .activate  (PE546_acount[7:0]               ), //i
    .weight    (PE447_bcount[7:0]               ), //i
    .valid     (PE547_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE547_acount[7:0]               ), //o
    .bcount    (PE547_bcount[7:0]               ), //o
    .PE_OUT    (PE547_PE_OUT[31:0]              ), //o
    .finish    (PE547_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE548 (
    .activate  (PE547_acount[7:0]               ), //i
    .weight    (PE448_bcount[7:0]               ), //i
    .valid     (PE548_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE548_acount[7:0]               ), //o
    .bcount    (PE548_bcount[7:0]               ), //o
    .PE_OUT    (PE548_PE_OUT[31:0]              ), //o
    .finish    (PE548_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE549 (
    .activate  (PE548_acount[7:0]               ), //i
    .weight    (PE449_bcount[7:0]               ), //i
    .valid     (PE549_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE549_acount[7:0]               ), //o
    .bcount    (PE549_bcount[7:0]               ), //o
    .PE_OUT    (PE549_PE_OUT[31:0]              ), //o
    .finish    (PE549_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE550 (
    .activate  (PE549_acount[7:0]               ), //i
    .weight    (PE450_bcount[7:0]               ), //i
    .valid     (PE550_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE550_acount[7:0]               ), //o
    .bcount    (PE550_bcount[7:0]               ), //o
    .PE_OUT    (PE550_PE_OUT[31:0]              ), //o
    .finish    (PE550_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE551 (
    .activate  (PE550_acount[7:0]               ), //i
    .weight    (PE451_bcount[7:0]               ), //i
    .valid     (PE551_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE551_acount[7:0]               ), //o
    .bcount    (PE551_bcount[7:0]               ), //o
    .PE_OUT    (PE551_PE_OUT[31:0]              ), //o
    .finish    (PE551_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE552 (
    .activate  (PE551_acount[7:0]               ), //i
    .weight    (PE452_bcount[7:0]               ), //i
    .valid     (PE552_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE552_acount[7:0]               ), //o
    .bcount    (PE552_bcount[7:0]               ), //o
    .PE_OUT    (PE552_PE_OUT[31:0]              ), //o
    .finish    (PE552_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE553 (
    .activate  (PE552_acount[7:0]               ), //i
    .weight    (PE453_bcount[7:0]               ), //i
    .valid     (PE553_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE553_acount[7:0]               ), //o
    .bcount    (PE553_bcount[7:0]               ), //o
    .PE_OUT    (PE553_PE_OUT[31:0]              ), //o
    .finish    (PE553_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE554 (
    .activate  (PE553_acount[7:0]               ), //i
    .weight    (PE454_bcount[7:0]               ), //i
    .valid     (PE554_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE554_acount[7:0]               ), //o
    .bcount    (PE554_bcount[7:0]               ), //o
    .PE_OUT    (PE554_PE_OUT[31:0]              ), //o
    .finish    (PE554_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE555 (
    .activate  (PE554_acount[7:0]               ), //i
    .weight    (PE455_bcount[7:0]               ), //i
    .valid     (PE555_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE555_acount[7:0]               ), //o
    .bcount    (PE555_bcount[7:0]               ), //o
    .PE_OUT    (PE555_PE_OUT[31:0]              ), //o
    .finish    (PE555_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE556 (
    .activate  (PE555_acount[7:0]               ), //i
    .weight    (PE456_bcount[7:0]               ), //i
    .valid     (PE556_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE556_acount[7:0]               ), //o
    .bcount    (PE556_bcount[7:0]               ), //o
    .PE_OUT    (PE556_PE_OUT[31:0]              ), //o
    .finish    (PE556_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE557 (
    .activate  (PE556_acount[7:0]               ), //i
    .weight    (PE457_bcount[7:0]               ), //i
    .valid     (PE557_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE557_acount[7:0]               ), //o
    .bcount    (PE557_bcount[7:0]               ), //o
    .PE_OUT    (PE557_PE_OUT[31:0]              ), //o
    .finish    (PE557_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE558 (
    .activate  (PE557_acount[7:0]               ), //i
    .weight    (PE458_bcount[7:0]               ), //i
    .valid     (PE558_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE558_acount[7:0]               ), //o
    .bcount    (PE558_bcount[7:0]               ), //o
    .PE_OUT    (PE558_PE_OUT[31:0]              ), //o
    .finish    (PE558_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE559 (
    .activate  (PE558_acount[7:0]               ), //i
    .weight    (PE459_bcount[7:0]               ), //i
    .valid     (PE559_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE559_acount[7:0]               ), //o
    .bcount    (PE559_bcount[7:0]               ), //o
    .PE_OUT    (PE559_PE_OUT[31:0]              ), //o
    .finish    (PE559_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE560 (
    .activate  (PE559_acount[7:0]               ), //i
    .weight    (PE460_bcount[7:0]               ), //i
    .valid     (PE560_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE560_acount[7:0]               ), //o
    .bcount    (PE560_bcount[7:0]               ), //o
    .PE_OUT    (PE560_PE_OUT[31:0]              ), //o
    .finish    (PE560_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE561 (
    .activate  (PE560_acount[7:0]               ), //i
    .weight    (PE461_bcount[7:0]               ), //i
    .valid     (PE561_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE561_acount[7:0]               ), //o
    .bcount    (PE561_bcount[7:0]               ), //o
    .PE_OUT    (PE561_PE_OUT[31:0]              ), //o
    .finish    (PE561_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE562 (
    .activate  (PE561_acount[7:0]               ), //i
    .weight    (PE462_bcount[7:0]               ), //i
    .valid     (PE562_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE562_acount[7:0]               ), //o
    .bcount    (PE562_bcount[7:0]               ), //o
    .PE_OUT    (PE562_PE_OUT[31:0]              ), //o
    .finish    (PE562_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE563 (
    .activate  (PE562_acount[7:0]               ), //i
    .weight    (PE463_bcount[7:0]               ), //i
    .valid     (PE563_valid                     ), //i
    .signCount (io_signCount_regNextWhen_5[15:0]), //i
    .acount    (PE563_acount[7:0]               ), //o
    .bcount    (PE563_bcount[7:0]               ), //o
    .PE_OUT    (PE563_PE_OUT[31:0]              ), //o
    .finish    (PE563_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE60 (
    .activate  (io_MatrixA_6[7:0]               ), //i
    .weight    (PE50_bcount[7:0]                ), //i
    .valid     (PE60_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE60_acount[7:0]                ), //o
    .bcount    (PE60_bcount[7:0]                ), //o
    .PE_OUT    (PE60_PE_OUT[31:0]               ), //o
    .finish    (PE60_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE61 (
    .activate  (PE60_acount[7:0]                ), //i
    .weight    (PE51_bcount[7:0]                ), //i
    .valid     (PE61_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE61_acount[7:0]                ), //o
    .bcount    (PE61_bcount[7:0]                ), //o
    .PE_OUT    (PE61_PE_OUT[31:0]               ), //o
    .finish    (PE61_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE62 (
    .activate  (PE61_acount[7:0]                ), //i
    .weight    (PE52_bcount[7:0]                ), //i
    .valid     (PE62_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE62_acount[7:0]                ), //o
    .bcount    (PE62_bcount[7:0]                ), //o
    .PE_OUT    (PE62_PE_OUT[31:0]               ), //o
    .finish    (PE62_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE63 (
    .activate  (PE62_acount[7:0]                ), //i
    .weight    (PE53_bcount[7:0]                ), //i
    .valid     (PE63_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE63_acount[7:0]                ), //o
    .bcount    (PE63_bcount[7:0]                ), //o
    .PE_OUT    (PE63_PE_OUT[31:0]               ), //o
    .finish    (PE63_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE64 (
    .activate  (PE63_acount[7:0]                ), //i
    .weight    (PE54_bcount[7:0]                ), //i
    .valid     (PE64_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE64_acount[7:0]                ), //o
    .bcount    (PE64_bcount[7:0]                ), //o
    .PE_OUT    (PE64_PE_OUT[31:0]               ), //o
    .finish    (PE64_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE65 (
    .activate  (PE64_acount[7:0]                ), //i
    .weight    (PE55_bcount[7:0]                ), //i
    .valid     (PE65_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE65_acount[7:0]                ), //o
    .bcount    (PE65_bcount[7:0]                ), //o
    .PE_OUT    (PE65_PE_OUT[31:0]               ), //o
    .finish    (PE65_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE66 (
    .activate  (PE65_acount[7:0]                ), //i
    .weight    (PE56_bcount[7:0]                ), //i
    .valid     (PE66_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE66_acount[7:0]                ), //o
    .bcount    (PE66_bcount[7:0]                ), //o
    .PE_OUT    (PE66_PE_OUT[31:0]               ), //o
    .finish    (PE66_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE67 (
    .activate  (PE66_acount[7:0]                ), //i
    .weight    (PE57_bcount[7:0]                ), //i
    .valid     (PE67_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE67_acount[7:0]                ), //o
    .bcount    (PE67_bcount[7:0]                ), //o
    .PE_OUT    (PE67_PE_OUT[31:0]               ), //o
    .finish    (PE67_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE68 (
    .activate  (PE67_acount[7:0]                ), //i
    .weight    (PE58_bcount[7:0]                ), //i
    .valid     (PE68_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE68_acount[7:0]                ), //o
    .bcount    (PE68_bcount[7:0]                ), //o
    .PE_OUT    (PE68_PE_OUT[31:0]               ), //o
    .finish    (PE68_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE69 (
    .activate  (PE68_acount[7:0]                ), //i
    .weight    (PE59_bcount[7:0]                ), //i
    .valid     (PE69_valid                      ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE69_acount[7:0]                ), //o
    .bcount    (PE69_bcount[7:0]                ), //o
    .PE_OUT    (PE69_PE_OUT[31:0]               ), //o
    .finish    (PE69_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE610 (
    .activate  (PE69_acount[7:0]                ), //i
    .weight    (PE510_bcount[7:0]               ), //i
    .valid     (PE610_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE610_acount[7:0]               ), //o
    .bcount    (PE610_bcount[7:0]               ), //o
    .PE_OUT    (PE610_PE_OUT[31:0]              ), //o
    .finish    (PE610_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE611 (
    .activate  (PE610_acount[7:0]               ), //i
    .weight    (PE511_bcount[7:0]               ), //i
    .valid     (PE611_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE611_acount[7:0]               ), //o
    .bcount    (PE611_bcount[7:0]               ), //o
    .PE_OUT    (PE611_PE_OUT[31:0]              ), //o
    .finish    (PE611_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE612 (
    .activate  (PE611_acount[7:0]               ), //i
    .weight    (PE512_bcount[7:0]               ), //i
    .valid     (PE612_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE612_acount[7:0]               ), //o
    .bcount    (PE612_bcount[7:0]               ), //o
    .PE_OUT    (PE612_PE_OUT[31:0]              ), //o
    .finish    (PE612_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE613 (
    .activate  (PE612_acount[7:0]               ), //i
    .weight    (PE513_bcount[7:0]               ), //i
    .valid     (PE613_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE613_acount[7:0]               ), //o
    .bcount    (PE613_bcount[7:0]               ), //o
    .PE_OUT    (PE613_PE_OUT[31:0]              ), //o
    .finish    (PE613_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE614 (
    .activate  (PE613_acount[7:0]               ), //i
    .weight    (PE514_bcount[7:0]               ), //i
    .valid     (PE614_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE614_acount[7:0]               ), //o
    .bcount    (PE614_bcount[7:0]               ), //o
    .PE_OUT    (PE614_PE_OUT[31:0]              ), //o
    .finish    (PE614_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE615 (
    .activate  (PE614_acount[7:0]               ), //i
    .weight    (PE515_bcount[7:0]               ), //i
    .valid     (PE615_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE615_acount[7:0]               ), //o
    .bcount    (PE615_bcount[7:0]               ), //o
    .PE_OUT    (PE615_PE_OUT[31:0]              ), //o
    .finish    (PE615_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE616 (
    .activate  (PE615_acount[7:0]               ), //i
    .weight    (PE516_bcount[7:0]               ), //i
    .valid     (PE616_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE616_acount[7:0]               ), //o
    .bcount    (PE616_bcount[7:0]               ), //o
    .PE_OUT    (PE616_PE_OUT[31:0]              ), //o
    .finish    (PE616_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE617 (
    .activate  (PE616_acount[7:0]               ), //i
    .weight    (PE517_bcount[7:0]               ), //i
    .valid     (PE617_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE617_acount[7:0]               ), //o
    .bcount    (PE617_bcount[7:0]               ), //o
    .PE_OUT    (PE617_PE_OUT[31:0]              ), //o
    .finish    (PE617_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE618 (
    .activate  (PE617_acount[7:0]               ), //i
    .weight    (PE518_bcount[7:0]               ), //i
    .valid     (PE618_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE618_acount[7:0]               ), //o
    .bcount    (PE618_bcount[7:0]               ), //o
    .PE_OUT    (PE618_PE_OUT[31:0]              ), //o
    .finish    (PE618_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE619 (
    .activate  (PE618_acount[7:0]               ), //i
    .weight    (PE519_bcount[7:0]               ), //i
    .valid     (PE619_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE619_acount[7:0]               ), //o
    .bcount    (PE619_bcount[7:0]               ), //o
    .PE_OUT    (PE619_PE_OUT[31:0]              ), //o
    .finish    (PE619_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE620 (
    .activate  (PE619_acount[7:0]               ), //i
    .weight    (PE520_bcount[7:0]               ), //i
    .valid     (PE620_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE620_acount[7:0]               ), //o
    .bcount    (PE620_bcount[7:0]               ), //o
    .PE_OUT    (PE620_PE_OUT[31:0]              ), //o
    .finish    (PE620_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE621 (
    .activate  (PE620_acount[7:0]               ), //i
    .weight    (PE521_bcount[7:0]               ), //i
    .valid     (PE621_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE621_acount[7:0]               ), //o
    .bcount    (PE621_bcount[7:0]               ), //o
    .PE_OUT    (PE621_PE_OUT[31:0]              ), //o
    .finish    (PE621_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE622 (
    .activate  (PE621_acount[7:0]               ), //i
    .weight    (PE522_bcount[7:0]               ), //i
    .valid     (PE622_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE622_acount[7:0]               ), //o
    .bcount    (PE622_bcount[7:0]               ), //o
    .PE_OUT    (PE622_PE_OUT[31:0]              ), //o
    .finish    (PE622_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE623 (
    .activate  (PE622_acount[7:0]               ), //i
    .weight    (PE523_bcount[7:0]               ), //i
    .valid     (PE623_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE623_acount[7:0]               ), //o
    .bcount    (PE623_bcount[7:0]               ), //o
    .PE_OUT    (PE623_PE_OUT[31:0]              ), //o
    .finish    (PE623_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE624 (
    .activate  (PE623_acount[7:0]               ), //i
    .weight    (PE524_bcount[7:0]               ), //i
    .valid     (PE624_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE624_acount[7:0]               ), //o
    .bcount    (PE624_bcount[7:0]               ), //o
    .PE_OUT    (PE624_PE_OUT[31:0]              ), //o
    .finish    (PE624_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE625 (
    .activate  (PE624_acount[7:0]               ), //i
    .weight    (PE525_bcount[7:0]               ), //i
    .valid     (PE625_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE625_acount[7:0]               ), //o
    .bcount    (PE625_bcount[7:0]               ), //o
    .PE_OUT    (PE625_PE_OUT[31:0]              ), //o
    .finish    (PE625_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE626 (
    .activate  (PE625_acount[7:0]               ), //i
    .weight    (PE526_bcount[7:0]               ), //i
    .valid     (PE626_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE626_acount[7:0]               ), //o
    .bcount    (PE626_bcount[7:0]               ), //o
    .PE_OUT    (PE626_PE_OUT[31:0]              ), //o
    .finish    (PE626_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE627 (
    .activate  (PE626_acount[7:0]               ), //i
    .weight    (PE527_bcount[7:0]               ), //i
    .valid     (PE627_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE627_acount[7:0]               ), //o
    .bcount    (PE627_bcount[7:0]               ), //o
    .PE_OUT    (PE627_PE_OUT[31:0]              ), //o
    .finish    (PE627_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE628 (
    .activate  (PE627_acount[7:0]               ), //i
    .weight    (PE528_bcount[7:0]               ), //i
    .valid     (PE628_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE628_acount[7:0]               ), //o
    .bcount    (PE628_bcount[7:0]               ), //o
    .PE_OUT    (PE628_PE_OUT[31:0]              ), //o
    .finish    (PE628_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE629 (
    .activate  (PE628_acount[7:0]               ), //i
    .weight    (PE529_bcount[7:0]               ), //i
    .valid     (PE629_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE629_acount[7:0]               ), //o
    .bcount    (PE629_bcount[7:0]               ), //o
    .PE_OUT    (PE629_PE_OUT[31:0]              ), //o
    .finish    (PE629_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE630 (
    .activate  (PE629_acount[7:0]               ), //i
    .weight    (PE530_bcount[7:0]               ), //i
    .valid     (PE630_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE630_acount[7:0]               ), //o
    .bcount    (PE630_bcount[7:0]               ), //o
    .PE_OUT    (PE630_PE_OUT[31:0]              ), //o
    .finish    (PE630_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE631 (
    .activate  (PE630_acount[7:0]               ), //i
    .weight    (PE531_bcount[7:0]               ), //i
    .valid     (PE631_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE631_acount[7:0]               ), //o
    .bcount    (PE631_bcount[7:0]               ), //o
    .PE_OUT    (PE631_PE_OUT[31:0]              ), //o
    .finish    (PE631_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE632 (
    .activate  (PE631_acount[7:0]               ), //i
    .weight    (PE532_bcount[7:0]               ), //i
    .valid     (PE632_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE632_acount[7:0]               ), //o
    .bcount    (PE632_bcount[7:0]               ), //o
    .PE_OUT    (PE632_PE_OUT[31:0]              ), //o
    .finish    (PE632_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE633 (
    .activate  (PE632_acount[7:0]               ), //i
    .weight    (PE533_bcount[7:0]               ), //i
    .valid     (PE633_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE633_acount[7:0]               ), //o
    .bcount    (PE633_bcount[7:0]               ), //o
    .PE_OUT    (PE633_PE_OUT[31:0]              ), //o
    .finish    (PE633_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE634 (
    .activate  (PE633_acount[7:0]               ), //i
    .weight    (PE534_bcount[7:0]               ), //i
    .valid     (PE634_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE634_acount[7:0]               ), //o
    .bcount    (PE634_bcount[7:0]               ), //o
    .PE_OUT    (PE634_PE_OUT[31:0]              ), //o
    .finish    (PE634_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE635 (
    .activate  (PE634_acount[7:0]               ), //i
    .weight    (PE535_bcount[7:0]               ), //i
    .valid     (PE635_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE635_acount[7:0]               ), //o
    .bcount    (PE635_bcount[7:0]               ), //o
    .PE_OUT    (PE635_PE_OUT[31:0]              ), //o
    .finish    (PE635_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE636 (
    .activate  (PE635_acount[7:0]               ), //i
    .weight    (PE536_bcount[7:0]               ), //i
    .valid     (PE636_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE636_acount[7:0]               ), //o
    .bcount    (PE636_bcount[7:0]               ), //o
    .PE_OUT    (PE636_PE_OUT[31:0]              ), //o
    .finish    (PE636_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE637 (
    .activate  (PE636_acount[7:0]               ), //i
    .weight    (PE537_bcount[7:0]               ), //i
    .valid     (PE637_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE637_acount[7:0]               ), //o
    .bcount    (PE637_bcount[7:0]               ), //o
    .PE_OUT    (PE637_PE_OUT[31:0]              ), //o
    .finish    (PE637_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE638 (
    .activate  (PE637_acount[7:0]               ), //i
    .weight    (PE538_bcount[7:0]               ), //i
    .valid     (PE638_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE638_acount[7:0]               ), //o
    .bcount    (PE638_bcount[7:0]               ), //o
    .PE_OUT    (PE638_PE_OUT[31:0]              ), //o
    .finish    (PE638_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE639 (
    .activate  (PE638_acount[7:0]               ), //i
    .weight    (PE539_bcount[7:0]               ), //i
    .valid     (PE639_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE639_acount[7:0]               ), //o
    .bcount    (PE639_bcount[7:0]               ), //o
    .PE_OUT    (PE639_PE_OUT[31:0]              ), //o
    .finish    (PE639_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE640 (
    .activate  (PE639_acount[7:0]               ), //i
    .weight    (PE540_bcount[7:0]               ), //i
    .valid     (PE640_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE640_acount[7:0]               ), //o
    .bcount    (PE640_bcount[7:0]               ), //o
    .PE_OUT    (PE640_PE_OUT[31:0]              ), //o
    .finish    (PE640_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE641 (
    .activate  (PE640_acount[7:0]               ), //i
    .weight    (PE541_bcount[7:0]               ), //i
    .valid     (PE641_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE641_acount[7:0]               ), //o
    .bcount    (PE641_bcount[7:0]               ), //o
    .PE_OUT    (PE641_PE_OUT[31:0]              ), //o
    .finish    (PE641_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE642 (
    .activate  (PE641_acount[7:0]               ), //i
    .weight    (PE542_bcount[7:0]               ), //i
    .valid     (PE642_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE642_acount[7:0]               ), //o
    .bcount    (PE642_bcount[7:0]               ), //o
    .PE_OUT    (PE642_PE_OUT[31:0]              ), //o
    .finish    (PE642_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE643 (
    .activate  (PE642_acount[7:0]               ), //i
    .weight    (PE543_bcount[7:0]               ), //i
    .valid     (PE643_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE643_acount[7:0]               ), //o
    .bcount    (PE643_bcount[7:0]               ), //o
    .PE_OUT    (PE643_PE_OUT[31:0]              ), //o
    .finish    (PE643_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE644 (
    .activate  (PE643_acount[7:0]               ), //i
    .weight    (PE544_bcount[7:0]               ), //i
    .valid     (PE644_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE644_acount[7:0]               ), //o
    .bcount    (PE644_bcount[7:0]               ), //o
    .PE_OUT    (PE644_PE_OUT[31:0]              ), //o
    .finish    (PE644_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE645 (
    .activate  (PE644_acount[7:0]               ), //i
    .weight    (PE545_bcount[7:0]               ), //i
    .valid     (PE645_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE645_acount[7:0]               ), //o
    .bcount    (PE645_bcount[7:0]               ), //o
    .PE_OUT    (PE645_PE_OUT[31:0]              ), //o
    .finish    (PE645_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE646 (
    .activate  (PE645_acount[7:0]               ), //i
    .weight    (PE546_bcount[7:0]               ), //i
    .valid     (PE646_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE646_acount[7:0]               ), //o
    .bcount    (PE646_bcount[7:0]               ), //o
    .PE_OUT    (PE646_PE_OUT[31:0]              ), //o
    .finish    (PE646_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE647 (
    .activate  (PE646_acount[7:0]               ), //i
    .weight    (PE547_bcount[7:0]               ), //i
    .valid     (PE647_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE647_acount[7:0]               ), //o
    .bcount    (PE647_bcount[7:0]               ), //o
    .PE_OUT    (PE647_PE_OUT[31:0]              ), //o
    .finish    (PE647_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE648 (
    .activate  (PE647_acount[7:0]               ), //i
    .weight    (PE548_bcount[7:0]               ), //i
    .valid     (PE648_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE648_acount[7:0]               ), //o
    .bcount    (PE648_bcount[7:0]               ), //o
    .PE_OUT    (PE648_PE_OUT[31:0]              ), //o
    .finish    (PE648_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE649 (
    .activate  (PE648_acount[7:0]               ), //i
    .weight    (PE549_bcount[7:0]               ), //i
    .valid     (PE649_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE649_acount[7:0]               ), //o
    .bcount    (PE649_bcount[7:0]               ), //o
    .PE_OUT    (PE649_PE_OUT[31:0]              ), //o
    .finish    (PE649_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE650 (
    .activate  (PE649_acount[7:0]               ), //i
    .weight    (PE550_bcount[7:0]               ), //i
    .valid     (PE650_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE650_acount[7:0]               ), //o
    .bcount    (PE650_bcount[7:0]               ), //o
    .PE_OUT    (PE650_PE_OUT[31:0]              ), //o
    .finish    (PE650_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE651 (
    .activate  (PE650_acount[7:0]               ), //i
    .weight    (PE551_bcount[7:0]               ), //i
    .valid     (PE651_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE651_acount[7:0]               ), //o
    .bcount    (PE651_bcount[7:0]               ), //o
    .PE_OUT    (PE651_PE_OUT[31:0]              ), //o
    .finish    (PE651_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE652 (
    .activate  (PE651_acount[7:0]               ), //i
    .weight    (PE552_bcount[7:0]               ), //i
    .valid     (PE652_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE652_acount[7:0]               ), //o
    .bcount    (PE652_bcount[7:0]               ), //o
    .PE_OUT    (PE652_PE_OUT[31:0]              ), //o
    .finish    (PE652_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE653 (
    .activate  (PE652_acount[7:0]               ), //i
    .weight    (PE553_bcount[7:0]               ), //i
    .valid     (PE653_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE653_acount[7:0]               ), //o
    .bcount    (PE653_bcount[7:0]               ), //o
    .PE_OUT    (PE653_PE_OUT[31:0]              ), //o
    .finish    (PE653_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE654 (
    .activate  (PE653_acount[7:0]               ), //i
    .weight    (PE554_bcount[7:0]               ), //i
    .valid     (PE654_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE654_acount[7:0]               ), //o
    .bcount    (PE654_bcount[7:0]               ), //o
    .PE_OUT    (PE654_PE_OUT[31:0]              ), //o
    .finish    (PE654_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE655 (
    .activate  (PE654_acount[7:0]               ), //i
    .weight    (PE555_bcount[7:0]               ), //i
    .valid     (PE655_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE655_acount[7:0]               ), //o
    .bcount    (PE655_bcount[7:0]               ), //o
    .PE_OUT    (PE655_PE_OUT[31:0]              ), //o
    .finish    (PE655_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE656 (
    .activate  (PE655_acount[7:0]               ), //i
    .weight    (PE556_bcount[7:0]               ), //i
    .valid     (PE656_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE656_acount[7:0]               ), //o
    .bcount    (PE656_bcount[7:0]               ), //o
    .PE_OUT    (PE656_PE_OUT[31:0]              ), //o
    .finish    (PE656_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE657 (
    .activate  (PE656_acount[7:0]               ), //i
    .weight    (PE557_bcount[7:0]               ), //i
    .valid     (PE657_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE657_acount[7:0]               ), //o
    .bcount    (PE657_bcount[7:0]               ), //o
    .PE_OUT    (PE657_PE_OUT[31:0]              ), //o
    .finish    (PE657_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE658 (
    .activate  (PE657_acount[7:0]               ), //i
    .weight    (PE558_bcount[7:0]               ), //i
    .valid     (PE658_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE658_acount[7:0]               ), //o
    .bcount    (PE658_bcount[7:0]               ), //o
    .PE_OUT    (PE658_PE_OUT[31:0]              ), //o
    .finish    (PE658_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE659 (
    .activate  (PE658_acount[7:0]               ), //i
    .weight    (PE559_bcount[7:0]               ), //i
    .valid     (PE659_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE659_acount[7:0]               ), //o
    .bcount    (PE659_bcount[7:0]               ), //o
    .PE_OUT    (PE659_PE_OUT[31:0]              ), //o
    .finish    (PE659_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE660 (
    .activate  (PE659_acount[7:0]               ), //i
    .weight    (PE560_bcount[7:0]               ), //i
    .valid     (PE660_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE660_acount[7:0]               ), //o
    .bcount    (PE660_bcount[7:0]               ), //o
    .PE_OUT    (PE660_PE_OUT[31:0]              ), //o
    .finish    (PE660_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE661 (
    .activate  (PE660_acount[7:0]               ), //i
    .weight    (PE561_bcount[7:0]               ), //i
    .valid     (PE661_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE661_acount[7:0]               ), //o
    .bcount    (PE661_bcount[7:0]               ), //o
    .PE_OUT    (PE661_PE_OUT[31:0]              ), //o
    .finish    (PE661_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE662 (
    .activate  (PE661_acount[7:0]               ), //i
    .weight    (PE562_bcount[7:0]               ), //i
    .valid     (PE662_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE662_acount[7:0]               ), //o
    .bcount    (PE662_bcount[7:0]               ), //o
    .PE_OUT    (PE662_PE_OUT[31:0]              ), //o
    .finish    (PE662_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE663 (
    .activate  (PE662_acount[7:0]               ), //i
    .weight    (PE563_bcount[7:0]               ), //i
    .valid     (PE663_valid                     ), //i
    .signCount (io_signCount_regNextWhen_6[15:0]), //i
    .acount    (PE663_acount[7:0]               ), //o
    .bcount    (PE663_bcount[7:0]               ), //o
    .PE_OUT    (PE663_PE_OUT[31:0]              ), //o
    .finish    (PE663_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE70 (
    .activate  (io_MatrixA_7[7:0]               ), //i
    .weight    (PE60_bcount[7:0]                ), //i
    .valid     (PE70_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE70_acount[7:0]                ), //o
    .bcount    (PE70_bcount[7:0]                ), //o
    .PE_OUT    (PE70_PE_OUT[31:0]               ), //o
    .finish    (PE70_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE71 (
    .activate  (PE70_acount[7:0]                ), //i
    .weight    (PE61_bcount[7:0]                ), //i
    .valid     (PE71_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE71_acount[7:0]                ), //o
    .bcount    (PE71_bcount[7:0]                ), //o
    .PE_OUT    (PE71_PE_OUT[31:0]               ), //o
    .finish    (PE71_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE72 (
    .activate  (PE71_acount[7:0]                ), //i
    .weight    (PE62_bcount[7:0]                ), //i
    .valid     (PE72_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE72_acount[7:0]                ), //o
    .bcount    (PE72_bcount[7:0]                ), //o
    .PE_OUT    (PE72_PE_OUT[31:0]               ), //o
    .finish    (PE72_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE73 (
    .activate  (PE72_acount[7:0]                ), //i
    .weight    (PE63_bcount[7:0]                ), //i
    .valid     (PE73_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE73_acount[7:0]                ), //o
    .bcount    (PE73_bcount[7:0]                ), //o
    .PE_OUT    (PE73_PE_OUT[31:0]               ), //o
    .finish    (PE73_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE74 (
    .activate  (PE73_acount[7:0]                ), //i
    .weight    (PE64_bcount[7:0]                ), //i
    .valid     (PE74_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE74_acount[7:0]                ), //o
    .bcount    (PE74_bcount[7:0]                ), //o
    .PE_OUT    (PE74_PE_OUT[31:0]               ), //o
    .finish    (PE74_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE75 (
    .activate  (PE74_acount[7:0]                ), //i
    .weight    (PE65_bcount[7:0]                ), //i
    .valid     (PE75_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE75_acount[7:0]                ), //o
    .bcount    (PE75_bcount[7:0]                ), //o
    .PE_OUT    (PE75_PE_OUT[31:0]               ), //o
    .finish    (PE75_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE76 (
    .activate  (PE75_acount[7:0]                ), //i
    .weight    (PE66_bcount[7:0]                ), //i
    .valid     (PE76_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE76_acount[7:0]                ), //o
    .bcount    (PE76_bcount[7:0]                ), //o
    .PE_OUT    (PE76_PE_OUT[31:0]               ), //o
    .finish    (PE76_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE77 (
    .activate  (PE76_acount[7:0]                ), //i
    .weight    (PE67_bcount[7:0]                ), //i
    .valid     (PE77_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE77_acount[7:0]                ), //o
    .bcount    (PE77_bcount[7:0]                ), //o
    .PE_OUT    (PE77_PE_OUT[31:0]               ), //o
    .finish    (PE77_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE78 (
    .activate  (PE77_acount[7:0]                ), //i
    .weight    (PE68_bcount[7:0]                ), //i
    .valid     (PE78_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE78_acount[7:0]                ), //o
    .bcount    (PE78_bcount[7:0]                ), //o
    .PE_OUT    (PE78_PE_OUT[31:0]               ), //o
    .finish    (PE78_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE79 (
    .activate  (PE78_acount[7:0]                ), //i
    .weight    (PE69_bcount[7:0]                ), //i
    .valid     (PE79_valid                      ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE79_acount[7:0]                ), //o
    .bcount    (PE79_bcount[7:0]                ), //o
    .PE_OUT    (PE79_PE_OUT[31:0]               ), //o
    .finish    (PE79_finish                     ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE710 (
    .activate  (PE79_acount[7:0]                ), //i
    .weight    (PE610_bcount[7:0]               ), //i
    .valid     (PE710_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE710_acount[7:0]               ), //o
    .bcount    (PE710_bcount[7:0]               ), //o
    .PE_OUT    (PE710_PE_OUT[31:0]              ), //o
    .finish    (PE710_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE711 (
    .activate  (PE710_acount[7:0]               ), //i
    .weight    (PE611_bcount[7:0]               ), //i
    .valid     (PE711_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE711_acount[7:0]               ), //o
    .bcount    (PE711_bcount[7:0]               ), //o
    .PE_OUT    (PE711_PE_OUT[31:0]              ), //o
    .finish    (PE711_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE712 (
    .activate  (PE711_acount[7:0]               ), //i
    .weight    (PE612_bcount[7:0]               ), //i
    .valid     (PE712_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE712_acount[7:0]               ), //o
    .bcount    (PE712_bcount[7:0]               ), //o
    .PE_OUT    (PE712_PE_OUT[31:0]              ), //o
    .finish    (PE712_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE713 (
    .activate  (PE712_acount[7:0]               ), //i
    .weight    (PE613_bcount[7:0]               ), //i
    .valid     (PE713_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE713_acount[7:0]               ), //o
    .bcount    (PE713_bcount[7:0]               ), //o
    .PE_OUT    (PE713_PE_OUT[31:0]              ), //o
    .finish    (PE713_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE714 (
    .activate  (PE713_acount[7:0]               ), //i
    .weight    (PE614_bcount[7:0]               ), //i
    .valid     (PE714_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE714_acount[7:0]               ), //o
    .bcount    (PE714_bcount[7:0]               ), //o
    .PE_OUT    (PE714_PE_OUT[31:0]              ), //o
    .finish    (PE714_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE715 (
    .activate  (PE714_acount[7:0]               ), //i
    .weight    (PE615_bcount[7:0]               ), //i
    .valid     (PE715_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE715_acount[7:0]               ), //o
    .bcount    (PE715_bcount[7:0]               ), //o
    .PE_OUT    (PE715_PE_OUT[31:0]              ), //o
    .finish    (PE715_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE716 (
    .activate  (PE715_acount[7:0]               ), //i
    .weight    (PE616_bcount[7:0]               ), //i
    .valid     (PE716_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE716_acount[7:0]               ), //o
    .bcount    (PE716_bcount[7:0]               ), //o
    .PE_OUT    (PE716_PE_OUT[31:0]              ), //o
    .finish    (PE716_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE717 (
    .activate  (PE716_acount[7:0]               ), //i
    .weight    (PE617_bcount[7:0]               ), //i
    .valid     (PE717_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE717_acount[7:0]               ), //o
    .bcount    (PE717_bcount[7:0]               ), //o
    .PE_OUT    (PE717_PE_OUT[31:0]              ), //o
    .finish    (PE717_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE718 (
    .activate  (PE717_acount[7:0]               ), //i
    .weight    (PE618_bcount[7:0]               ), //i
    .valid     (PE718_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE718_acount[7:0]               ), //o
    .bcount    (PE718_bcount[7:0]               ), //o
    .PE_OUT    (PE718_PE_OUT[31:0]              ), //o
    .finish    (PE718_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE719 (
    .activate  (PE718_acount[7:0]               ), //i
    .weight    (PE619_bcount[7:0]               ), //i
    .valid     (PE719_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE719_acount[7:0]               ), //o
    .bcount    (PE719_bcount[7:0]               ), //o
    .PE_OUT    (PE719_PE_OUT[31:0]              ), //o
    .finish    (PE719_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE720 (
    .activate  (PE719_acount[7:0]               ), //i
    .weight    (PE620_bcount[7:0]               ), //i
    .valid     (PE720_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE720_acount[7:0]               ), //o
    .bcount    (PE720_bcount[7:0]               ), //o
    .PE_OUT    (PE720_PE_OUT[31:0]              ), //o
    .finish    (PE720_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE721 (
    .activate  (PE720_acount[7:0]               ), //i
    .weight    (PE621_bcount[7:0]               ), //i
    .valid     (PE721_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE721_acount[7:0]               ), //o
    .bcount    (PE721_bcount[7:0]               ), //o
    .PE_OUT    (PE721_PE_OUT[31:0]              ), //o
    .finish    (PE721_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE722 (
    .activate  (PE721_acount[7:0]               ), //i
    .weight    (PE622_bcount[7:0]               ), //i
    .valid     (PE722_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE722_acount[7:0]               ), //o
    .bcount    (PE722_bcount[7:0]               ), //o
    .PE_OUT    (PE722_PE_OUT[31:0]              ), //o
    .finish    (PE722_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE723 (
    .activate  (PE722_acount[7:0]               ), //i
    .weight    (PE623_bcount[7:0]               ), //i
    .valid     (PE723_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE723_acount[7:0]               ), //o
    .bcount    (PE723_bcount[7:0]               ), //o
    .PE_OUT    (PE723_PE_OUT[31:0]              ), //o
    .finish    (PE723_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE724 (
    .activate  (PE723_acount[7:0]               ), //i
    .weight    (PE624_bcount[7:0]               ), //i
    .valid     (PE724_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE724_acount[7:0]               ), //o
    .bcount    (PE724_bcount[7:0]               ), //o
    .PE_OUT    (PE724_PE_OUT[31:0]              ), //o
    .finish    (PE724_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE725 (
    .activate  (PE724_acount[7:0]               ), //i
    .weight    (PE625_bcount[7:0]               ), //i
    .valid     (PE725_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE725_acount[7:0]               ), //o
    .bcount    (PE725_bcount[7:0]               ), //o
    .PE_OUT    (PE725_PE_OUT[31:0]              ), //o
    .finish    (PE725_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE726 (
    .activate  (PE725_acount[7:0]               ), //i
    .weight    (PE626_bcount[7:0]               ), //i
    .valid     (PE726_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE726_acount[7:0]               ), //o
    .bcount    (PE726_bcount[7:0]               ), //o
    .PE_OUT    (PE726_PE_OUT[31:0]              ), //o
    .finish    (PE726_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE727 (
    .activate  (PE726_acount[7:0]               ), //i
    .weight    (PE627_bcount[7:0]               ), //i
    .valid     (PE727_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE727_acount[7:0]               ), //o
    .bcount    (PE727_bcount[7:0]               ), //o
    .PE_OUT    (PE727_PE_OUT[31:0]              ), //o
    .finish    (PE727_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE728 (
    .activate  (PE727_acount[7:0]               ), //i
    .weight    (PE628_bcount[7:0]               ), //i
    .valid     (PE728_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE728_acount[7:0]               ), //o
    .bcount    (PE728_bcount[7:0]               ), //o
    .PE_OUT    (PE728_PE_OUT[31:0]              ), //o
    .finish    (PE728_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE729 (
    .activate  (PE728_acount[7:0]               ), //i
    .weight    (PE629_bcount[7:0]               ), //i
    .valid     (PE729_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE729_acount[7:0]               ), //o
    .bcount    (PE729_bcount[7:0]               ), //o
    .PE_OUT    (PE729_PE_OUT[31:0]              ), //o
    .finish    (PE729_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE730 (
    .activate  (PE729_acount[7:0]               ), //i
    .weight    (PE630_bcount[7:0]               ), //i
    .valid     (PE730_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE730_acount[7:0]               ), //o
    .bcount    (PE730_bcount[7:0]               ), //o
    .PE_OUT    (PE730_PE_OUT[31:0]              ), //o
    .finish    (PE730_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE731 (
    .activate  (PE730_acount[7:0]               ), //i
    .weight    (PE631_bcount[7:0]               ), //i
    .valid     (PE731_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE731_acount[7:0]               ), //o
    .bcount    (PE731_bcount[7:0]               ), //o
    .PE_OUT    (PE731_PE_OUT[31:0]              ), //o
    .finish    (PE731_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE732 (
    .activate  (PE731_acount[7:0]               ), //i
    .weight    (PE632_bcount[7:0]               ), //i
    .valid     (PE732_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE732_acount[7:0]               ), //o
    .bcount    (PE732_bcount[7:0]               ), //o
    .PE_OUT    (PE732_PE_OUT[31:0]              ), //o
    .finish    (PE732_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE733 (
    .activate  (PE732_acount[7:0]               ), //i
    .weight    (PE633_bcount[7:0]               ), //i
    .valid     (PE733_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE733_acount[7:0]               ), //o
    .bcount    (PE733_bcount[7:0]               ), //o
    .PE_OUT    (PE733_PE_OUT[31:0]              ), //o
    .finish    (PE733_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE734 (
    .activate  (PE733_acount[7:0]               ), //i
    .weight    (PE634_bcount[7:0]               ), //i
    .valid     (PE734_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE734_acount[7:0]               ), //o
    .bcount    (PE734_bcount[7:0]               ), //o
    .PE_OUT    (PE734_PE_OUT[31:0]              ), //o
    .finish    (PE734_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE735 (
    .activate  (PE734_acount[7:0]               ), //i
    .weight    (PE635_bcount[7:0]               ), //i
    .valid     (PE735_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE735_acount[7:0]               ), //o
    .bcount    (PE735_bcount[7:0]               ), //o
    .PE_OUT    (PE735_PE_OUT[31:0]              ), //o
    .finish    (PE735_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE736 (
    .activate  (PE735_acount[7:0]               ), //i
    .weight    (PE636_bcount[7:0]               ), //i
    .valid     (PE736_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE736_acount[7:0]               ), //o
    .bcount    (PE736_bcount[7:0]               ), //o
    .PE_OUT    (PE736_PE_OUT[31:0]              ), //o
    .finish    (PE736_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE737 (
    .activate  (PE736_acount[7:0]               ), //i
    .weight    (PE637_bcount[7:0]               ), //i
    .valid     (PE737_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE737_acount[7:0]               ), //o
    .bcount    (PE737_bcount[7:0]               ), //o
    .PE_OUT    (PE737_PE_OUT[31:0]              ), //o
    .finish    (PE737_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE738 (
    .activate  (PE737_acount[7:0]               ), //i
    .weight    (PE638_bcount[7:0]               ), //i
    .valid     (PE738_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE738_acount[7:0]               ), //o
    .bcount    (PE738_bcount[7:0]               ), //o
    .PE_OUT    (PE738_PE_OUT[31:0]              ), //o
    .finish    (PE738_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE739 (
    .activate  (PE738_acount[7:0]               ), //i
    .weight    (PE639_bcount[7:0]               ), //i
    .valid     (PE739_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE739_acount[7:0]               ), //o
    .bcount    (PE739_bcount[7:0]               ), //o
    .PE_OUT    (PE739_PE_OUT[31:0]              ), //o
    .finish    (PE739_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE740 (
    .activate  (PE739_acount[7:0]               ), //i
    .weight    (PE640_bcount[7:0]               ), //i
    .valid     (PE740_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE740_acount[7:0]               ), //o
    .bcount    (PE740_bcount[7:0]               ), //o
    .PE_OUT    (PE740_PE_OUT[31:0]              ), //o
    .finish    (PE740_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE741 (
    .activate  (PE740_acount[7:0]               ), //i
    .weight    (PE641_bcount[7:0]               ), //i
    .valid     (PE741_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE741_acount[7:0]               ), //o
    .bcount    (PE741_bcount[7:0]               ), //o
    .PE_OUT    (PE741_PE_OUT[31:0]              ), //o
    .finish    (PE741_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE742 (
    .activate  (PE741_acount[7:0]               ), //i
    .weight    (PE642_bcount[7:0]               ), //i
    .valid     (PE742_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE742_acount[7:0]               ), //o
    .bcount    (PE742_bcount[7:0]               ), //o
    .PE_OUT    (PE742_PE_OUT[31:0]              ), //o
    .finish    (PE742_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE743 (
    .activate  (PE742_acount[7:0]               ), //i
    .weight    (PE643_bcount[7:0]               ), //i
    .valid     (PE743_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE743_acount[7:0]               ), //o
    .bcount    (PE743_bcount[7:0]               ), //o
    .PE_OUT    (PE743_PE_OUT[31:0]              ), //o
    .finish    (PE743_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE744 (
    .activate  (PE743_acount[7:0]               ), //i
    .weight    (PE644_bcount[7:0]               ), //i
    .valid     (PE744_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE744_acount[7:0]               ), //o
    .bcount    (PE744_bcount[7:0]               ), //o
    .PE_OUT    (PE744_PE_OUT[31:0]              ), //o
    .finish    (PE744_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE745 (
    .activate  (PE744_acount[7:0]               ), //i
    .weight    (PE645_bcount[7:0]               ), //i
    .valid     (PE745_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE745_acount[7:0]               ), //o
    .bcount    (PE745_bcount[7:0]               ), //o
    .PE_OUT    (PE745_PE_OUT[31:0]              ), //o
    .finish    (PE745_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE746 (
    .activate  (PE745_acount[7:0]               ), //i
    .weight    (PE646_bcount[7:0]               ), //i
    .valid     (PE746_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE746_acount[7:0]               ), //o
    .bcount    (PE746_bcount[7:0]               ), //o
    .PE_OUT    (PE746_PE_OUT[31:0]              ), //o
    .finish    (PE746_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE747 (
    .activate  (PE746_acount[7:0]               ), //i
    .weight    (PE647_bcount[7:0]               ), //i
    .valid     (PE747_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE747_acount[7:0]               ), //o
    .bcount    (PE747_bcount[7:0]               ), //o
    .PE_OUT    (PE747_PE_OUT[31:0]              ), //o
    .finish    (PE747_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE748 (
    .activate  (PE747_acount[7:0]               ), //i
    .weight    (PE648_bcount[7:0]               ), //i
    .valid     (PE748_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE748_acount[7:0]               ), //o
    .bcount    (PE748_bcount[7:0]               ), //o
    .PE_OUT    (PE748_PE_OUT[31:0]              ), //o
    .finish    (PE748_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE749 (
    .activate  (PE748_acount[7:0]               ), //i
    .weight    (PE649_bcount[7:0]               ), //i
    .valid     (PE749_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE749_acount[7:0]               ), //o
    .bcount    (PE749_bcount[7:0]               ), //o
    .PE_OUT    (PE749_PE_OUT[31:0]              ), //o
    .finish    (PE749_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE750 (
    .activate  (PE749_acount[7:0]               ), //i
    .weight    (PE650_bcount[7:0]               ), //i
    .valid     (PE750_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE750_acount[7:0]               ), //o
    .bcount    (PE750_bcount[7:0]               ), //o
    .PE_OUT    (PE750_PE_OUT[31:0]              ), //o
    .finish    (PE750_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE751 (
    .activate  (PE750_acount[7:0]               ), //i
    .weight    (PE651_bcount[7:0]               ), //i
    .valid     (PE751_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE751_acount[7:0]               ), //o
    .bcount    (PE751_bcount[7:0]               ), //o
    .PE_OUT    (PE751_PE_OUT[31:0]              ), //o
    .finish    (PE751_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE752 (
    .activate  (PE751_acount[7:0]               ), //i
    .weight    (PE652_bcount[7:0]               ), //i
    .valid     (PE752_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE752_acount[7:0]               ), //o
    .bcount    (PE752_bcount[7:0]               ), //o
    .PE_OUT    (PE752_PE_OUT[31:0]              ), //o
    .finish    (PE752_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE753 (
    .activate  (PE752_acount[7:0]               ), //i
    .weight    (PE653_bcount[7:0]               ), //i
    .valid     (PE753_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE753_acount[7:0]               ), //o
    .bcount    (PE753_bcount[7:0]               ), //o
    .PE_OUT    (PE753_PE_OUT[31:0]              ), //o
    .finish    (PE753_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE754 (
    .activate  (PE753_acount[7:0]               ), //i
    .weight    (PE654_bcount[7:0]               ), //i
    .valid     (PE754_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE754_acount[7:0]               ), //o
    .bcount    (PE754_bcount[7:0]               ), //o
    .PE_OUT    (PE754_PE_OUT[31:0]              ), //o
    .finish    (PE754_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE755 (
    .activate  (PE754_acount[7:0]               ), //i
    .weight    (PE655_bcount[7:0]               ), //i
    .valid     (PE755_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE755_acount[7:0]               ), //o
    .bcount    (PE755_bcount[7:0]               ), //o
    .PE_OUT    (PE755_PE_OUT[31:0]              ), //o
    .finish    (PE755_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE756 (
    .activate  (PE755_acount[7:0]               ), //i
    .weight    (PE656_bcount[7:0]               ), //i
    .valid     (PE756_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE756_acount[7:0]               ), //o
    .bcount    (PE756_bcount[7:0]               ), //o
    .PE_OUT    (PE756_PE_OUT[31:0]              ), //o
    .finish    (PE756_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE757 (
    .activate  (PE756_acount[7:0]               ), //i
    .weight    (PE657_bcount[7:0]               ), //i
    .valid     (PE757_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE757_acount[7:0]               ), //o
    .bcount    (PE757_bcount[7:0]               ), //o
    .PE_OUT    (PE757_PE_OUT[31:0]              ), //o
    .finish    (PE757_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE758 (
    .activate  (PE757_acount[7:0]               ), //i
    .weight    (PE658_bcount[7:0]               ), //i
    .valid     (PE758_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE758_acount[7:0]               ), //o
    .bcount    (PE758_bcount[7:0]               ), //o
    .PE_OUT    (PE758_PE_OUT[31:0]              ), //o
    .finish    (PE758_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE759 (
    .activate  (PE758_acount[7:0]               ), //i
    .weight    (PE659_bcount[7:0]               ), //i
    .valid     (PE759_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE759_acount[7:0]               ), //o
    .bcount    (PE759_bcount[7:0]               ), //o
    .PE_OUT    (PE759_PE_OUT[31:0]              ), //o
    .finish    (PE759_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE760 (
    .activate  (PE759_acount[7:0]               ), //i
    .weight    (PE660_bcount[7:0]               ), //i
    .valid     (PE760_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE760_acount[7:0]               ), //o
    .bcount    (PE760_bcount[7:0]               ), //o
    .PE_OUT    (PE760_PE_OUT[31:0]              ), //o
    .finish    (PE760_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE761 (
    .activate  (PE760_acount[7:0]               ), //i
    .weight    (PE661_bcount[7:0]               ), //i
    .valid     (PE761_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE761_acount[7:0]               ), //o
    .bcount    (PE761_bcount[7:0]               ), //o
    .PE_OUT    (PE761_PE_OUT[31:0]              ), //o
    .finish    (PE761_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE762 (
    .activate  (PE761_acount[7:0]               ), //i
    .weight    (PE662_bcount[7:0]               ), //i
    .valid     (PE762_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE762_acount[7:0]               ), //o
    .bcount    (PE762_bcount[7:0]               ), //o
    .PE_OUT    (PE762_PE_OUT[31:0]              ), //o
    .finish    (PE762_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  PE PE763 (
    .activate  (PE762_acount[7:0]               ), //i
    .weight    (PE663_bcount[7:0]               ), //i
    .valid     (PE763_valid                     ), //i
    .signCount (io_signCount_regNextWhen_7[15:0]), //i
    .acount    (PE763_acount[7:0]               ), //o
    .bcount    (PE763_bcount[7:0]               ), //o
    .PE_OUT    (PE763_PE_OUT[31:0]              ), //o
    .finish    (PE763_finish                    ), //o
    .clk       (clk                             ), //i
    .reset     (reset                           )  //i
  );
  always @(*) begin
    MatrixC_0 = 32'h0;
    if(PE00_finish) begin
      MatrixC_0 = PE00_PE_OUT;
    end
    if(PE01_finish) begin
      MatrixC_0 = PE01_PE_OUT;
    end
    if(PE02_finish) begin
      MatrixC_0 = PE02_PE_OUT;
    end
    if(PE03_finish) begin
      MatrixC_0 = PE03_PE_OUT;
    end
    if(PE04_finish) begin
      MatrixC_0 = PE04_PE_OUT;
    end
    if(PE05_finish) begin
      MatrixC_0 = PE05_PE_OUT;
    end
    if(PE06_finish) begin
      MatrixC_0 = PE06_PE_OUT;
    end
    if(PE07_finish) begin
      MatrixC_0 = PE07_PE_OUT;
    end
    if(PE08_finish) begin
      MatrixC_0 = PE08_PE_OUT;
    end
    if(PE09_finish) begin
      MatrixC_0 = PE09_PE_OUT;
    end
    if(PE010_finish) begin
      MatrixC_0 = PE010_PE_OUT;
    end
    if(PE011_finish) begin
      MatrixC_0 = PE011_PE_OUT;
    end
    if(PE012_finish) begin
      MatrixC_0 = PE012_PE_OUT;
    end
    if(PE013_finish) begin
      MatrixC_0 = PE013_PE_OUT;
    end
    if(PE014_finish) begin
      MatrixC_0 = PE014_PE_OUT;
    end
    if(PE015_finish) begin
      MatrixC_0 = PE015_PE_OUT;
    end
    if(PE016_finish) begin
      MatrixC_0 = PE016_PE_OUT;
    end
    if(PE017_finish) begin
      MatrixC_0 = PE017_PE_OUT;
    end
    if(PE018_finish) begin
      MatrixC_0 = PE018_PE_OUT;
    end
    if(PE019_finish) begin
      MatrixC_0 = PE019_PE_OUT;
    end
    if(PE020_finish) begin
      MatrixC_0 = PE020_PE_OUT;
    end
    if(PE021_finish) begin
      MatrixC_0 = PE021_PE_OUT;
    end
    if(PE022_finish) begin
      MatrixC_0 = PE022_PE_OUT;
    end
    if(PE023_finish) begin
      MatrixC_0 = PE023_PE_OUT;
    end
    if(PE024_finish) begin
      MatrixC_0 = PE024_PE_OUT;
    end
    if(PE025_finish) begin
      MatrixC_0 = PE025_PE_OUT;
    end
    if(PE026_finish) begin
      MatrixC_0 = PE026_PE_OUT;
    end
    if(PE027_finish) begin
      MatrixC_0 = PE027_PE_OUT;
    end
    if(PE028_finish) begin
      MatrixC_0 = PE028_PE_OUT;
    end
    if(PE029_finish) begin
      MatrixC_0 = PE029_PE_OUT;
    end
    if(PE030_finish) begin
      MatrixC_0 = PE030_PE_OUT;
    end
    if(PE031_finish) begin
      MatrixC_0 = PE031_PE_OUT;
    end
    if(PE032_finish) begin
      MatrixC_0 = PE032_PE_OUT;
    end
    if(PE033_finish) begin
      MatrixC_0 = PE033_PE_OUT;
    end
    if(PE034_finish) begin
      MatrixC_0 = PE034_PE_OUT;
    end
    if(PE035_finish) begin
      MatrixC_0 = PE035_PE_OUT;
    end
    if(PE036_finish) begin
      MatrixC_0 = PE036_PE_OUT;
    end
    if(PE037_finish) begin
      MatrixC_0 = PE037_PE_OUT;
    end
    if(PE038_finish) begin
      MatrixC_0 = PE038_PE_OUT;
    end
    if(PE039_finish) begin
      MatrixC_0 = PE039_PE_OUT;
    end
    if(PE040_finish) begin
      MatrixC_0 = PE040_PE_OUT;
    end
    if(PE041_finish) begin
      MatrixC_0 = PE041_PE_OUT;
    end
    if(PE042_finish) begin
      MatrixC_0 = PE042_PE_OUT;
    end
    if(PE043_finish) begin
      MatrixC_0 = PE043_PE_OUT;
    end
    if(PE044_finish) begin
      MatrixC_0 = PE044_PE_OUT;
    end
    if(PE045_finish) begin
      MatrixC_0 = PE045_PE_OUT;
    end
    if(PE046_finish) begin
      MatrixC_0 = PE046_PE_OUT;
    end
    if(PE047_finish) begin
      MatrixC_0 = PE047_PE_OUT;
    end
    if(PE048_finish) begin
      MatrixC_0 = PE048_PE_OUT;
    end
    if(PE049_finish) begin
      MatrixC_0 = PE049_PE_OUT;
    end
    if(PE050_finish) begin
      MatrixC_0 = PE050_PE_OUT;
    end
    if(PE051_finish) begin
      MatrixC_0 = PE051_PE_OUT;
    end
    if(PE052_finish) begin
      MatrixC_0 = PE052_PE_OUT;
    end
    if(PE053_finish) begin
      MatrixC_0 = PE053_PE_OUT;
    end
    if(PE054_finish) begin
      MatrixC_0 = PE054_PE_OUT;
    end
    if(PE055_finish) begin
      MatrixC_0 = PE055_PE_OUT;
    end
    if(PE056_finish) begin
      MatrixC_0 = PE056_PE_OUT;
    end
    if(PE057_finish) begin
      MatrixC_0 = PE057_PE_OUT;
    end
    if(PE058_finish) begin
      MatrixC_0 = PE058_PE_OUT;
    end
    if(PE059_finish) begin
      MatrixC_0 = PE059_PE_OUT;
    end
    if(PE060_finish) begin
      MatrixC_0 = PE060_PE_OUT;
    end
    if(PE061_finish) begin
      MatrixC_0 = PE061_PE_OUT;
    end
    if(PE062_finish) begin
      MatrixC_0 = PE062_PE_OUT;
    end
    if(PE063_finish) begin
      MatrixC_0 = PE063_PE_OUT;
    end
  end

  always @(*) begin
    _zz_C_Valid_0[0] = PE00_finish;
    _zz_C_Valid_0[1] = PE01_finish;
    _zz_C_Valid_0[2] = PE02_finish;
    _zz_C_Valid_0[3] = PE03_finish;
    _zz_C_Valid_0[4] = PE04_finish;
    _zz_C_Valid_0[5] = PE05_finish;
    _zz_C_Valid_0[6] = PE06_finish;
    _zz_C_Valid_0[7] = PE07_finish;
    _zz_C_Valid_0[8] = PE08_finish;
    _zz_C_Valid_0[9] = PE09_finish;
    _zz_C_Valid_0[10] = PE010_finish;
    _zz_C_Valid_0[11] = PE011_finish;
    _zz_C_Valid_0[12] = PE012_finish;
    _zz_C_Valid_0[13] = PE013_finish;
    _zz_C_Valid_0[14] = PE014_finish;
    _zz_C_Valid_0[15] = PE015_finish;
    _zz_C_Valid_0[16] = PE016_finish;
    _zz_C_Valid_0[17] = PE017_finish;
    _zz_C_Valid_0[18] = PE018_finish;
    _zz_C_Valid_0[19] = PE019_finish;
    _zz_C_Valid_0[20] = PE020_finish;
    _zz_C_Valid_0[21] = PE021_finish;
    _zz_C_Valid_0[22] = PE022_finish;
    _zz_C_Valid_0[23] = PE023_finish;
    _zz_C_Valid_0[24] = PE024_finish;
    _zz_C_Valid_0[25] = PE025_finish;
    _zz_C_Valid_0[26] = PE026_finish;
    _zz_C_Valid_0[27] = PE027_finish;
    _zz_C_Valid_0[28] = PE028_finish;
    _zz_C_Valid_0[29] = PE029_finish;
    _zz_C_Valid_0[30] = PE030_finish;
    _zz_C_Valid_0[31] = PE031_finish;
    _zz_C_Valid_0[32] = PE032_finish;
    _zz_C_Valid_0[33] = PE033_finish;
    _zz_C_Valid_0[34] = PE034_finish;
    _zz_C_Valid_0[35] = PE035_finish;
    _zz_C_Valid_0[36] = PE036_finish;
    _zz_C_Valid_0[37] = PE037_finish;
    _zz_C_Valid_0[38] = PE038_finish;
    _zz_C_Valid_0[39] = PE039_finish;
    _zz_C_Valid_0[40] = PE040_finish;
    _zz_C_Valid_0[41] = PE041_finish;
    _zz_C_Valid_0[42] = PE042_finish;
    _zz_C_Valid_0[43] = PE043_finish;
    _zz_C_Valid_0[44] = PE044_finish;
    _zz_C_Valid_0[45] = PE045_finish;
    _zz_C_Valid_0[46] = PE046_finish;
    _zz_C_Valid_0[47] = PE047_finish;
    _zz_C_Valid_0[48] = PE048_finish;
    _zz_C_Valid_0[49] = PE049_finish;
    _zz_C_Valid_0[50] = PE050_finish;
    _zz_C_Valid_0[51] = PE051_finish;
    _zz_C_Valid_0[52] = PE052_finish;
    _zz_C_Valid_0[53] = PE053_finish;
    _zz_C_Valid_0[54] = PE054_finish;
    _zz_C_Valid_0[55] = PE055_finish;
    _zz_C_Valid_0[56] = PE056_finish;
    _zz_C_Valid_0[57] = PE057_finish;
    _zz_C_Valid_0[58] = PE058_finish;
    _zz_C_Valid_0[59] = PE059_finish;
    _zz_C_Valid_0[60] = PE060_finish;
    _zz_C_Valid_0[61] = PE061_finish;
    _zz_C_Valid_0[62] = PE062_finish;
    _zz_C_Valid_0[63] = PE063_finish;
  end

  assign C_Valid_0 = (|_zz_C_Valid_0);
  always @(*) begin
    MatrixC_1 = 32'h0;
    if(PE10_finish) begin
      MatrixC_1 = PE10_PE_OUT;
    end
    if(PE11_finish) begin
      MatrixC_1 = PE11_PE_OUT;
    end
    if(PE12_finish) begin
      MatrixC_1 = PE12_PE_OUT;
    end
    if(PE13_finish) begin
      MatrixC_1 = PE13_PE_OUT;
    end
    if(PE14_finish) begin
      MatrixC_1 = PE14_PE_OUT;
    end
    if(PE15_finish) begin
      MatrixC_1 = PE15_PE_OUT;
    end
    if(PE16_finish) begin
      MatrixC_1 = PE16_PE_OUT;
    end
    if(PE17_finish) begin
      MatrixC_1 = PE17_PE_OUT;
    end
    if(PE18_finish) begin
      MatrixC_1 = PE18_PE_OUT;
    end
    if(PE19_finish) begin
      MatrixC_1 = PE19_PE_OUT;
    end
    if(PE110_finish) begin
      MatrixC_1 = PE110_PE_OUT;
    end
    if(PE111_finish) begin
      MatrixC_1 = PE111_PE_OUT;
    end
    if(PE112_finish) begin
      MatrixC_1 = PE112_PE_OUT;
    end
    if(PE113_finish) begin
      MatrixC_1 = PE113_PE_OUT;
    end
    if(PE114_finish) begin
      MatrixC_1 = PE114_PE_OUT;
    end
    if(PE115_finish) begin
      MatrixC_1 = PE115_PE_OUT;
    end
    if(PE116_finish) begin
      MatrixC_1 = PE116_PE_OUT;
    end
    if(PE117_finish) begin
      MatrixC_1 = PE117_PE_OUT;
    end
    if(PE118_finish) begin
      MatrixC_1 = PE118_PE_OUT;
    end
    if(PE119_finish) begin
      MatrixC_1 = PE119_PE_OUT;
    end
    if(PE120_finish) begin
      MatrixC_1 = PE120_PE_OUT;
    end
    if(PE121_finish) begin
      MatrixC_1 = PE121_PE_OUT;
    end
    if(PE122_finish) begin
      MatrixC_1 = PE122_PE_OUT;
    end
    if(PE123_finish) begin
      MatrixC_1 = PE123_PE_OUT;
    end
    if(PE124_finish) begin
      MatrixC_1 = PE124_PE_OUT;
    end
    if(PE125_finish) begin
      MatrixC_1 = PE125_PE_OUT;
    end
    if(PE126_finish) begin
      MatrixC_1 = PE126_PE_OUT;
    end
    if(PE127_finish) begin
      MatrixC_1 = PE127_PE_OUT;
    end
    if(PE128_finish) begin
      MatrixC_1 = PE128_PE_OUT;
    end
    if(PE129_finish) begin
      MatrixC_1 = PE129_PE_OUT;
    end
    if(PE130_finish) begin
      MatrixC_1 = PE130_PE_OUT;
    end
    if(PE131_finish) begin
      MatrixC_1 = PE131_PE_OUT;
    end
    if(PE132_finish) begin
      MatrixC_1 = PE132_PE_OUT;
    end
    if(PE133_finish) begin
      MatrixC_1 = PE133_PE_OUT;
    end
    if(PE134_finish) begin
      MatrixC_1 = PE134_PE_OUT;
    end
    if(PE135_finish) begin
      MatrixC_1 = PE135_PE_OUT;
    end
    if(PE136_finish) begin
      MatrixC_1 = PE136_PE_OUT;
    end
    if(PE137_finish) begin
      MatrixC_1 = PE137_PE_OUT;
    end
    if(PE138_finish) begin
      MatrixC_1 = PE138_PE_OUT;
    end
    if(PE139_finish) begin
      MatrixC_1 = PE139_PE_OUT;
    end
    if(PE140_finish) begin
      MatrixC_1 = PE140_PE_OUT;
    end
    if(PE141_finish) begin
      MatrixC_1 = PE141_PE_OUT;
    end
    if(PE142_finish) begin
      MatrixC_1 = PE142_PE_OUT;
    end
    if(PE143_finish) begin
      MatrixC_1 = PE143_PE_OUT;
    end
    if(PE144_finish) begin
      MatrixC_1 = PE144_PE_OUT;
    end
    if(PE145_finish) begin
      MatrixC_1 = PE145_PE_OUT;
    end
    if(PE146_finish) begin
      MatrixC_1 = PE146_PE_OUT;
    end
    if(PE147_finish) begin
      MatrixC_1 = PE147_PE_OUT;
    end
    if(PE148_finish) begin
      MatrixC_1 = PE148_PE_OUT;
    end
    if(PE149_finish) begin
      MatrixC_1 = PE149_PE_OUT;
    end
    if(PE150_finish) begin
      MatrixC_1 = PE150_PE_OUT;
    end
    if(PE151_finish) begin
      MatrixC_1 = PE151_PE_OUT;
    end
    if(PE152_finish) begin
      MatrixC_1 = PE152_PE_OUT;
    end
    if(PE153_finish) begin
      MatrixC_1 = PE153_PE_OUT;
    end
    if(PE154_finish) begin
      MatrixC_1 = PE154_PE_OUT;
    end
    if(PE155_finish) begin
      MatrixC_1 = PE155_PE_OUT;
    end
    if(PE156_finish) begin
      MatrixC_1 = PE156_PE_OUT;
    end
    if(PE157_finish) begin
      MatrixC_1 = PE157_PE_OUT;
    end
    if(PE158_finish) begin
      MatrixC_1 = PE158_PE_OUT;
    end
    if(PE159_finish) begin
      MatrixC_1 = PE159_PE_OUT;
    end
    if(PE160_finish) begin
      MatrixC_1 = PE160_PE_OUT;
    end
    if(PE161_finish) begin
      MatrixC_1 = PE161_PE_OUT;
    end
    if(PE162_finish) begin
      MatrixC_1 = PE162_PE_OUT;
    end
    if(PE163_finish) begin
      MatrixC_1 = PE163_PE_OUT;
    end
  end

  always @(*) begin
    _zz_C_Valid_1[0] = PE10_finish;
    _zz_C_Valid_1[1] = PE11_finish;
    _zz_C_Valid_1[2] = PE12_finish;
    _zz_C_Valid_1[3] = PE13_finish;
    _zz_C_Valid_1[4] = PE14_finish;
    _zz_C_Valid_1[5] = PE15_finish;
    _zz_C_Valid_1[6] = PE16_finish;
    _zz_C_Valid_1[7] = PE17_finish;
    _zz_C_Valid_1[8] = PE18_finish;
    _zz_C_Valid_1[9] = PE19_finish;
    _zz_C_Valid_1[10] = PE110_finish;
    _zz_C_Valid_1[11] = PE111_finish;
    _zz_C_Valid_1[12] = PE112_finish;
    _zz_C_Valid_1[13] = PE113_finish;
    _zz_C_Valid_1[14] = PE114_finish;
    _zz_C_Valid_1[15] = PE115_finish;
    _zz_C_Valid_1[16] = PE116_finish;
    _zz_C_Valid_1[17] = PE117_finish;
    _zz_C_Valid_1[18] = PE118_finish;
    _zz_C_Valid_1[19] = PE119_finish;
    _zz_C_Valid_1[20] = PE120_finish;
    _zz_C_Valid_1[21] = PE121_finish;
    _zz_C_Valid_1[22] = PE122_finish;
    _zz_C_Valid_1[23] = PE123_finish;
    _zz_C_Valid_1[24] = PE124_finish;
    _zz_C_Valid_1[25] = PE125_finish;
    _zz_C_Valid_1[26] = PE126_finish;
    _zz_C_Valid_1[27] = PE127_finish;
    _zz_C_Valid_1[28] = PE128_finish;
    _zz_C_Valid_1[29] = PE129_finish;
    _zz_C_Valid_1[30] = PE130_finish;
    _zz_C_Valid_1[31] = PE131_finish;
    _zz_C_Valid_1[32] = PE132_finish;
    _zz_C_Valid_1[33] = PE133_finish;
    _zz_C_Valid_1[34] = PE134_finish;
    _zz_C_Valid_1[35] = PE135_finish;
    _zz_C_Valid_1[36] = PE136_finish;
    _zz_C_Valid_1[37] = PE137_finish;
    _zz_C_Valid_1[38] = PE138_finish;
    _zz_C_Valid_1[39] = PE139_finish;
    _zz_C_Valid_1[40] = PE140_finish;
    _zz_C_Valid_1[41] = PE141_finish;
    _zz_C_Valid_1[42] = PE142_finish;
    _zz_C_Valid_1[43] = PE143_finish;
    _zz_C_Valid_1[44] = PE144_finish;
    _zz_C_Valid_1[45] = PE145_finish;
    _zz_C_Valid_1[46] = PE146_finish;
    _zz_C_Valid_1[47] = PE147_finish;
    _zz_C_Valid_1[48] = PE148_finish;
    _zz_C_Valid_1[49] = PE149_finish;
    _zz_C_Valid_1[50] = PE150_finish;
    _zz_C_Valid_1[51] = PE151_finish;
    _zz_C_Valid_1[52] = PE152_finish;
    _zz_C_Valid_1[53] = PE153_finish;
    _zz_C_Valid_1[54] = PE154_finish;
    _zz_C_Valid_1[55] = PE155_finish;
    _zz_C_Valid_1[56] = PE156_finish;
    _zz_C_Valid_1[57] = PE157_finish;
    _zz_C_Valid_1[58] = PE158_finish;
    _zz_C_Valid_1[59] = PE159_finish;
    _zz_C_Valid_1[60] = PE160_finish;
    _zz_C_Valid_1[61] = PE161_finish;
    _zz_C_Valid_1[62] = PE162_finish;
    _zz_C_Valid_1[63] = PE163_finish;
  end

  assign C_Valid_1 = (|_zz_C_Valid_1);
  always @(*) begin
    MatrixC_2 = 32'h0;
    if(PE20_finish) begin
      MatrixC_2 = PE20_PE_OUT;
    end
    if(PE21_finish) begin
      MatrixC_2 = PE21_PE_OUT;
    end
    if(PE22_finish) begin
      MatrixC_2 = PE22_PE_OUT;
    end
    if(PE23_finish) begin
      MatrixC_2 = PE23_PE_OUT;
    end
    if(PE24_finish) begin
      MatrixC_2 = PE24_PE_OUT;
    end
    if(PE25_finish) begin
      MatrixC_2 = PE25_PE_OUT;
    end
    if(PE26_finish) begin
      MatrixC_2 = PE26_PE_OUT;
    end
    if(PE27_finish) begin
      MatrixC_2 = PE27_PE_OUT;
    end
    if(PE28_finish) begin
      MatrixC_2 = PE28_PE_OUT;
    end
    if(PE29_finish) begin
      MatrixC_2 = PE29_PE_OUT;
    end
    if(PE210_finish) begin
      MatrixC_2 = PE210_PE_OUT;
    end
    if(PE211_finish) begin
      MatrixC_2 = PE211_PE_OUT;
    end
    if(PE212_finish) begin
      MatrixC_2 = PE212_PE_OUT;
    end
    if(PE213_finish) begin
      MatrixC_2 = PE213_PE_OUT;
    end
    if(PE214_finish) begin
      MatrixC_2 = PE214_PE_OUT;
    end
    if(PE215_finish) begin
      MatrixC_2 = PE215_PE_OUT;
    end
    if(PE216_finish) begin
      MatrixC_2 = PE216_PE_OUT;
    end
    if(PE217_finish) begin
      MatrixC_2 = PE217_PE_OUT;
    end
    if(PE218_finish) begin
      MatrixC_2 = PE218_PE_OUT;
    end
    if(PE219_finish) begin
      MatrixC_2 = PE219_PE_OUT;
    end
    if(PE220_finish) begin
      MatrixC_2 = PE220_PE_OUT;
    end
    if(PE221_finish) begin
      MatrixC_2 = PE221_PE_OUT;
    end
    if(PE222_finish) begin
      MatrixC_2 = PE222_PE_OUT;
    end
    if(PE223_finish) begin
      MatrixC_2 = PE223_PE_OUT;
    end
    if(PE224_finish) begin
      MatrixC_2 = PE224_PE_OUT;
    end
    if(PE225_finish) begin
      MatrixC_2 = PE225_PE_OUT;
    end
    if(PE226_finish) begin
      MatrixC_2 = PE226_PE_OUT;
    end
    if(PE227_finish) begin
      MatrixC_2 = PE227_PE_OUT;
    end
    if(PE228_finish) begin
      MatrixC_2 = PE228_PE_OUT;
    end
    if(PE229_finish) begin
      MatrixC_2 = PE229_PE_OUT;
    end
    if(PE230_finish) begin
      MatrixC_2 = PE230_PE_OUT;
    end
    if(PE231_finish) begin
      MatrixC_2 = PE231_PE_OUT;
    end
    if(PE232_finish) begin
      MatrixC_2 = PE232_PE_OUT;
    end
    if(PE233_finish) begin
      MatrixC_2 = PE233_PE_OUT;
    end
    if(PE234_finish) begin
      MatrixC_2 = PE234_PE_OUT;
    end
    if(PE235_finish) begin
      MatrixC_2 = PE235_PE_OUT;
    end
    if(PE236_finish) begin
      MatrixC_2 = PE236_PE_OUT;
    end
    if(PE237_finish) begin
      MatrixC_2 = PE237_PE_OUT;
    end
    if(PE238_finish) begin
      MatrixC_2 = PE238_PE_OUT;
    end
    if(PE239_finish) begin
      MatrixC_2 = PE239_PE_OUT;
    end
    if(PE240_finish) begin
      MatrixC_2 = PE240_PE_OUT;
    end
    if(PE241_finish) begin
      MatrixC_2 = PE241_PE_OUT;
    end
    if(PE242_finish) begin
      MatrixC_2 = PE242_PE_OUT;
    end
    if(PE243_finish) begin
      MatrixC_2 = PE243_PE_OUT;
    end
    if(PE244_finish) begin
      MatrixC_2 = PE244_PE_OUT;
    end
    if(PE245_finish) begin
      MatrixC_2 = PE245_PE_OUT;
    end
    if(PE246_finish) begin
      MatrixC_2 = PE246_PE_OUT;
    end
    if(PE247_finish) begin
      MatrixC_2 = PE247_PE_OUT;
    end
    if(PE248_finish) begin
      MatrixC_2 = PE248_PE_OUT;
    end
    if(PE249_finish) begin
      MatrixC_2 = PE249_PE_OUT;
    end
    if(PE250_finish) begin
      MatrixC_2 = PE250_PE_OUT;
    end
    if(PE251_finish) begin
      MatrixC_2 = PE251_PE_OUT;
    end
    if(PE252_finish) begin
      MatrixC_2 = PE252_PE_OUT;
    end
    if(PE253_finish) begin
      MatrixC_2 = PE253_PE_OUT;
    end
    if(PE254_finish) begin
      MatrixC_2 = PE254_PE_OUT;
    end
    if(PE255_finish) begin
      MatrixC_2 = PE255_PE_OUT;
    end
    if(PE256_finish) begin
      MatrixC_2 = PE256_PE_OUT;
    end
    if(PE257_finish) begin
      MatrixC_2 = PE257_PE_OUT;
    end
    if(PE258_finish) begin
      MatrixC_2 = PE258_PE_OUT;
    end
    if(PE259_finish) begin
      MatrixC_2 = PE259_PE_OUT;
    end
    if(PE260_finish) begin
      MatrixC_2 = PE260_PE_OUT;
    end
    if(PE261_finish) begin
      MatrixC_2 = PE261_PE_OUT;
    end
    if(PE262_finish) begin
      MatrixC_2 = PE262_PE_OUT;
    end
    if(PE263_finish) begin
      MatrixC_2 = PE263_PE_OUT;
    end
  end

  always @(*) begin
    _zz_C_Valid_2[0] = PE20_finish;
    _zz_C_Valid_2[1] = PE21_finish;
    _zz_C_Valid_2[2] = PE22_finish;
    _zz_C_Valid_2[3] = PE23_finish;
    _zz_C_Valid_2[4] = PE24_finish;
    _zz_C_Valid_2[5] = PE25_finish;
    _zz_C_Valid_2[6] = PE26_finish;
    _zz_C_Valid_2[7] = PE27_finish;
    _zz_C_Valid_2[8] = PE28_finish;
    _zz_C_Valid_2[9] = PE29_finish;
    _zz_C_Valid_2[10] = PE210_finish;
    _zz_C_Valid_2[11] = PE211_finish;
    _zz_C_Valid_2[12] = PE212_finish;
    _zz_C_Valid_2[13] = PE213_finish;
    _zz_C_Valid_2[14] = PE214_finish;
    _zz_C_Valid_2[15] = PE215_finish;
    _zz_C_Valid_2[16] = PE216_finish;
    _zz_C_Valid_2[17] = PE217_finish;
    _zz_C_Valid_2[18] = PE218_finish;
    _zz_C_Valid_2[19] = PE219_finish;
    _zz_C_Valid_2[20] = PE220_finish;
    _zz_C_Valid_2[21] = PE221_finish;
    _zz_C_Valid_2[22] = PE222_finish;
    _zz_C_Valid_2[23] = PE223_finish;
    _zz_C_Valid_2[24] = PE224_finish;
    _zz_C_Valid_2[25] = PE225_finish;
    _zz_C_Valid_2[26] = PE226_finish;
    _zz_C_Valid_2[27] = PE227_finish;
    _zz_C_Valid_2[28] = PE228_finish;
    _zz_C_Valid_2[29] = PE229_finish;
    _zz_C_Valid_2[30] = PE230_finish;
    _zz_C_Valid_2[31] = PE231_finish;
    _zz_C_Valid_2[32] = PE232_finish;
    _zz_C_Valid_2[33] = PE233_finish;
    _zz_C_Valid_2[34] = PE234_finish;
    _zz_C_Valid_2[35] = PE235_finish;
    _zz_C_Valid_2[36] = PE236_finish;
    _zz_C_Valid_2[37] = PE237_finish;
    _zz_C_Valid_2[38] = PE238_finish;
    _zz_C_Valid_2[39] = PE239_finish;
    _zz_C_Valid_2[40] = PE240_finish;
    _zz_C_Valid_2[41] = PE241_finish;
    _zz_C_Valid_2[42] = PE242_finish;
    _zz_C_Valid_2[43] = PE243_finish;
    _zz_C_Valid_2[44] = PE244_finish;
    _zz_C_Valid_2[45] = PE245_finish;
    _zz_C_Valid_2[46] = PE246_finish;
    _zz_C_Valid_2[47] = PE247_finish;
    _zz_C_Valid_2[48] = PE248_finish;
    _zz_C_Valid_2[49] = PE249_finish;
    _zz_C_Valid_2[50] = PE250_finish;
    _zz_C_Valid_2[51] = PE251_finish;
    _zz_C_Valid_2[52] = PE252_finish;
    _zz_C_Valid_2[53] = PE253_finish;
    _zz_C_Valid_2[54] = PE254_finish;
    _zz_C_Valid_2[55] = PE255_finish;
    _zz_C_Valid_2[56] = PE256_finish;
    _zz_C_Valid_2[57] = PE257_finish;
    _zz_C_Valid_2[58] = PE258_finish;
    _zz_C_Valid_2[59] = PE259_finish;
    _zz_C_Valid_2[60] = PE260_finish;
    _zz_C_Valid_2[61] = PE261_finish;
    _zz_C_Valid_2[62] = PE262_finish;
    _zz_C_Valid_2[63] = PE263_finish;
  end

  assign C_Valid_2 = (|_zz_C_Valid_2);
  always @(*) begin
    MatrixC_3 = 32'h0;
    if(PE30_finish) begin
      MatrixC_3 = PE30_PE_OUT;
    end
    if(PE31_finish) begin
      MatrixC_3 = PE31_PE_OUT;
    end
    if(PE32_finish) begin
      MatrixC_3 = PE32_PE_OUT;
    end
    if(PE33_finish) begin
      MatrixC_3 = PE33_PE_OUT;
    end
    if(PE34_finish) begin
      MatrixC_3 = PE34_PE_OUT;
    end
    if(PE35_finish) begin
      MatrixC_3 = PE35_PE_OUT;
    end
    if(PE36_finish) begin
      MatrixC_3 = PE36_PE_OUT;
    end
    if(PE37_finish) begin
      MatrixC_3 = PE37_PE_OUT;
    end
    if(PE38_finish) begin
      MatrixC_3 = PE38_PE_OUT;
    end
    if(PE39_finish) begin
      MatrixC_3 = PE39_PE_OUT;
    end
    if(PE310_finish) begin
      MatrixC_3 = PE310_PE_OUT;
    end
    if(PE311_finish) begin
      MatrixC_3 = PE311_PE_OUT;
    end
    if(PE312_finish) begin
      MatrixC_3 = PE312_PE_OUT;
    end
    if(PE313_finish) begin
      MatrixC_3 = PE313_PE_OUT;
    end
    if(PE314_finish) begin
      MatrixC_3 = PE314_PE_OUT;
    end
    if(PE315_finish) begin
      MatrixC_3 = PE315_PE_OUT;
    end
    if(PE316_finish) begin
      MatrixC_3 = PE316_PE_OUT;
    end
    if(PE317_finish) begin
      MatrixC_3 = PE317_PE_OUT;
    end
    if(PE318_finish) begin
      MatrixC_3 = PE318_PE_OUT;
    end
    if(PE319_finish) begin
      MatrixC_3 = PE319_PE_OUT;
    end
    if(PE320_finish) begin
      MatrixC_3 = PE320_PE_OUT;
    end
    if(PE321_finish) begin
      MatrixC_3 = PE321_PE_OUT;
    end
    if(PE322_finish) begin
      MatrixC_3 = PE322_PE_OUT;
    end
    if(PE323_finish) begin
      MatrixC_3 = PE323_PE_OUT;
    end
    if(PE324_finish) begin
      MatrixC_3 = PE324_PE_OUT;
    end
    if(PE325_finish) begin
      MatrixC_3 = PE325_PE_OUT;
    end
    if(PE326_finish) begin
      MatrixC_3 = PE326_PE_OUT;
    end
    if(PE327_finish) begin
      MatrixC_3 = PE327_PE_OUT;
    end
    if(PE328_finish) begin
      MatrixC_3 = PE328_PE_OUT;
    end
    if(PE329_finish) begin
      MatrixC_3 = PE329_PE_OUT;
    end
    if(PE330_finish) begin
      MatrixC_3 = PE330_PE_OUT;
    end
    if(PE331_finish) begin
      MatrixC_3 = PE331_PE_OUT;
    end
    if(PE332_finish) begin
      MatrixC_3 = PE332_PE_OUT;
    end
    if(PE333_finish) begin
      MatrixC_3 = PE333_PE_OUT;
    end
    if(PE334_finish) begin
      MatrixC_3 = PE334_PE_OUT;
    end
    if(PE335_finish) begin
      MatrixC_3 = PE335_PE_OUT;
    end
    if(PE336_finish) begin
      MatrixC_3 = PE336_PE_OUT;
    end
    if(PE337_finish) begin
      MatrixC_3 = PE337_PE_OUT;
    end
    if(PE338_finish) begin
      MatrixC_3 = PE338_PE_OUT;
    end
    if(PE339_finish) begin
      MatrixC_3 = PE339_PE_OUT;
    end
    if(PE340_finish) begin
      MatrixC_3 = PE340_PE_OUT;
    end
    if(PE341_finish) begin
      MatrixC_3 = PE341_PE_OUT;
    end
    if(PE342_finish) begin
      MatrixC_3 = PE342_PE_OUT;
    end
    if(PE343_finish) begin
      MatrixC_3 = PE343_PE_OUT;
    end
    if(PE344_finish) begin
      MatrixC_3 = PE344_PE_OUT;
    end
    if(PE345_finish) begin
      MatrixC_3 = PE345_PE_OUT;
    end
    if(PE346_finish) begin
      MatrixC_3 = PE346_PE_OUT;
    end
    if(PE347_finish) begin
      MatrixC_3 = PE347_PE_OUT;
    end
    if(PE348_finish) begin
      MatrixC_3 = PE348_PE_OUT;
    end
    if(PE349_finish) begin
      MatrixC_3 = PE349_PE_OUT;
    end
    if(PE350_finish) begin
      MatrixC_3 = PE350_PE_OUT;
    end
    if(PE351_finish) begin
      MatrixC_3 = PE351_PE_OUT;
    end
    if(PE352_finish) begin
      MatrixC_3 = PE352_PE_OUT;
    end
    if(PE353_finish) begin
      MatrixC_3 = PE353_PE_OUT;
    end
    if(PE354_finish) begin
      MatrixC_3 = PE354_PE_OUT;
    end
    if(PE355_finish) begin
      MatrixC_3 = PE355_PE_OUT;
    end
    if(PE356_finish) begin
      MatrixC_3 = PE356_PE_OUT;
    end
    if(PE357_finish) begin
      MatrixC_3 = PE357_PE_OUT;
    end
    if(PE358_finish) begin
      MatrixC_3 = PE358_PE_OUT;
    end
    if(PE359_finish) begin
      MatrixC_3 = PE359_PE_OUT;
    end
    if(PE360_finish) begin
      MatrixC_3 = PE360_PE_OUT;
    end
    if(PE361_finish) begin
      MatrixC_3 = PE361_PE_OUT;
    end
    if(PE362_finish) begin
      MatrixC_3 = PE362_PE_OUT;
    end
    if(PE363_finish) begin
      MatrixC_3 = PE363_PE_OUT;
    end
  end

  always @(*) begin
    _zz_C_Valid_3[0] = PE30_finish;
    _zz_C_Valid_3[1] = PE31_finish;
    _zz_C_Valid_3[2] = PE32_finish;
    _zz_C_Valid_3[3] = PE33_finish;
    _zz_C_Valid_3[4] = PE34_finish;
    _zz_C_Valid_3[5] = PE35_finish;
    _zz_C_Valid_3[6] = PE36_finish;
    _zz_C_Valid_3[7] = PE37_finish;
    _zz_C_Valid_3[8] = PE38_finish;
    _zz_C_Valid_3[9] = PE39_finish;
    _zz_C_Valid_3[10] = PE310_finish;
    _zz_C_Valid_3[11] = PE311_finish;
    _zz_C_Valid_3[12] = PE312_finish;
    _zz_C_Valid_3[13] = PE313_finish;
    _zz_C_Valid_3[14] = PE314_finish;
    _zz_C_Valid_3[15] = PE315_finish;
    _zz_C_Valid_3[16] = PE316_finish;
    _zz_C_Valid_3[17] = PE317_finish;
    _zz_C_Valid_3[18] = PE318_finish;
    _zz_C_Valid_3[19] = PE319_finish;
    _zz_C_Valid_3[20] = PE320_finish;
    _zz_C_Valid_3[21] = PE321_finish;
    _zz_C_Valid_3[22] = PE322_finish;
    _zz_C_Valid_3[23] = PE323_finish;
    _zz_C_Valid_3[24] = PE324_finish;
    _zz_C_Valid_3[25] = PE325_finish;
    _zz_C_Valid_3[26] = PE326_finish;
    _zz_C_Valid_3[27] = PE327_finish;
    _zz_C_Valid_3[28] = PE328_finish;
    _zz_C_Valid_3[29] = PE329_finish;
    _zz_C_Valid_3[30] = PE330_finish;
    _zz_C_Valid_3[31] = PE331_finish;
    _zz_C_Valid_3[32] = PE332_finish;
    _zz_C_Valid_3[33] = PE333_finish;
    _zz_C_Valid_3[34] = PE334_finish;
    _zz_C_Valid_3[35] = PE335_finish;
    _zz_C_Valid_3[36] = PE336_finish;
    _zz_C_Valid_3[37] = PE337_finish;
    _zz_C_Valid_3[38] = PE338_finish;
    _zz_C_Valid_3[39] = PE339_finish;
    _zz_C_Valid_3[40] = PE340_finish;
    _zz_C_Valid_3[41] = PE341_finish;
    _zz_C_Valid_3[42] = PE342_finish;
    _zz_C_Valid_3[43] = PE343_finish;
    _zz_C_Valid_3[44] = PE344_finish;
    _zz_C_Valid_3[45] = PE345_finish;
    _zz_C_Valid_3[46] = PE346_finish;
    _zz_C_Valid_3[47] = PE347_finish;
    _zz_C_Valid_3[48] = PE348_finish;
    _zz_C_Valid_3[49] = PE349_finish;
    _zz_C_Valid_3[50] = PE350_finish;
    _zz_C_Valid_3[51] = PE351_finish;
    _zz_C_Valid_3[52] = PE352_finish;
    _zz_C_Valid_3[53] = PE353_finish;
    _zz_C_Valid_3[54] = PE354_finish;
    _zz_C_Valid_3[55] = PE355_finish;
    _zz_C_Valid_3[56] = PE356_finish;
    _zz_C_Valid_3[57] = PE357_finish;
    _zz_C_Valid_3[58] = PE358_finish;
    _zz_C_Valid_3[59] = PE359_finish;
    _zz_C_Valid_3[60] = PE360_finish;
    _zz_C_Valid_3[61] = PE361_finish;
    _zz_C_Valid_3[62] = PE362_finish;
    _zz_C_Valid_3[63] = PE363_finish;
  end

  assign C_Valid_3 = (|_zz_C_Valid_3);
  always @(*) begin
    MatrixC_4 = 32'h0;
    if(PE40_finish) begin
      MatrixC_4 = PE40_PE_OUT;
    end
    if(PE41_finish) begin
      MatrixC_4 = PE41_PE_OUT;
    end
    if(PE42_finish) begin
      MatrixC_4 = PE42_PE_OUT;
    end
    if(PE43_finish) begin
      MatrixC_4 = PE43_PE_OUT;
    end
    if(PE44_finish) begin
      MatrixC_4 = PE44_PE_OUT;
    end
    if(PE45_finish) begin
      MatrixC_4 = PE45_PE_OUT;
    end
    if(PE46_finish) begin
      MatrixC_4 = PE46_PE_OUT;
    end
    if(PE47_finish) begin
      MatrixC_4 = PE47_PE_OUT;
    end
    if(PE48_finish) begin
      MatrixC_4 = PE48_PE_OUT;
    end
    if(PE49_finish) begin
      MatrixC_4 = PE49_PE_OUT;
    end
    if(PE410_finish) begin
      MatrixC_4 = PE410_PE_OUT;
    end
    if(PE411_finish) begin
      MatrixC_4 = PE411_PE_OUT;
    end
    if(PE412_finish) begin
      MatrixC_4 = PE412_PE_OUT;
    end
    if(PE413_finish) begin
      MatrixC_4 = PE413_PE_OUT;
    end
    if(PE414_finish) begin
      MatrixC_4 = PE414_PE_OUT;
    end
    if(PE415_finish) begin
      MatrixC_4 = PE415_PE_OUT;
    end
    if(PE416_finish) begin
      MatrixC_4 = PE416_PE_OUT;
    end
    if(PE417_finish) begin
      MatrixC_4 = PE417_PE_OUT;
    end
    if(PE418_finish) begin
      MatrixC_4 = PE418_PE_OUT;
    end
    if(PE419_finish) begin
      MatrixC_4 = PE419_PE_OUT;
    end
    if(PE420_finish) begin
      MatrixC_4 = PE420_PE_OUT;
    end
    if(PE421_finish) begin
      MatrixC_4 = PE421_PE_OUT;
    end
    if(PE422_finish) begin
      MatrixC_4 = PE422_PE_OUT;
    end
    if(PE423_finish) begin
      MatrixC_4 = PE423_PE_OUT;
    end
    if(PE424_finish) begin
      MatrixC_4 = PE424_PE_OUT;
    end
    if(PE425_finish) begin
      MatrixC_4 = PE425_PE_OUT;
    end
    if(PE426_finish) begin
      MatrixC_4 = PE426_PE_OUT;
    end
    if(PE427_finish) begin
      MatrixC_4 = PE427_PE_OUT;
    end
    if(PE428_finish) begin
      MatrixC_4 = PE428_PE_OUT;
    end
    if(PE429_finish) begin
      MatrixC_4 = PE429_PE_OUT;
    end
    if(PE430_finish) begin
      MatrixC_4 = PE430_PE_OUT;
    end
    if(PE431_finish) begin
      MatrixC_4 = PE431_PE_OUT;
    end
    if(PE432_finish) begin
      MatrixC_4 = PE432_PE_OUT;
    end
    if(PE433_finish) begin
      MatrixC_4 = PE433_PE_OUT;
    end
    if(PE434_finish) begin
      MatrixC_4 = PE434_PE_OUT;
    end
    if(PE435_finish) begin
      MatrixC_4 = PE435_PE_OUT;
    end
    if(PE436_finish) begin
      MatrixC_4 = PE436_PE_OUT;
    end
    if(PE437_finish) begin
      MatrixC_4 = PE437_PE_OUT;
    end
    if(PE438_finish) begin
      MatrixC_4 = PE438_PE_OUT;
    end
    if(PE439_finish) begin
      MatrixC_4 = PE439_PE_OUT;
    end
    if(PE440_finish) begin
      MatrixC_4 = PE440_PE_OUT;
    end
    if(PE441_finish) begin
      MatrixC_4 = PE441_PE_OUT;
    end
    if(PE442_finish) begin
      MatrixC_4 = PE442_PE_OUT;
    end
    if(PE443_finish) begin
      MatrixC_4 = PE443_PE_OUT;
    end
    if(PE444_finish) begin
      MatrixC_4 = PE444_PE_OUT;
    end
    if(PE445_finish) begin
      MatrixC_4 = PE445_PE_OUT;
    end
    if(PE446_finish) begin
      MatrixC_4 = PE446_PE_OUT;
    end
    if(PE447_finish) begin
      MatrixC_4 = PE447_PE_OUT;
    end
    if(PE448_finish) begin
      MatrixC_4 = PE448_PE_OUT;
    end
    if(PE449_finish) begin
      MatrixC_4 = PE449_PE_OUT;
    end
    if(PE450_finish) begin
      MatrixC_4 = PE450_PE_OUT;
    end
    if(PE451_finish) begin
      MatrixC_4 = PE451_PE_OUT;
    end
    if(PE452_finish) begin
      MatrixC_4 = PE452_PE_OUT;
    end
    if(PE453_finish) begin
      MatrixC_4 = PE453_PE_OUT;
    end
    if(PE454_finish) begin
      MatrixC_4 = PE454_PE_OUT;
    end
    if(PE455_finish) begin
      MatrixC_4 = PE455_PE_OUT;
    end
    if(PE456_finish) begin
      MatrixC_4 = PE456_PE_OUT;
    end
    if(PE457_finish) begin
      MatrixC_4 = PE457_PE_OUT;
    end
    if(PE458_finish) begin
      MatrixC_4 = PE458_PE_OUT;
    end
    if(PE459_finish) begin
      MatrixC_4 = PE459_PE_OUT;
    end
    if(PE460_finish) begin
      MatrixC_4 = PE460_PE_OUT;
    end
    if(PE461_finish) begin
      MatrixC_4 = PE461_PE_OUT;
    end
    if(PE462_finish) begin
      MatrixC_4 = PE462_PE_OUT;
    end
    if(PE463_finish) begin
      MatrixC_4 = PE463_PE_OUT;
    end
  end

  always @(*) begin
    _zz_C_Valid_4[0] = PE40_finish;
    _zz_C_Valid_4[1] = PE41_finish;
    _zz_C_Valid_4[2] = PE42_finish;
    _zz_C_Valid_4[3] = PE43_finish;
    _zz_C_Valid_4[4] = PE44_finish;
    _zz_C_Valid_4[5] = PE45_finish;
    _zz_C_Valid_4[6] = PE46_finish;
    _zz_C_Valid_4[7] = PE47_finish;
    _zz_C_Valid_4[8] = PE48_finish;
    _zz_C_Valid_4[9] = PE49_finish;
    _zz_C_Valid_4[10] = PE410_finish;
    _zz_C_Valid_4[11] = PE411_finish;
    _zz_C_Valid_4[12] = PE412_finish;
    _zz_C_Valid_4[13] = PE413_finish;
    _zz_C_Valid_4[14] = PE414_finish;
    _zz_C_Valid_4[15] = PE415_finish;
    _zz_C_Valid_4[16] = PE416_finish;
    _zz_C_Valid_4[17] = PE417_finish;
    _zz_C_Valid_4[18] = PE418_finish;
    _zz_C_Valid_4[19] = PE419_finish;
    _zz_C_Valid_4[20] = PE420_finish;
    _zz_C_Valid_4[21] = PE421_finish;
    _zz_C_Valid_4[22] = PE422_finish;
    _zz_C_Valid_4[23] = PE423_finish;
    _zz_C_Valid_4[24] = PE424_finish;
    _zz_C_Valid_4[25] = PE425_finish;
    _zz_C_Valid_4[26] = PE426_finish;
    _zz_C_Valid_4[27] = PE427_finish;
    _zz_C_Valid_4[28] = PE428_finish;
    _zz_C_Valid_4[29] = PE429_finish;
    _zz_C_Valid_4[30] = PE430_finish;
    _zz_C_Valid_4[31] = PE431_finish;
    _zz_C_Valid_4[32] = PE432_finish;
    _zz_C_Valid_4[33] = PE433_finish;
    _zz_C_Valid_4[34] = PE434_finish;
    _zz_C_Valid_4[35] = PE435_finish;
    _zz_C_Valid_4[36] = PE436_finish;
    _zz_C_Valid_4[37] = PE437_finish;
    _zz_C_Valid_4[38] = PE438_finish;
    _zz_C_Valid_4[39] = PE439_finish;
    _zz_C_Valid_4[40] = PE440_finish;
    _zz_C_Valid_4[41] = PE441_finish;
    _zz_C_Valid_4[42] = PE442_finish;
    _zz_C_Valid_4[43] = PE443_finish;
    _zz_C_Valid_4[44] = PE444_finish;
    _zz_C_Valid_4[45] = PE445_finish;
    _zz_C_Valid_4[46] = PE446_finish;
    _zz_C_Valid_4[47] = PE447_finish;
    _zz_C_Valid_4[48] = PE448_finish;
    _zz_C_Valid_4[49] = PE449_finish;
    _zz_C_Valid_4[50] = PE450_finish;
    _zz_C_Valid_4[51] = PE451_finish;
    _zz_C_Valid_4[52] = PE452_finish;
    _zz_C_Valid_4[53] = PE453_finish;
    _zz_C_Valid_4[54] = PE454_finish;
    _zz_C_Valid_4[55] = PE455_finish;
    _zz_C_Valid_4[56] = PE456_finish;
    _zz_C_Valid_4[57] = PE457_finish;
    _zz_C_Valid_4[58] = PE458_finish;
    _zz_C_Valid_4[59] = PE459_finish;
    _zz_C_Valid_4[60] = PE460_finish;
    _zz_C_Valid_4[61] = PE461_finish;
    _zz_C_Valid_4[62] = PE462_finish;
    _zz_C_Valid_4[63] = PE463_finish;
  end

  assign C_Valid_4 = (|_zz_C_Valid_4);
  always @(*) begin
    MatrixC_5 = 32'h0;
    if(PE50_finish) begin
      MatrixC_5 = PE50_PE_OUT;
    end
    if(PE51_finish) begin
      MatrixC_5 = PE51_PE_OUT;
    end
    if(PE52_finish) begin
      MatrixC_5 = PE52_PE_OUT;
    end
    if(PE53_finish) begin
      MatrixC_5 = PE53_PE_OUT;
    end
    if(PE54_finish) begin
      MatrixC_5 = PE54_PE_OUT;
    end
    if(PE55_finish) begin
      MatrixC_5 = PE55_PE_OUT;
    end
    if(PE56_finish) begin
      MatrixC_5 = PE56_PE_OUT;
    end
    if(PE57_finish) begin
      MatrixC_5 = PE57_PE_OUT;
    end
    if(PE58_finish) begin
      MatrixC_5 = PE58_PE_OUT;
    end
    if(PE59_finish) begin
      MatrixC_5 = PE59_PE_OUT;
    end
    if(PE510_finish) begin
      MatrixC_5 = PE510_PE_OUT;
    end
    if(PE511_finish) begin
      MatrixC_5 = PE511_PE_OUT;
    end
    if(PE512_finish) begin
      MatrixC_5 = PE512_PE_OUT;
    end
    if(PE513_finish) begin
      MatrixC_5 = PE513_PE_OUT;
    end
    if(PE514_finish) begin
      MatrixC_5 = PE514_PE_OUT;
    end
    if(PE515_finish) begin
      MatrixC_5 = PE515_PE_OUT;
    end
    if(PE516_finish) begin
      MatrixC_5 = PE516_PE_OUT;
    end
    if(PE517_finish) begin
      MatrixC_5 = PE517_PE_OUT;
    end
    if(PE518_finish) begin
      MatrixC_5 = PE518_PE_OUT;
    end
    if(PE519_finish) begin
      MatrixC_5 = PE519_PE_OUT;
    end
    if(PE520_finish) begin
      MatrixC_5 = PE520_PE_OUT;
    end
    if(PE521_finish) begin
      MatrixC_5 = PE521_PE_OUT;
    end
    if(PE522_finish) begin
      MatrixC_5 = PE522_PE_OUT;
    end
    if(PE523_finish) begin
      MatrixC_5 = PE523_PE_OUT;
    end
    if(PE524_finish) begin
      MatrixC_5 = PE524_PE_OUT;
    end
    if(PE525_finish) begin
      MatrixC_5 = PE525_PE_OUT;
    end
    if(PE526_finish) begin
      MatrixC_5 = PE526_PE_OUT;
    end
    if(PE527_finish) begin
      MatrixC_5 = PE527_PE_OUT;
    end
    if(PE528_finish) begin
      MatrixC_5 = PE528_PE_OUT;
    end
    if(PE529_finish) begin
      MatrixC_5 = PE529_PE_OUT;
    end
    if(PE530_finish) begin
      MatrixC_5 = PE530_PE_OUT;
    end
    if(PE531_finish) begin
      MatrixC_5 = PE531_PE_OUT;
    end
    if(PE532_finish) begin
      MatrixC_5 = PE532_PE_OUT;
    end
    if(PE533_finish) begin
      MatrixC_5 = PE533_PE_OUT;
    end
    if(PE534_finish) begin
      MatrixC_5 = PE534_PE_OUT;
    end
    if(PE535_finish) begin
      MatrixC_5 = PE535_PE_OUT;
    end
    if(PE536_finish) begin
      MatrixC_5 = PE536_PE_OUT;
    end
    if(PE537_finish) begin
      MatrixC_5 = PE537_PE_OUT;
    end
    if(PE538_finish) begin
      MatrixC_5 = PE538_PE_OUT;
    end
    if(PE539_finish) begin
      MatrixC_5 = PE539_PE_OUT;
    end
    if(PE540_finish) begin
      MatrixC_5 = PE540_PE_OUT;
    end
    if(PE541_finish) begin
      MatrixC_5 = PE541_PE_OUT;
    end
    if(PE542_finish) begin
      MatrixC_5 = PE542_PE_OUT;
    end
    if(PE543_finish) begin
      MatrixC_5 = PE543_PE_OUT;
    end
    if(PE544_finish) begin
      MatrixC_5 = PE544_PE_OUT;
    end
    if(PE545_finish) begin
      MatrixC_5 = PE545_PE_OUT;
    end
    if(PE546_finish) begin
      MatrixC_5 = PE546_PE_OUT;
    end
    if(PE547_finish) begin
      MatrixC_5 = PE547_PE_OUT;
    end
    if(PE548_finish) begin
      MatrixC_5 = PE548_PE_OUT;
    end
    if(PE549_finish) begin
      MatrixC_5 = PE549_PE_OUT;
    end
    if(PE550_finish) begin
      MatrixC_5 = PE550_PE_OUT;
    end
    if(PE551_finish) begin
      MatrixC_5 = PE551_PE_OUT;
    end
    if(PE552_finish) begin
      MatrixC_5 = PE552_PE_OUT;
    end
    if(PE553_finish) begin
      MatrixC_5 = PE553_PE_OUT;
    end
    if(PE554_finish) begin
      MatrixC_5 = PE554_PE_OUT;
    end
    if(PE555_finish) begin
      MatrixC_5 = PE555_PE_OUT;
    end
    if(PE556_finish) begin
      MatrixC_5 = PE556_PE_OUT;
    end
    if(PE557_finish) begin
      MatrixC_5 = PE557_PE_OUT;
    end
    if(PE558_finish) begin
      MatrixC_5 = PE558_PE_OUT;
    end
    if(PE559_finish) begin
      MatrixC_5 = PE559_PE_OUT;
    end
    if(PE560_finish) begin
      MatrixC_5 = PE560_PE_OUT;
    end
    if(PE561_finish) begin
      MatrixC_5 = PE561_PE_OUT;
    end
    if(PE562_finish) begin
      MatrixC_5 = PE562_PE_OUT;
    end
    if(PE563_finish) begin
      MatrixC_5 = PE563_PE_OUT;
    end
  end

  always @(*) begin
    _zz_C_Valid_5[0] = PE50_finish;
    _zz_C_Valid_5[1] = PE51_finish;
    _zz_C_Valid_5[2] = PE52_finish;
    _zz_C_Valid_5[3] = PE53_finish;
    _zz_C_Valid_5[4] = PE54_finish;
    _zz_C_Valid_5[5] = PE55_finish;
    _zz_C_Valid_5[6] = PE56_finish;
    _zz_C_Valid_5[7] = PE57_finish;
    _zz_C_Valid_5[8] = PE58_finish;
    _zz_C_Valid_5[9] = PE59_finish;
    _zz_C_Valid_5[10] = PE510_finish;
    _zz_C_Valid_5[11] = PE511_finish;
    _zz_C_Valid_5[12] = PE512_finish;
    _zz_C_Valid_5[13] = PE513_finish;
    _zz_C_Valid_5[14] = PE514_finish;
    _zz_C_Valid_5[15] = PE515_finish;
    _zz_C_Valid_5[16] = PE516_finish;
    _zz_C_Valid_5[17] = PE517_finish;
    _zz_C_Valid_5[18] = PE518_finish;
    _zz_C_Valid_5[19] = PE519_finish;
    _zz_C_Valid_5[20] = PE520_finish;
    _zz_C_Valid_5[21] = PE521_finish;
    _zz_C_Valid_5[22] = PE522_finish;
    _zz_C_Valid_5[23] = PE523_finish;
    _zz_C_Valid_5[24] = PE524_finish;
    _zz_C_Valid_5[25] = PE525_finish;
    _zz_C_Valid_5[26] = PE526_finish;
    _zz_C_Valid_5[27] = PE527_finish;
    _zz_C_Valid_5[28] = PE528_finish;
    _zz_C_Valid_5[29] = PE529_finish;
    _zz_C_Valid_5[30] = PE530_finish;
    _zz_C_Valid_5[31] = PE531_finish;
    _zz_C_Valid_5[32] = PE532_finish;
    _zz_C_Valid_5[33] = PE533_finish;
    _zz_C_Valid_5[34] = PE534_finish;
    _zz_C_Valid_5[35] = PE535_finish;
    _zz_C_Valid_5[36] = PE536_finish;
    _zz_C_Valid_5[37] = PE537_finish;
    _zz_C_Valid_5[38] = PE538_finish;
    _zz_C_Valid_5[39] = PE539_finish;
    _zz_C_Valid_5[40] = PE540_finish;
    _zz_C_Valid_5[41] = PE541_finish;
    _zz_C_Valid_5[42] = PE542_finish;
    _zz_C_Valid_5[43] = PE543_finish;
    _zz_C_Valid_5[44] = PE544_finish;
    _zz_C_Valid_5[45] = PE545_finish;
    _zz_C_Valid_5[46] = PE546_finish;
    _zz_C_Valid_5[47] = PE547_finish;
    _zz_C_Valid_5[48] = PE548_finish;
    _zz_C_Valid_5[49] = PE549_finish;
    _zz_C_Valid_5[50] = PE550_finish;
    _zz_C_Valid_5[51] = PE551_finish;
    _zz_C_Valid_5[52] = PE552_finish;
    _zz_C_Valid_5[53] = PE553_finish;
    _zz_C_Valid_5[54] = PE554_finish;
    _zz_C_Valid_5[55] = PE555_finish;
    _zz_C_Valid_5[56] = PE556_finish;
    _zz_C_Valid_5[57] = PE557_finish;
    _zz_C_Valid_5[58] = PE558_finish;
    _zz_C_Valid_5[59] = PE559_finish;
    _zz_C_Valid_5[60] = PE560_finish;
    _zz_C_Valid_5[61] = PE561_finish;
    _zz_C_Valid_5[62] = PE562_finish;
    _zz_C_Valid_5[63] = PE563_finish;
  end

  assign C_Valid_5 = (|_zz_C_Valid_5);
  always @(*) begin
    MatrixC_6 = 32'h0;
    if(PE60_finish) begin
      MatrixC_6 = PE60_PE_OUT;
    end
    if(PE61_finish) begin
      MatrixC_6 = PE61_PE_OUT;
    end
    if(PE62_finish) begin
      MatrixC_6 = PE62_PE_OUT;
    end
    if(PE63_finish) begin
      MatrixC_6 = PE63_PE_OUT;
    end
    if(PE64_finish) begin
      MatrixC_6 = PE64_PE_OUT;
    end
    if(PE65_finish) begin
      MatrixC_6 = PE65_PE_OUT;
    end
    if(PE66_finish) begin
      MatrixC_6 = PE66_PE_OUT;
    end
    if(PE67_finish) begin
      MatrixC_6 = PE67_PE_OUT;
    end
    if(PE68_finish) begin
      MatrixC_6 = PE68_PE_OUT;
    end
    if(PE69_finish) begin
      MatrixC_6 = PE69_PE_OUT;
    end
    if(PE610_finish) begin
      MatrixC_6 = PE610_PE_OUT;
    end
    if(PE611_finish) begin
      MatrixC_6 = PE611_PE_OUT;
    end
    if(PE612_finish) begin
      MatrixC_6 = PE612_PE_OUT;
    end
    if(PE613_finish) begin
      MatrixC_6 = PE613_PE_OUT;
    end
    if(PE614_finish) begin
      MatrixC_6 = PE614_PE_OUT;
    end
    if(PE615_finish) begin
      MatrixC_6 = PE615_PE_OUT;
    end
    if(PE616_finish) begin
      MatrixC_6 = PE616_PE_OUT;
    end
    if(PE617_finish) begin
      MatrixC_6 = PE617_PE_OUT;
    end
    if(PE618_finish) begin
      MatrixC_6 = PE618_PE_OUT;
    end
    if(PE619_finish) begin
      MatrixC_6 = PE619_PE_OUT;
    end
    if(PE620_finish) begin
      MatrixC_6 = PE620_PE_OUT;
    end
    if(PE621_finish) begin
      MatrixC_6 = PE621_PE_OUT;
    end
    if(PE622_finish) begin
      MatrixC_6 = PE622_PE_OUT;
    end
    if(PE623_finish) begin
      MatrixC_6 = PE623_PE_OUT;
    end
    if(PE624_finish) begin
      MatrixC_6 = PE624_PE_OUT;
    end
    if(PE625_finish) begin
      MatrixC_6 = PE625_PE_OUT;
    end
    if(PE626_finish) begin
      MatrixC_6 = PE626_PE_OUT;
    end
    if(PE627_finish) begin
      MatrixC_6 = PE627_PE_OUT;
    end
    if(PE628_finish) begin
      MatrixC_6 = PE628_PE_OUT;
    end
    if(PE629_finish) begin
      MatrixC_6 = PE629_PE_OUT;
    end
    if(PE630_finish) begin
      MatrixC_6 = PE630_PE_OUT;
    end
    if(PE631_finish) begin
      MatrixC_6 = PE631_PE_OUT;
    end
    if(PE632_finish) begin
      MatrixC_6 = PE632_PE_OUT;
    end
    if(PE633_finish) begin
      MatrixC_6 = PE633_PE_OUT;
    end
    if(PE634_finish) begin
      MatrixC_6 = PE634_PE_OUT;
    end
    if(PE635_finish) begin
      MatrixC_6 = PE635_PE_OUT;
    end
    if(PE636_finish) begin
      MatrixC_6 = PE636_PE_OUT;
    end
    if(PE637_finish) begin
      MatrixC_6 = PE637_PE_OUT;
    end
    if(PE638_finish) begin
      MatrixC_6 = PE638_PE_OUT;
    end
    if(PE639_finish) begin
      MatrixC_6 = PE639_PE_OUT;
    end
    if(PE640_finish) begin
      MatrixC_6 = PE640_PE_OUT;
    end
    if(PE641_finish) begin
      MatrixC_6 = PE641_PE_OUT;
    end
    if(PE642_finish) begin
      MatrixC_6 = PE642_PE_OUT;
    end
    if(PE643_finish) begin
      MatrixC_6 = PE643_PE_OUT;
    end
    if(PE644_finish) begin
      MatrixC_6 = PE644_PE_OUT;
    end
    if(PE645_finish) begin
      MatrixC_6 = PE645_PE_OUT;
    end
    if(PE646_finish) begin
      MatrixC_6 = PE646_PE_OUT;
    end
    if(PE647_finish) begin
      MatrixC_6 = PE647_PE_OUT;
    end
    if(PE648_finish) begin
      MatrixC_6 = PE648_PE_OUT;
    end
    if(PE649_finish) begin
      MatrixC_6 = PE649_PE_OUT;
    end
    if(PE650_finish) begin
      MatrixC_6 = PE650_PE_OUT;
    end
    if(PE651_finish) begin
      MatrixC_6 = PE651_PE_OUT;
    end
    if(PE652_finish) begin
      MatrixC_6 = PE652_PE_OUT;
    end
    if(PE653_finish) begin
      MatrixC_6 = PE653_PE_OUT;
    end
    if(PE654_finish) begin
      MatrixC_6 = PE654_PE_OUT;
    end
    if(PE655_finish) begin
      MatrixC_6 = PE655_PE_OUT;
    end
    if(PE656_finish) begin
      MatrixC_6 = PE656_PE_OUT;
    end
    if(PE657_finish) begin
      MatrixC_6 = PE657_PE_OUT;
    end
    if(PE658_finish) begin
      MatrixC_6 = PE658_PE_OUT;
    end
    if(PE659_finish) begin
      MatrixC_6 = PE659_PE_OUT;
    end
    if(PE660_finish) begin
      MatrixC_6 = PE660_PE_OUT;
    end
    if(PE661_finish) begin
      MatrixC_6 = PE661_PE_OUT;
    end
    if(PE662_finish) begin
      MatrixC_6 = PE662_PE_OUT;
    end
    if(PE663_finish) begin
      MatrixC_6 = PE663_PE_OUT;
    end
  end

  always @(*) begin
    _zz_C_Valid_6[0] = PE60_finish;
    _zz_C_Valid_6[1] = PE61_finish;
    _zz_C_Valid_6[2] = PE62_finish;
    _zz_C_Valid_6[3] = PE63_finish;
    _zz_C_Valid_6[4] = PE64_finish;
    _zz_C_Valid_6[5] = PE65_finish;
    _zz_C_Valid_6[6] = PE66_finish;
    _zz_C_Valid_6[7] = PE67_finish;
    _zz_C_Valid_6[8] = PE68_finish;
    _zz_C_Valid_6[9] = PE69_finish;
    _zz_C_Valid_6[10] = PE610_finish;
    _zz_C_Valid_6[11] = PE611_finish;
    _zz_C_Valid_6[12] = PE612_finish;
    _zz_C_Valid_6[13] = PE613_finish;
    _zz_C_Valid_6[14] = PE614_finish;
    _zz_C_Valid_6[15] = PE615_finish;
    _zz_C_Valid_6[16] = PE616_finish;
    _zz_C_Valid_6[17] = PE617_finish;
    _zz_C_Valid_6[18] = PE618_finish;
    _zz_C_Valid_6[19] = PE619_finish;
    _zz_C_Valid_6[20] = PE620_finish;
    _zz_C_Valid_6[21] = PE621_finish;
    _zz_C_Valid_6[22] = PE622_finish;
    _zz_C_Valid_6[23] = PE623_finish;
    _zz_C_Valid_6[24] = PE624_finish;
    _zz_C_Valid_6[25] = PE625_finish;
    _zz_C_Valid_6[26] = PE626_finish;
    _zz_C_Valid_6[27] = PE627_finish;
    _zz_C_Valid_6[28] = PE628_finish;
    _zz_C_Valid_6[29] = PE629_finish;
    _zz_C_Valid_6[30] = PE630_finish;
    _zz_C_Valid_6[31] = PE631_finish;
    _zz_C_Valid_6[32] = PE632_finish;
    _zz_C_Valid_6[33] = PE633_finish;
    _zz_C_Valid_6[34] = PE634_finish;
    _zz_C_Valid_6[35] = PE635_finish;
    _zz_C_Valid_6[36] = PE636_finish;
    _zz_C_Valid_6[37] = PE637_finish;
    _zz_C_Valid_6[38] = PE638_finish;
    _zz_C_Valid_6[39] = PE639_finish;
    _zz_C_Valid_6[40] = PE640_finish;
    _zz_C_Valid_6[41] = PE641_finish;
    _zz_C_Valid_6[42] = PE642_finish;
    _zz_C_Valid_6[43] = PE643_finish;
    _zz_C_Valid_6[44] = PE644_finish;
    _zz_C_Valid_6[45] = PE645_finish;
    _zz_C_Valid_6[46] = PE646_finish;
    _zz_C_Valid_6[47] = PE647_finish;
    _zz_C_Valid_6[48] = PE648_finish;
    _zz_C_Valid_6[49] = PE649_finish;
    _zz_C_Valid_6[50] = PE650_finish;
    _zz_C_Valid_6[51] = PE651_finish;
    _zz_C_Valid_6[52] = PE652_finish;
    _zz_C_Valid_6[53] = PE653_finish;
    _zz_C_Valid_6[54] = PE654_finish;
    _zz_C_Valid_6[55] = PE655_finish;
    _zz_C_Valid_6[56] = PE656_finish;
    _zz_C_Valid_6[57] = PE657_finish;
    _zz_C_Valid_6[58] = PE658_finish;
    _zz_C_Valid_6[59] = PE659_finish;
    _zz_C_Valid_6[60] = PE660_finish;
    _zz_C_Valid_6[61] = PE661_finish;
    _zz_C_Valid_6[62] = PE662_finish;
    _zz_C_Valid_6[63] = PE663_finish;
  end

  assign C_Valid_6 = (|_zz_C_Valid_6);
  always @(*) begin
    MatrixC_7 = 32'h0;
    if(PE70_finish) begin
      MatrixC_7 = PE70_PE_OUT;
    end
    if(PE71_finish) begin
      MatrixC_7 = PE71_PE_OUT;
    end
    if(PE72_finish) begin
      MatrixC_7 = PE72_PE_OUT;
    end
    if(PE73_finish) begin
      MatrixC_7 = PE73_PE_OUT;
    end
    if(PE74_finish) begin
      MatrixC_7 = PE74_PE_OUT;
    end
    if(PE75_finish) begin
      MatrixC_7 = PE75_PE_OUT;
    end
    if(PE76_finish) begin
      MatrixC_7 = PE76_PE_OUT;
    end
    if(PE77_finish) begin
      MatrixC_7 = PE77_PE_OUT;
    end
    if(PE78_finish) begin
      MatrixC_7 = PE78_PE_OUT;
    end
    if(PE79_finish) begin
      MatrixC_7 = PE79_PE_OUT;
    end
    if(PE710_finish) begin
      MatrixC_7 = PE710_PE_OUT;
    end
    if(PE711_finish) begin
      MatrixC_7 = PE711_PE_OUT;
    end
    if(PE712_finish) begin
      MatrixC_7 = PE712_PE_OUT;
    end
    if(PE713_finish) begin
      MatrixC_7 = PE713_PE_OUT;
    end
    if(PE714_finish) begin
      MatrixC_7 = PE714_PE_OUT;
    end
    if(PE715_finish) begin
      MatrixC_7 = PE715_PE_OUT;
    end
    if(PE716_finish) begin
      MatrixC_7 = PE716_PE_OUT;
    end
    if(PE717_finish) begin
      MatrixC_7 = PE717_PE_OUT;
    end
    if(PE718_finish) begin
      MatrixC_7 = PE718_PE_OUT;
    end
    if(PE719_finish) begin
      MatrixC_7 = PE719_PE_OUT;
    end
    if(PE720_finish) begin
      MatrixC_7 = PE720_PE_OUT;
    end
    if(PE721_finish) begin
      MatrixC_7 = PE721_PE_OUT;
    end
    if(PE722_finish) begin
      MatrixC_7 = PE722_PE_OUT;
    end
    if(PE723_finish) begin
      MatrixC_7 = PE723_PE_OUT;
    end
    if(PE724_finish) begin
      MatrixC_7 = PE724_PE_OUT;
    end
    if(PE725_finish) begin
      MatrixC_7 = PE725_PE_OUT;
    end
    if(PE726_finish) begin
      MatrixC_7 = PE726_PE_OUT;
    end
    if(PE727_finish) begin
      MatrixC_7 = PE727_PE_OUT;
    end
    if(PE728_finish) begin
      MatrixC_7 = PE728_PE_OUT;
    end
    if(PE729_finish) begin
      MatrixC_7 = PE729_PE_OUT;
    end
    if(PE730_finish) begin
      MatrixC_7 = PE730_PE_OUT;
    end
    if(PE731_finish) begin
      MatrixC_7 = PE731_PE_OUT;
    end
    if(PE732_finish) begin
      MatrixC_7 = PE732_PE_OUT;
    end
    if(PE733_finish) begin
      MatrixC_7 = PE733_PE_OUT;
    end
    if(PE734_finish) begin
      MatrixC_7 = PE734_PE_OUT;
    end
    if(PE735_finish) begin
      MatrixC_7 = PE735_PE_OUT;
    end
    if(PE736_finish) begin
      MatrixC_7 = PE736_PE_OUT;
    end
    if(PE737_finish) begin
      MatrixC_7 = PE737_PE_OUT;
    end
    if(PE738_finish) begin
      MatrixC_7 = PE738_PE_OUT;
    end
    if(PE739_finish) begin
      MatrixC_7 = PE739_PE_OUT;
    end
    if(PE740_finish) begin
      MatrixC_7 = PE740_PE_OUT;
    end
    if(PE741_finish) begin
      MatrixC_7 = PE741_PE_OUT;
    end
    if(PE742_finish) begin
      MatrixC_7 = PE742_PE_OUT;
    end
    if(PE743_finish) begin
      MatrixC_7 = PE743_PE_OUT;
    end
    if(PE744_finish) begin
      MatrixC_7 = PE744_PE_OUT;
    end
    if(PE745_finish) begin
      MatrixC_7 = PE745_PE_OUT;
    end
    if(PE746_finish) begin
      MatrixC_7 = PE746_PE_OUT;
    end
    if(PE747_finish) begin
      MatrixC_7 = PE747_PE_OUT;
    end
    if(PE748_finish) begin
      MatrixC_7 = PE748_PE_OUT;
    end
    if(PE749_finish) begin
      MatrixC_7 = PE749_PE_OUT;
    end
    if(PE750_finish) begin
      MatrixC_7 = PE750_PE_OUT;
    end
    if(PE751_finish) begin
      MatrixC_7 = PE751_PE_OUT;
    end
    if(PE752_finish) begin
      MatrixC_7 = PE752_PE_OUT;
    end
    if(PE753_finish) begin
      MatrixC_7 = PE753_PE_OUT;
    end
    if(PE754_finish) begin
      MatrixC_7 = PE754_PE_OUT;
    end
    if(PE755_finish) begin
      MatrixC_7 = PE755_PE_OUT;
    end
    if(PE756_finish) begin
      MatrixC_7 = PE756_PE_OUT;
    end
    if(PE757_finish) begin
      MatrixC_7 = PE757_PE_OUT;
    end
    if(PE758_finish) begin
      MatrixC_7 = PE758_PE_OUT;
    end
    if(PE759_finish) begin
      MatrixC_7 = PE759_PE_OUT;
    end
    if(PE760_finish) begin
      MatrixC_7 = PE760_PE_OUT;
    end
    if(PE761_finish) begin
      MatrixC_7 = PE761_PE_OUT;
    end
    if(PE762_finish) begin
      MatrixC_7 = PE762_PE_OUT;
    end
    if(PE763_finish) begin
      MatrixC_7 = PE763_PE_OUT;
    end
  end

  always @(*) begin
    _zz_C_Valid_7[0] = PE70_finish;
    _zz_C_Valid_7[1] = PE71_finish;
    _zz_C_Valid_7[2] = PE72_finish;
    _zz_C_Valid_7[3] = PE73_finish;
    _zz_C_Valid_7[4] = PE74_finish;
    _zz_C_Valid_7[5] = PE75_finish;
    _zz_C_Valid_7[6] = PE76_finish;
    _zz_C_Valid_7[7] = PE77_finish;
    _zz_C_Valid_7[8] = PE78_finish;
    _zz_C_Valid_7[9] = PE79_finish;
    _zz_C_Valid_7[10] = PE710_finish;
    _zz_C_Valid_7[11] = PE711_finish;
    _zz_C_Valid_7[12] = PE712_finish;
    _zz_C_Valid_7[13] = PE713_finish;
    _zz_C_Valid_7[14] = PE714_finish;
    _zz_C_Valid_7[15] = PE715_finish;
    _zz_C_Valid_7[16] = PE716_finish;
    _zz_C_Valid_7[17] = PE717_finish;
    _zz_C_Valid_7[18] = PE718_finish;
    _zz_C_Valid_7[19] = PE719_finish;
    _zz_C_Valid_7[20] = PE720_finish;
    _zz_C_Valid_7[21] = PE721_finish;
    _zz_C_Valid_7[22] = PE722_finish;
    _zz_C_Valid_7[23] = PE723_finish;
    _zz_C_Valid_7[24] = PE724_finish;
    _zz_C_Valid_7[25] = PE725_finish;
    _zz_C_Valid_7[26] = PE726_finish;
    _zz_C_Valid_7[27] = PE727_finish;
    _zz_C_Valid_7[28] = PE728_finish;
    _zz_C_Valid_7[29] = PE729_finish;
    _zz_C_Valid_7[30] = PE730_finish;
    _zz_C_Valid_7[31] = PE731_finish;
    _zz_C_Valid_7[32] = PE732_finish;
    _zz_C_Valid_7[33] = PE733_finish;
    _zz_C_Valid_7[34] = PE734_finish;
    _zz_C_Valid_7[35] = PE735_finish;
    _zz_C_Valid_7[36] = PE736_finish;
    _zz_C_Valid_7[37] = PE737_finish;
    _zz_C_Valid_7[38] = PE738_finish;
    _zz_C_Valid_7[39] = PE739_finish;
    _zz_C_Valid_7[40] = PE740_finish;
    _zz_C_Valid_7[41] = PE741_finish;
    _zz_C_Valid_7[42] = PE742_finish;
    _zz_C_Valid_7[43] = PE743_finish;
    _zz_C_Valid_7[44] = PE744_finish;
    _zz_C_Valid_7[45] = PE745_finish;
    _zz_C_Valid_7[46] = PE746_finish;
    _zz_C_Valid_7[47] = PE747_finish;
    _zz_C_Valid_7[48] = PE748_finish;
    _zz_C_Valid_7[49] = PE749_finish;
    _zz_C_Valid_7[50] = PE750_finish;
    _zz_C_Valid_7[51] = PE751_finish;
    _zz_C_Valid_7[52] = PE752_finish;
    _zz_C_Valid_7[53] = PE753_finish;
    _zz_C_Valid_7[54] = PE754_finish;
    _zz_C_Valid_7[55] = PE755_finish;
    _zz_C_Valid_7[56] = PE756_finish;
    _zz_C_Valid_7[57] = PE757_finish;
    _zz_C_Valid_7[58] = PE758_finish;
    _zz_C_Valid_7[59] = PE759_finish;
    _zz_C_Valid_7[60] = PE760_finish;
    _zz_C_Valid_7[61] = PE761_finish;
    _zz_C_Valid_7[62] = PE762_finish;
    _zz_C_Valid_7[63] = PE763_finish;
  end

  assign C_Valid_7 = (|_zz_C_Valid_7);
  assign PE00_valid = (io_A_Valid_0 && io_B_Valid_0);
  assign PE01_valid = (io_A_Valid_0_delay_1 && io_B_Valid_1);
  assign PE02_valid = (io_A_Valid_0_delay_2 && io_B_Valid_2);
  assign PE03_valid = (io_A_Valid_0_delay_3 && io_B_Valid_3);
  assign PE04_valid = (io_A_Valid_0_delay_4 && io_B_Valid_4);
  assign PE05_valid = (io_A_Valid_0_delay_5 && io_B_Valid_5);
  assign PE06_valid = (io_A_Valid_0_delay_6 && io_B_Valid_6);
  assign PE07_valid = (io_A_Valid_0_delay_7 && io_B_Valid_7);
  assign PE08_valid = (io_A_Valid_0_delay_8 && io_B_Valid_8);
  assign PE09_valid = (io_A_Valid_0_delay_9 && io_B_Valid_9);
  assign PE010_valid = (io_A_Valid_0_delay_10 && io_B_Valid_10);
  assign PE011_valid = (io_A_Valid_0_delay_11 && io_B_Valid_11);
  assign PE012_valid = (io_A_Valid_0_delay_12 && io_B_Valid_12);
  assign PE013_valid = (io_A_Valid_0_delay_13 && io_B_Valid_13);
  assign PE014_valid = (io_A_Valid_0_delay_14 && io_B_Valid_14);
  assign PE015_valid = (io_A_Valid_0_delay_15 && io_B_Valid_15);
  assign PE016_valid = (io_A_Valid_0_delay_16 && io_B_Valid_16);
  assign PE017_valid = (io_A_Valid_0_delay_17 && io_B_Valid_17);
  assign PE018_valid = (io_A_Valid_0_delay_18 && io_B_Valid_18);
  assign PE019_valid = (io_A_Valid_0_delay_19 && io_B_Valid_19);
  assign PE020_valid = (io_A_Valid_0_delay_20 && io_B_Valid_20);
  assign PE021_valid = (io_A_Valid_0_delay_21 && io_B_Valid_21);
  assign PE022_valid = (io_A_Valid_0_delay_22 && io_B_Valid_22);
  assign PE023_valid = (io_A_Valid_0_delay_23 && io_B_Valid_23);
  assign PE024_valid = (io_A_Valid_0_delay_24 && io_B_Valid_24);
  assign PE025_valid = (io_A_Valid_0_delay_25 && io_B_Valid_25);
  assign PE026_valid = (io_A_Valid_0_delay_26 && io_B_Valid_26);
  assign PE027_valid = (io_A_Valid_0_delay_27 && io_B_Valid_27);
  assign PE028_valid = (io_A_Valid_0_delay_28 && io_B_Valid_28);
  assign PE029_valid = (io_A_Valid_0_delay_29 && io_B_Valid_29);
  assign PE030_valid = (io_A_Valid_0_delay_30 && io_B_Valid_30);
  assign PE031_valid = (io_A_Valid_0_delay_31 && io_B_Valid_31);
  assign PE032_valid = (io_A_Valid_0_delay_32 && io_B_Valid_32);
  assign PE033_valid = (io_A_Valid_0_delay_33 && io_B_Valid_33);
  assign PE034_valid = (io_A_Valid_0_delay_34 && io_B_Valid_34);
  assign PE035_valid = (io_A_Valid_0_delay_35 && io_B_Valid_35);
  assign PE036_valid = (io_A_Valid_0_delay_36 && io_B_Valid_36);
  assign PE037_valid = (io_A_Valid_0_delay_37 && io_B_Valid_37);
  assign PE038_valid = (io_A_Valid_0_delay_38 && io_B_Valid_38);
  assign PE039_valid = (io_A_Valid_0_delay_39 && io_B_Valid_39);
  assign PE040_valid = (io_A_Valid_0_delay_40 && io_B_Valid_40);
  assign PE041_valid = (io_A_Valid_0_delay_41 && io_B_Valid_41);
  assign PE042_valid = (io_A_Valid_0_delay_42 && io_B_Valid_42);
  assign PE043_valid = (io_A_Valid_0_delay_43 && io_B_Valid_43);
  assign PE044_valid = (io_A_Valid_0_delay_44 && io_B_Valid_44);
  assign PE045_valid = (io_A_Valid_0_delay_45 && io_B_Valid_45);
  assign PE046_valid = (io_A_Valid_0_delay_46 && io_B_Valid_46);
  assign PE047_valid = (io_A_Valid_0_delay_47 && io_B_Valid_47);
  assign PE048_valid = (io_A_Valid_0_delay_48 && io_B_Valid_48);
  assign PE049_valid = (io_A_Valid_0_delay_49 && io_B_Valid_49);
  assign PE050_valid = (io_A_Valid_0_delay_50 && io_B_Valid_50);
  assign PE051_valid = (io_A_Valid_0_delay_51 && io_B_Valid_51);
  assign PE052_valid = (io_A_Valid_0_delay_52 && io_B_Valid_52);
  assign PE053_valid = (io_A_Valid_0_delay_53 && io_B_Valid_53);
  assign PE054_valid = (io_A_Valid_0_delay_54 && io_B_Valid_54);
  assign PE055_valid = (io_A_Valid_0_delay_55 && io_B_Valid_55);
  assign PE056_valid = (io_A_Valid_0_delay_56 && io_B_Valid_56);
  assign PE057_valid = (io_A_Valid_0_delay_57 && io_B_Valid_57);
  assign PE058_valid = (io_A_Valid_0_delay_58 && io_B_Valid_58);
  assign PE059_valid = (io_A_Valid_0_delay_59 && io_B_Valid_59);
  assign PE060_valid = (io_A_Valid_0_delay_60 && io_B_Valid_60);
  assign PE061_valid = (io_A_Valid_0_delay_61 && io_B_Valid_61);
  assign PE062_valid = (io_A_Valid_0_delay_62 && io_B_Valid_62);
  assign PE063_valid = (io_A_Valid_0_delay_63 && io_B_Valid_63);
  assign PE10_valid = (io_A_Valid_1 && io_B_Valid_0_delay_1);
  assign PE11_valid = (io_A_Valid_1_delay_1 && io_B_Valid_1_delay_1);
  assign PE12_valid = (io_A_Valid_1_delay_2 && io_B_Valid_2_delay_1);
  assign PE13_valid = (io_A_Valid_1_delay_3 && io_B_Valid_3_delay_1);
  assign PE14_valid = (io_A_Valid_1_delay_4 && io_B_Valid_4_delay_1);
  assign PE15_valid = (io_A_Valid_1_delay_5 && io_B_Valid_5_delay_1);
  assign PE16_valid = (io_A_Valid_1_delay_6 && io_B_Valid_6_delay_1);
  assign PE17_valid = (io_A_Valid_1_delay_7 && io_B_Valid_7_delay_1);
  assign PE18_valid = (io_A_Valid_1_delay_8 && io_B_Valid_8_delay_1);
  assign PE19_valid = (io_A_Valid_1_delay_9 && io_B_Valid_9_delay_1);
  assign PE110_valid = (io_A_Valid_1_delay_10 && io_B_Valid_10_delay_1);
  assign PE111_valid = (io_A_Valid_1_delay_11 && io_B_Valid_11_delay_1);
  assign PE112_valid = (io_A_Valid_1_delay_12 && io_B_Valid_12_delay_1);
  assign PE113_valid = (io_A_Valid_1_delay_13 && io_B_Valid_13_delay_1);
  assign PE114_valid = (io_A_Valid_1_delay_14 && io_B_Valid_14_delay_1);
  assign PE115_valid = (io_A_Valid_1_delay_15 && io_B_Valid_15_delay_1);
  assign PE116_valid = (io_A_Valid_1_delay_16 && io_B_Valid_16_delay_1);
  assign PE117_valid = (io_A_Valid_1_delay_17 && io_B_Valid_17_delay_1);
  assign PE118_valid = (io_A_Valid_1_delay_18 && io_B_Valid_18_delay_1);
  assign PE119_valid = (io_A_Valid_1_delay_19 && io_B_Valid_19_delay_1);
  assign PE120_valid = (io_A_Valid_1_delay_20 && io_B_Valid_20_delay_1);
  assign PE121_valid = (io_A_Valid_1_delay_21 && io_B_Valid_21_delay_1);
  assign PE122_valid = (io_A_Valid_1_delay_22 && io_B_Valid_22_delay_1);
  assign PE123_valid = (io_A_Valid_1_delay_23 && io_B_Valid_23_delay_1);
  assign PE124_valid = (io_A_Valid_1_delay_24 && io_B_Valid_24_delay_1);
  assign PE125_valid = (io_A_Valid_1_delay_25 && io_B_Valid_25_delay_1);
  assign PE126_valid = (io_A_Valid_1_delay_26 && io_B_Valid_26_delay_1);
  assign PE127_valid = (io_A_Valid_1_delay_27 && io_B_Valid_27_delay_1);
  assign PE128_valid = (io_A_Valid_1_delay_28 && io_B_Valid_28_delay_1);
  assign PE129_valid = (io_A_Valid_1_delay_29 && io_B_Valid_29_delay_1);
  assign PE130_valid = (io_A_Valid_1_delay_30 && io_B_Valid_30_delay_1);
  assign PE131_valid = (io_A_Valid_1_delay_31 && io_B_Valid_31_delay_1);
  assign PE132_valid = (io_A_Valid_1_delay_32 && io_B_Valid_32_delay_1);
  assign PE133_valid = (io_A_Valid_1_delay_33 && io_B_Valid_33_delay_1);
  assign PE134_valid = (io_A_Valid_1_delay_34 && io_B_Valid_34_delay_1);
  assign PE135_valid = (io_A_Valid_1_delay_35 && io_B_Valid_35_delay_1);
  assign PE136_valid = (io_A_Valid_1_delay_36 && io_B_Valid_36_delay_1);
  assign PE137_valid = (io_A_Valid_1_delay_37 && io_B_Valid_37_delay_1);
  assign PE138_valid = (io_A_Valid_1_delay_38 && io_B_Valid_38_delay_1);
  assign PE139_valid = (io_A_Valid_1_delay_39 && io_B_Valid_39_delay_1);
  assign PE140_valid = (io_A_Valid_1_delay_40 && io_B_Valid_40_delay_1);
  assign PE141_valid = (io_A_Valid_1_delay_41 && io_B_Valid_41_delay_1);
  assign PE142_valid = (io_A_Valid_1_delay_42 && io_B_Valid_42_delay_1);
  assign PE143_valid = (io_A_Valid_1_delay_43 && io_B_Valid_43_delay_1);
  assign PE144_valid = (io_A_Valid_1_delay_44 && io_B_Valid_44_delay_1);
  assign PE145_valid = (io_A_Valid_1_delay_45 && io_B_Valid_45_delay_1);
  assign PE146_valid = (io_A_Valid_1_delay_46 && io_B_Valid_46_delay_1);
  assign PE147_valid = (io_A_Valid_1_delay_47 && io_B_Valid_47_delay_1);
  assign PE148_valid = (io_A_Valid_1_delay_48 && io_B_Valid_48_delay_1);
  assign PE149_valid = (io_A_Valid_1_delay_49 && io_B_Valid_49_delay_1);
  assign PE150_valid = (io_A_Valid_1_delay_50 && io_B_Valid_50_delay_1);
  assign PE151_valid = (io_A_Valid_1_delay_51 && io_B_Valid_51_delay_1);
  assign PE152_valid = (io_A_Valid_1_delay_52 && io_B_Valid_52_delay_1);
  assign PE153_valid = (io_A_Valid_1_delay_53 && io_B_Valid_53_delay_1);
  assign PE154_valid = (io_A_Valid_1_delay_54 && io_B_Valid_54_delay_1);
  assign PE155_valid = (io_A_Valid_1_delay_55 && io_B_Valid_55_delay_1);
  assign PE156_valid = (io_A_Valid_1_delay_56 && io_B_Valid_56_delay_1);
  assign PE157_valid = (io_A_Valid_1_delay_57 && io_B_Valid_57_delay_1);
  assign PE158_valid = (io_A_Valid_1_delay_58 && io_B_Valid_58_delay_1);
  assign PE159_valid = (io_A_Valid_1_delay_59 && io_B_Valid_59_delay_1);
  assign PE160_valid = (io_A_Valid_1_delay_60 && io_B_Valid_60_delay_1);
  assign PE161_valid = (io_A_Valid_1_delay_61 && io_B_Valid_61_delay_1);
  assign PE162_valid = (io_A_Valid_1_delay_62 && io_B_Valid_62_delay_1);
  assign PE163_valid = (io_A_Valid_1_delay_63 && io_B_Valid_63_delay_1);
  assign PE20_valid = (io_A_Valid_2 && io_B_Valid_0_delay_2);
  assign PE21_valid = (io_A_Valid_2_delay_1 && io_B_Valid_1_delay_2);
  assign PE22_valid = (io_A_Valid_2_delay_2 && io_B_Valid_2_delay_2);
  assign PE23_valid = (io_A_Valid_2_delay_3 && io_B_Valid_3_delay_2);
  assign PE24_valid = (io_A_Valid_2_delay_4 && io_B_Valid_4_delay_2);
  assign PE25_valid = (io_A_Valid_2_delay_5 && io_B_Valid_5_delay_2);
  assign PE26_valid = (io_A_Valid_2_delay_6 && io_B_Valid_6_delay_2);
  assign PE27_valid = (io_A_Valid_2_delay_7 && io_B_Valid_7_delay_2);
  assign PE28_valid = (io_A_Valid_2_delay_8 && io_B_Valid_8_delay_2);
  assign PE29_valid = (io_A_Valid_2_delay_9 && io_B_Valid_9_delay_2);
  assign PE210_valid = (io_A_Valid_2_delay_10 && io_B_Valid_10_delay_2);
  assign PE211_valid = (io_A_Valid_2_delay_11 && io_B_Valid_11_delay_2);
  assign PE212_valid = (io_A_Valid_2_delay_12 && io_B_Valid_12_delay_2);
  assign PE213_valid = (io_A_Valid_2_delay_13 && io_B_Valid_13_delay_2);
  assign PE214_valid = (io_A_Valid_2_delay_14 && io_B_Valid_14_delay_2);
  assign PE215_valid = (io_A_Valid_2_delay_15 && io_B_Valid_15_delay_2);
  assign PE216_valid = (io_A_Valid_2_delay_16 && io_B_Valid_16_delay_2);
  assign PE217_valid = (io_A_Valid_2_delay_17 && io_B_Valid_17_delay_2);
  assign PE218_valid = (io_A_Valid_2_delay_18 && io_B_Valid_18_delay_2);
  assign PE219_valid = (io_A_Valid_2_delay_19 && io_B_Valid_19_delay_2);
  assign PE220_valid = (io_A_Valid_2_delay_20 && io_B_Valid_20_delay_2);
  assign PE221_valid = (io_A_Valid_2_delay_21 && io_B_Valid_21_delay_2);
  assign PE222_valid = (io_A_Valid_2_delay_22 && io_B_Valid_22_delay_2);
  assign PE223_valid = (io_A_Valid_2_delay_23 && io_B_Valid_23_delay_2);
  assign PE224_valid = (io_A_Valid_2_delay_24 && io_B_Valid_24_delay_2);
  assign PE225_valid = (io_A_Valid_2_delay_25 && io_B_Valid_25_delay_2);
  assign PE226_valid = (io_A_Valid_2_delay_26 && io_B_Valid_26_delay_2);
  assign PE227_valid = (io_A_Valid_2_delay_27 && io_B_Valid_27_delay_2);
  assign PE228_valid = (io_A_Valid_2_delay_28 && io_B_Valid_28_delay_2);
  assign PE229_valid = (io_A_Valid_2_delay_29 && io_B_Valid_29_delay_2);
  assign PE230_valid = (io_A_Valid_2_delay_30 && io_B_Valid_30_delay_2);
  assign PE231_valid = (io_A_Valid_2_delay_31 && io_B_Valid_31_delay_2);
  assign PE232_valid = (io_A_Valid_2_delay_32 && io_B_Valid_32_delay_2);
  assign PE233_valid = (io_A_Valid_2_delay_33 && io_B_Valid_33_delay_2);
  assign PE234_valid = (io_A_Valid_2_delay_34 && io_B_Valid_34_delay_2);
  assign PE235_valid = (io_A_Valid_2_delay_35 && io_B_Valid_35_delay_2);
  assign PE236_valid = (io_A_Valid_2_delay_36 && io_B_Valid_36_delay_2);
  assign PE237_valid = (io_A_Valid_2_delay_37 && io_B_Valid_37_delay_2);
  assign PE238_valid = (io_A_Valid_2_delay_38 && io_B_Valid_38_delay_2);
  assign PE239_valid = (io_A_Valid_2_delay_39 && io_B_Valid_39_delay_2);
  assign PE240_valid = (io_A_Valid_2_delay_40 && io_B_Valid_40_delay_2);
  assign PE241_valid = (io_A_Valid_2_delay_41 && io_B_Valid_41_delay_2);
  assign PE242_valid = (io_A_Valid_2_delay_42 && io_B_Valid_42_delay_2);
  assign PE243_valid = (io_A_Valid_2_delay_43 && io_B_Valid_43_delay_2);
  assign PE244_valid = (io_A_Valid_2_delay_44 && io_B_Valid_44_delay_2);
  assign PE245_valid = (io_A_Valid_2_delay_45 && io_B_Valid_45_delay_2);
  assign PE246_valid = (io_A_Valid_2_delay_46 && io_B_Valid_46_delay_2);
  assign PE247_valid = (io_A_Valid_2_delay_47 && io_B_Valid_47_delay_2);
  assign PE248_valid = (io_A_Valid_2_delay_48 && io_B_Valid_48_delay_2);
  assign PE249_valid = (io_A_Valid_2_delay_49 && io_B_Valid_49_delay_2);
  assign PE250_valid = (io_A_Valid_2_delay_50 && io_B_Valid_50_delay_2);
  assign PE251_valid = (io_A_Valid_2_delay_51 && io_B_Valid_51_delay_2);
  assign PE252_valid = (io_A_Valid_2_delay_52 && io_B_Valid_52_delay_2);
  assign PE253_valid = (io_A_Valid_2_delay_53 && io_B_Valid_53_delay_2);
  assign PE254_valid = (io_A_Valid_2_delay_54 && io_B_Valid_54_delay_2);
  assign PE255_valid = (io_A_Valid_2_delay_55 && io_B_Valid_55_delay_2);
  assign PE256_valid = (io_A_Valid_2_delay_56 && io_B_Valid_56_delay_2);
  assign PE257_valid = (io_A_Valid_2_delay_57 && io_B_Valid_57_delay_2);
  assign PE258_valid = (io_A_Valid_2_delay_58 && io_B_Valid_58_delay_2);
  assign PE259_valid = (io_A_Valid_2_delay_59 && io_B_Valid_59_delay_2);
  assign PE260_valid = (io_A_Valid_2_delay_60 && io_B_Valid_60_delay_2);
  assign PE261_valid = (io_A_Valid_2_delay_61 && io_B_Valid_61_delay_2);
  assign PE262_valid = (io_A_Valid_2_delay_62 && io_B_Valid_62_delay_2);
  assign PE263_valid = (io_A_Valid_2_delay_63 && io_B_Valid_63_delay_2);
  assign PE30_valid = (io_A_Valid_3 && io_B_Valid_0_delay_3);
  assign PE31_valid = (io_A_Valid_3_delay_1 && io_B_Valid_1_delay_3);
  assign PE32_valid = (io_A_Valid_3_delay_2 && io_B_Valid_2_delay_3);
  assign PE33_valid = (io_A_Valid_3_delay_3 && io_B_Valid_3_delay_3);
  assign PE34_valid = (io_A_Valid_3_delay_4 && io_B_Valid_4_delay_3);
  assign PE35_valid = (io_A_Valid_3_delay_5 && io_B_Valid_5_delay_3);
  assign PE36_valid = (io_A_Valid_3_delay_6 && io_B_Valid_6_delay_3);
  assign PE37_valid = (io_A_Valid_3_delay_7 && io_B_Valid_7_delay_3);
  assign PE38_valid = (io_A_Valid_3_delay_8 && io_B_Valid_8_delay_3);
  assign PE39_valid = (io_A_Valid_3_delay_9 && io_B_Valid_9_delay_3);
  assign PE310_valid = (io_A_Valid_3_delay_10 && io_B_Valid_10_delay_3);
  assign PE311_valid = (io_A_Valid_3_delay_11 && io_B_Valid_11_delay_3);
  assign PE312_valid = (io_A_Valid_3_delay_12 && io_B_Valid_12_delay_3);
  assign PE313_valid = (io_A_Valid_3_delay_13 && io_B_Valid_13_delay_3);
  assign PE314_valid = (io_A_Valid_3_delay_14 && io_B_Valid_14_delay_3);
  assign PE315_valid = (io_A_Valid_3_delay_15 && io_B_Valid_15_delay_3);
  assign PE316_valid = (io_A_Valid_3_delay_16 && io_B_Valid_16_delay_3);
  assign PE317_valid = (io_A_Valid_3_delay_17 && io_B_Valid_17_delay_3);
  assign PE318_valid = (io_A_Valid_3_delay_18 && io_B_Valid_18_delay_3);
  assign PE319_valid = (io_A_Valid_3_delay_19 && io_B_Valid_19_delay_3);
  assign PE320_valid = (io_A_Valid_3_delay_20 && io_B_Valid_20_delay_3);
  assign PE321_valid = (io_A_Valid_3_delay_21 && io_B_Valid_21_delay_3);
  assign PE322_valid = (io_A_Valid_3_delay_22 && io_B_Valid_22_delay_3);
  assign PE323_valid = (io_A_Valid_3_delay_23 && io_B_Valid_23_delay_3);
  assign PE324_valid = (io_A_Valid_3_delay_24 && io_B_Valid_24_delay_3);
  assign PE325_valid = (io_A_Valid_3_delay_25 && io_B_Valid_25_delay_3);
  assign PE326_valid = (io_A_Valid_3_delay_26 && io_B_Valid_26_delay_3);
  assign PE327_valid = (io_A_Valid_3_delay_27 && io_B_Valid_27_delay_3);
  assign PE328_valid = (io_A_Valid_3_delay_28 && io_B_Valid_28_delay_3);
  assign PE329_valid = (io_A_Valid_3_delay_29 && io_B_Valid_29_delay_3);
  assign PE330_valid = (io_A_Valid_3_delay_30 && io_B_Valid_30_delay_3);
  assign PE331_valid = (io_A_Valid_3_delay_31 && io_B_Valid_31_delay_3);
  assign PE332_valid = (io_A_Valid_3_delay_32 && io_B_Valid_32_delay_3);
  assign PE333_valid = (io_A_Valid_3_delay_33 && io_B_Valid_33_delay_3);
  assign PE334_valid = (io_A_Valid_3_delay_34 && io_B_Valid_34_delay_3);
  assign PE335_valid = (io_A_Valid_3_delay_35 && io_B_Valid_35_delay_3);
  assign PE336_valid = (io_A_Valid_3_delay_36 && io_B_Valid_36_delay_3);
  assign PE337_valid = (io_A_Valid_3_delay_37 && io_B_Valid_37_delay_3);
  assign PE338_valid = (io_A_Valid_3_delay_38 && io_B_Valid_38_delay_3);
  assign PE339_valid = (io_A_Valid_3_delay_39 && io_B_Valid_39_delay_3);
  assign PE340_valid = (io_A_Valid_3_delay_40 && io_B_Valid_40_delay_3);
  assign PE341_valid = (io_A_Valid_3_delay_41 && io_B_Valid_41_delay_3);
  assign PE342_valid = (io_A_Valid_3_delay_42 && io_B_Valid_42_delay_3);
  assign PE343_valid = (io_A_Valid_3_delay_43 && io_B_Valid_43_delay_3);
  assign PE344_valid = (io_A_Valid_3_delay_44 && io_B_Valid_44_delay_3);
  assign PE345_valid = (io_A_Valid_3_delay_45 && io_B_Valid_45_delay_3);
  assign PE346_valid = (io_A_Valid_3_delay_46 && io_B_Valid_46_delay_3);
  assign PE347_valid = (io_A_Valid_3_delay_47 && io_B_Valid_47_delay_3);
  assign PE348_valid = (io_A_Valid_3_delay_48 && io_B_Valid_48_delay_3);
  assign PE349_valid = (io_A_Valid_3_delay_49 && io_B_Valid_49_delay_3);
  assign PE350_valid = (io_A_Valid_3_delay_50 && io_B_Valid_50_delay_3);
  assign PE351_valid = (io_A_Valid_3_delay_51 && io_B_Valid_51_delay_3);
  assign PE352_valid = (io_A_Valid_3_delay_52 && io_B_Valid_52_delay_3);
  assign PE353_valid = (io_A_Valid_3_delay_53 && io_B_Valid_53_delay_3);
  assign PE354_valid = (io_A_Valid_3_delay_54 && io_B_Valid_54_delay_3);
  assign PE355_valid = (io_A_Valid_3_delay_55 && io_B_Valid_55_delay_3);
  assign PE356_valid = (io_A_Valid_3_delay_56 && io_B_Valid_56_delay_3);
  assign PE357_valid = (io_A_Valid_3_delay_57 && io_B_Valid_57_delay_3);
  assign PE358_valid = (io_A_Valid_3_delay_58 && io_B_Valid_58_delay_3);
  assign PE359_valid = (io_A_Valid_3_delay_59 && io_B_Valid_59_delay_3);
  assign PE360_valid = (io_A_Valid_3_delay_60 && io_B_Valid_60_delay_3);
  assign PE361_valid = (io_A_Valid_3_delay_61 && io_B_Valid_61_delay_3);
  assign PE362_valid = (io_A_Valid_3_delay_62 && io_B_Valid_62_delay_3);
  assign PE363_valid = (io_A_Valid_3_delay_63 && io_B_Valid_63_delay_3);
  assign PE40_valid = (io_A_Valid_4 && io_B_Valid_0_delay_4);
  assign PE41_valid = (io_A_Valid_4_delay_1 && io_B_Valid_1_delay_4);
  assign PE42_valid = (io_A_Valid_4_delay_2 && io_B_Valid_2_delay_4);
  assign PE43_valid = (io_A_Valid_4_delay_3 && io_B_Valid_3_delay_4);
  assign PE44_valid = (io_A_Valid_4_delay_4 && io_B_Valid_4_delay_4);
  assign PE45_valid = (io_A_Valid_4_delay_5 && io_B_Valid_5_delay_4);
  assign PE46_valid = (io_A_Valid_4_delay_6 && io_B_Valid_6_delay_4);
  assign PE47_valid = (io_A_Valid_4_delay_7 && io_B_Valid_7_delay_4);
  assign PE48_valid = (io_A_Valid_4_delay_8 && io_B_Valid_8_delay_4);
  assign PE49_valid = (io_A_Valid_4_delay_9 && io_B_Valid_9_delay_4);
  assign PE410_valid = (io_A_Valid_4_delay_10 && io_B_Valid_10_delay_4);
  assign PE411_valid = (io_A_Valid_4_delay_11 && io_B_Valid_11_delay_4);
  assign PE412_valid = (io_A_Valid_4_delay_12 && io_B_Valid_12_delay_4);
  assign PE413_valid = (io_A_Valid_4_delay_13 && io_B_Valid_13_delay_4);
  assign PE414_valid = (io_A_Valid_4_delay_14 && io_B_Valid_14_delay_4);
  assign PE415_valid = (io_A_Valid_4_delay_15 && io_B_Valid_15_delay_4);
  assign PE416_valid = (io_A_Valid_4_delay_16 && io_B_Valid_16_delay_4);
  assign PE417_valid = (io_A_Valid_4_delay_17 && io_B_Valid_17_delay_4);
  assign PE418_valid = (io_A_Valid_4_delay_18 && io_B_Valid_18_delay_4);
  assign PE419_valid = (io_A_Valid_4_delay_19 && io_B_Valid_19_delay_4);
  assign PE420_valid = (io_A_Valid_4_delay_20 && io_B_Valid_20_delay_4);
  assign PE421_valid = (io_A_Valid_4_delay_21 && io_B_Valid_21_delay_4);
  assign PE422_valid = (io_A_Valid_4_delay_22 && io_B_Valid_22_delay_4);
  assign PE423_valid = (io_A_Valid_4_delay_23 && io_B_Valid_23_delay_4);
  assign PE424_valid = (io_A_Valid_4_delay_24 && io_B_Valid_24_delay_4);
  assign PE425_valid = (io_A_Valid_4_delay_25 && io_B_Valid_25_delay_4);
  assign PE426_valid = (io_A_Valid_4_delay_26 && io_B_Valid_26_delay_4);
  assign PE427_valid = (io_A_Valid_4_delay_27 && io_B_Valid_27_delay_4);
  assign PE428_valid = (io_A_Valid_4_delay_28 && io_B_Valid_28_delay_4);
  assign PE429_valid = (io_A_Valid_4_delay_29 && io_B_Valid_29_delay_4);
  assign PE430_valid = (io_A_Valid_4_delay_30 && io_B_Valid_30_delay_4);
  assign PE431_valid = (io_A_Valid_4_delay_31 && io_B_Valid_31_delay_4);
  assign PE432_valid = (io_A_Valid_4_delay_32 && io_B_Valid_32_delay_4);
  assign PE433_valid = (io_A_Valid_4_delay_33 && io_B_Valid_33_delay_4);
  assign PE434_valid = (io_A_Valid_4_delay_34 && io_B_Valid_34_delay_4);
  assign PE435_valid = (io_A_Valid_4_delay_35 && io_B_Valid_35_delay_4);
  assign PE436_valid = (io_A_Valid_4_delay_36 && io_B_Valid_36_delay_4);
  assign PE437_valid = (io_A_Valid_4_delay_37 && io_B_Valid_37_delay_4);
  assign PE438_valid = (io_A_Valid_4_delay_38 && io_B_Valid_38_delay_4);
  assign PE439_valid = (io_A_Valid_4_delay_39 && io_B_Valid_39_delay_4);
  assign PE440_valid = (io_A_Valid_4_delay_40 && io_B_Valid_40_delay_4);
  assign PE441_valid = (io_A_Valid_4_delay_41 && io_B_Valid_41_delay_4);
  assign PE442_valid = (io_A_Valid_4_delay_42 && io_B_Valid_42_delay_4);
  assign PE443_valid = (io_A_Valid_4_delay_43 && io_B_Valid_43_delay_4);
  assign PE444_valid = (io_A_Valid_4_delay_44 && io_B_Valid_44_delay_4);
  assign PE445_valid = (io_A_Valid_4_delay_45 && io_B_Valid_45_delay_4);
  assign PE446_valid = (io_A_Valid_4_delay_46 && io_B_Valid_46_delay_4);
  assign PE447_valid = (io_A_Valid_4_delay_47 && io_B_Valid_47_delay_4);
  assign PE448_valid = (io_A_Valid_4_delay_48 && io_B_Valid_48_delay_4);
  assign PE449_valid = (io_A_Valid_4_delay_49 && io_B_Valid_49_delay_4);
  assign PE450_valid = (io_A_Valid_4_delay_50 && io_B_Valid_50_delay_4);
  assign PE451_valid = (io_A_Valid_4_delay_51 && io_B_Valid_51_delay_4);
  assign PE452_valid = (io_A_Valid_4_delay_52 && io_B_Valid_52_delay_4);
  assign PE453_valid = (io_A_Valid_4_delay_53 && io_B_Valid_53_delay_4);
  assign PE454_valid = (io_A_Valid_4_delay_54 && io_B_Valid_54_delay_4);
  assign PE455_valid = (io_A_Valid_4_delay_55 && io_B_Valid_55_delay_4);
  assign PE456_valid = (io_A_Valid_4_delay_56 && io_B_Valid_56_delay_4);
  assign PE457_valid = (io_A_Valid_4_delay_57 && io_B_Valid_57_delay_4);
  assign PE458_valid = (io_A_Valid_4_delay_58 && io_B_Valid_58_delay_4);
  assign PE459_valid = (io_A_Valid_4_delay_59 && io_B_Valid_59_delay_4);
  assign PE460_valid = (io_A_Valid_4_delay_60 && io_B_Valid_60_delay_4);
  assign PE461_valid = (io_A_Valid_4_delay_61 && io_B_Valid_61_delay_4);
  assign PE462_valid = (io_A_Valid_4_delay_62 && io_B_Valid_62_delay_4);
  assign PE463_valid = (io_A_Valid_4_delay_63 && io_B_Valid_63_delay_4);
  assign PE50_valid = (io_A_Valid_5 && io_B_Valid_0_delay_5);
  assign PE51_valid = (io_A_Valid_5_delay_1 && io_B_Valid_1_delay_5);
  assign PE52_valid = (io_A_Valid_5_delay_2 && io_B_Valid_2_delay_5);
  assign PE53_valid = (io_A_Valid_5_delay_3 && io_B_Valid_3_delay_5);
  assign PE54_valid = (io_A_Valid_5_delay_4 && io_B_Valid_4_delay_5);
  assign PE55_valid = (io_A_Valid_5_delay_5 && io_B_Valid_5_delay_5);
  assign PE56_valid = (io_A_Valid_5_delay_6 && io_B_Valid_6_delay_5);
  assign PE57_valid = (io_A_Valid_5_delay_7 && io_B_Valid_7_delay_5);
  assign PE58_valid = (io_A_Valid_5_delay_8 && io_B_Valid_8_delay_5);
  assign PE59_valid = (io_A_Valid_5_delay_9 && io_B_Valid_9_delay_5);
  assign PE510_valid = (io_A_Valid_5_delay_10 && io_B_Valid_10_delay_5);
  assign PE511_valid = (io_A_Valid_5_delay_11 && io_B_Valid_11_delay_5);
  assign PE512_valid = (io_A_Valid_5_delay_12 && io_B_Valid_12_delay_5);
  assign PE513_valid = (io_A_Valid_5_delay_13 && io_B_Valid_13_delay_5);
  assign PE514_valid = (io_A_Valid_5_delay_14 && io_B_Valid_14_delay_5);
  assign PE515_valid = (io_A_Valid_5_delay_15 && io_B_Valid_15_delay_5);
  assign PE516_valid = (io_A_Valid_5_delay_16 && io_B_Valid_16_delay_5);
  assign PE517_valid = (io_A_Valid_5_delay_17 && io_B_Valid_17_delay_5);
  assign PE518_valid = (io_A_Valid_5_delay_18 && io_B_Valid_18_delay_5);
  assign PE519_valid = (io_A_Valid_5_delay_19 && io_B_Valid_19_delay_5);
  assign PE520_valid = (io_A_Valid_5_delay_20 && io_B_Valid_20_delay_5);
  assign PE521_valid = (io_A_Valid_5_delay_21 && io_B_Valid_21_delay_5);
  assign PE522_valid = (io_A_Valid_5_delay_22 && io_B_Valid_22_delay_5);
  assign PE523_valid = (io_A_Valid_5_delay_23 && io_B_Valid_23_delay_5);
  assign PE524_valid = (io_A_Valid_5_delay_24 && io_B_Valid_24_delay_5);
  assign PE525_valid = (io_A_Valid_5_delay_25 && io_B_Valid_25_delay_5);
  assign PE526_valid = (io_A_Valid_5_delay_26 && io_B_Valid_26_delay_5);
  assign PE527_valid = (io_A_Valid_5_delay_27 && io_B_Valid_27_delay_5);
  assign PE528_valid = (io_A_Valid_5_delay_28 && io_B_Valid_28_delay_5);
  assign PE529_valid = (io_A_Valid_5_delay_29 && io_B_Valid_29_delay_5);
  assign PE530_valid = (io_A_Valid_5_delay_30 && io_B_Valid_30_delay_5);
  assign PE531_valid = (io_A_Valid_5_delay_31 && io_B_Valid_31_delay_5);
  assign PE532_valid = (io_A_Valid_5_delay_32 && io_B_Valid_32_delay_5);
  assign PE533_valid = (io_A_Valid_5_delay_33 && io_B_Valid_33_delay_5);
  assign PE534_valid = (io_A_Valid_5_delay_34 && io_B_Valid_34_delay_5);
  assign PE535_valid = (io_A_Valid_5_delay_35 && io_B_Valid_35_delay_5);
  assign PE536_valid = (io_A_Valid_5_delay_36 && io_B_Valid_36_delay_5);
  assign PE537_valid = (io_A_Valid_5_delay_37 && io_B_Valid_37_delay_5);
  assign PE538_valid = (io_A_Valid_5_delay_38 && io_B_Valid_38_delay_5);
  assign PE539_valid = (io_A_Valid_5_delay_39 && io_B_Valid_39_delay_5);
  assign PE540_valid = (io_A_Valid_5_delay_40 && io_B_Valid_40_delay_5);
  assign PE541_valid = (io_A_Valid_5_delay_41 && io_B_Valid_41_delay_5);
  assign PE542_valid = (io_A_Valid_5_delay_42 && io_B_Valid_42_delay_5);
  assign PE543_valid = (io_A_Valid_5_delay_43 && io_B_Valid_43_delay_5);
  assign PE544_valid = (io_A_Valid_5_delay_44 && io_B_Valid_44_delay_5);
  assign PE545_valid = (io_A_Valid_5_delay_45 && io_B_Valid_45_delay_5);
  assign PE546_valid = (io_A_Valid_5_delay_46 && io_B_Valid_46_delay_5);
  assign PE547_valid = (io_A_Valid_5_delay_47 && io_B_Valid_47_delay_5);
  assign PE548_valid = (io_A_Valid_5_delay_48 && io_B_Valid_48_delay_5);
  assign PE549_valid = (io_A_Valid_5_delay_49 && io_B_Valid_49_delay_5);
  assign PE550_valid = (io_A_Valid_5_delay_50 && io_B_Valid_50_delay_5);
  assign PE551_valid = (io_A_Valid_5_delay_51 && io_B_Valid_51_delay_5);
  assign PE552_valid = (io_A_Valid_5_delay_52 && io_B_Valid_52_delay_5);
  assign PE553_valid = (io_A_Valid_5_delay_53 && io_B_Valid_53_delay_5);
  assign PE554_valid = (io_A_Valid_5_delay_54 && io_B_Valid_54_delay_5);
  assign PE555_valid = (io_A_Valid_5_delay_55 && io_B_Valid_55_delay_5);
  assign PE556_valid = (io_A_Valid_5_delay_56 && io_B_Valid_56_delay_5);
  assign PE557_valid = (io_A_Valid_5_delay_57 && io_B_Valid_57_delay_5);
  assign PE558_valid = (io_A_Valid_5_delay_58 && io_B_Valid_58_delay_5);
  assign PE559_valid = (io_A_Valid_5_delay_59 && io_B_Valid_59_delay_5);
  assign PE560_valid = (io_A_Valid_5_delay_60 && io_B_Valid_60_delay_5);
  assign PE561_valid = (io_A_Valid_5_delay_61 && io_B_Valid_61_delay_5);
  assign PE562_valid = (io_A_Valid_5_delay_62 && io_B_Valid_62_delay_5);
  assign PE563_valid = (io_A_Valid_5_delay_63 && io_B_Valid_63_delay_5);
  assign PE60_valid = (io_A_Valid_6 && io_B_Valid_0_delay_6);
  assign PE61_valid = (io_A_Valid_6_delay_1 && io_B_Valid_1_delay_6);
  assign PE62_valid = (io_A_Valid_6_delay_2 && io_B_Valid_2_delay_6);
  assign PE63_valid = (io_A_Valid_6_delay_3 && io_B_Valid_3_delay_6);
  assign PE64_valid = (io_A_Valid_6_delay_4 && io_B_Valid_4_delay_6);
  assign PE65_valid = (io_A_Valid_6_delay_5 && io_B_Valid_5_delay_6);
  assign PE66_valid = (io_A_Valid_6_delay_6 && io_B_Valid_6_delay_6);
  assign PE67_valid = (io_A_Valid_6_delay_7 && io_B_Valid_7_delay_6);
  assign PE68_valid = (io_A_Valid_6_delay_8 && io_B_Valid_8_delay_6);
  assign PE69_valid = (io_A_Valid_6_delay_9 && io_B_Valid_9_delay_6);
  assign PE610_valid = (io_A_Valid_6_delay_10 && io_B_Valid_10_delay_6);
  assign PE611_valid = (io_A_Valid_6_delay_11 && io_B_Valid_11_delay_6);
  assign PE612_valid = (io_A_Valid_6_delay_12 && io_B_Valid_12_delay_6);
  assign PE613_valid = (io_A_Valid_6_delay_13 && io_B_Valid_13_delay_6);
  assign PE614_valid = (io_A_Valid_6_delay_14 && io_B_Valid_14_delay_6);
  assign PE615_valid = (io_A_Valid_6_delay_15 && io_B_Valid_15_delay_6);
  assign PE616_valid = (io_A_Valid_6_delay_16 && io_B_Valid_16_delay_6);
  assign PE617_valid = (io_A_Valid_6_delay_17 && io_B_Valid_17_delay_6);
  assign PE618_valid = (io_A_Valid_6_delay_18 && io_B_Valid_18_delay_6);
  assign PE619_valid = (io_A_Valid_6_delay_19 && io_B_Valid_19_delay_6);
  assign PE620_valid = (io_A_Valid_6_delay_20 && io_B_Valid_20_delay_6);
  assign PE621_valid = (io_A_Valid_6_delay_21 && io_B_Valid_21_delay_6);
  assign PE622_valid = (io_A_Valid_6_delay_22 && io_B_Valid_22_delay_6);
  assign PE623_valid = (io_A_Valid_6_delay_23 && io_B_Valid_23_delay_6);
  assign PE624_valid = (io_A_Valid_6_delay_24 && io_B_Valid_24_delay_6);
  assign PE625_valid = (io_A_Valid_6_delay_25 && io_B_Valid_25_delay_6);
  assign PE626_valid = (io_A_Valid_6_delay_26 && io_B_Valid_26_delay_6);
  assign PE627_valid = (io_A_Valid_6_delay_27 && io_B_Valid_27_delay_6);
  assign PE628_valid = (io_A_Valid_6_delay_28 && io_B_Valid_28_delay_6);
  assign PE629_valid = (io_A_Valid_6_delay_29 && io_B_Valid_29_delay_6);
  assign PE630_valid = (io_A_Valid_6_delay_30 && io_B_Valid_30_delay_6);
  assign PE631_valid = (io_A_Valid_6_delay_31 && io_B_Valid_31_delay_6);
  assign PE632_valid = (io_A_Valid_6_delay_32 && io_B_Valid_32_delay_6);
  assign PE633_valid = (io_A_Valid_6_delay_33 && io_B_Valid_33_delay_6);
  assign PE634_valid = (io_A_Valid_6_delay_34 && io_B_Valid_34_delay_6);
  assign PE635_valid = (io_A_Valid_6_delay_35 && io_B_Valid_35_delay_6);
  assign PE636_valid = (io_A_Valid_6_delay_36 && io_B_Valid_36_delay_6);
  assign PE637_valid = (io_A_Valid_6_delay_37 && io_B_Valid_37_delay_6);
  assign PE638_valid = (io_A_Valid_6_delay_38 && io_B_Valid_38_delay_6);
  assign PE639_valid = (io_A_Valid_6_delay_39 && io_B_Valid_39_delay_6);
  assign PE640_valid = (io_A_Valid_6_delay_40 && io_B_Valid_40_delay_6);
  assign PE641_valid = (io_A_Valid_6_delay_41 && io_B_Valid_41_delay_6);
  assign PE642_valid = (io_A_Valid_6_delay_42 && io_B_Valid_42_delay_6);
  assign PE643_valid = (io_A_Valid_6_delay_43 && io_B_Valid_43_delay_6);
  assign PE644_valid = (io_A_Valid_6_delay_44 && io_B_Valid_44_delay_6);
  assign PE645_valid = (io_A_Valid_6_delay_45 && io_B_Valid_45_delay_6);
  assign PE646_valid = (io_A_Valid_6_delay_46 && io_B_Valid_46_delay_6);
  assign PE647_valid = (io_A_Valid_6_delay_47 && io_B_Valid_47_delay_6);
  assign PE648_valid = (io_A_Valid_6_delay_48 && io_B_Valid_48_delay_6);
  assign PE649_valid = (io_A_Valid_6_delay_49 && io_B_Valid_49_delay_6);
  assign PE650_valid = (io_A_Valid_6_delay_50 && io_B_Valid_50_delay_6);
  assign PE651_valid = (io_A_Valid_6_delay_51 && io_B_Valid_51_delay_6);
  assign PE652_valid = (io_A_Valid_6_delay_52 && io_B_Valid_52_delay_6);
  assign PE653_valid = (io_A_Valid_6_delay_53 && io_B_Valid_53_delay_6);
  assign PE654_valid = (io_A_Valid_6_delay_54 && io_B_Valid_54_delay_6);
  assign PE655_valid = (io_A_Valid_6_delay_55 && io_B_Valid_55_delay_6);
  assign PE656_valid = (io_A_Valid_6_delay_56 && io_B_Valid_56_delay_6);
  assign PE657_valid = (io_A_Valid_6_delay_57 && io_B_Valid_57_delay_6);
  assign PE658_valid = (io_A_Valid_6_delay_58 && io_B_Valid_58_delay_6);
  assign PE659_valid = (io_A_Valid_6_delay_59 && io_B_Valid_59_delay_6);
  assign PE660_valid = (io_A_Valid_6_delay_60 && io_B_Valid_60_delay_6);
  assign PE661_valid = (io_A_Valid_6_delay_61 && io_B_Valid_61_delay_6);
  assign PE662_valid = (io_A_Valid_6_delay_62 && io_B_Valid_62_delay_6);
  assign PE663_valid = (io_A_Valid_6_delay_63 && io_B_Valid_63_delay_6);
  assign PE70_valid = (io_A_Valid_7 && io_B_Valid_0_delay_7);
  assign PE71_valid = (io_A_Valid_7_delay_1 && io_B_Valid_1_delay_7);
  assign PE72_valid = (io_A_Valid_7_delay_2 && io_B_Valid_2_delay_7);
  assign PE73_valid = (io_A_Valid_7_delay_3 && io_B_Valid_3_delay_7);
  assign PE74_valid = (io_A_Valid_7_delay_4 && io_B_Valid_4_delay_7);
  assign PE75_valid = (io_A_Valid_7_delay_5 && io_B_Valid_5_delay_7);
  assign PE76_valid = (io_A_Valid_7_delay_6 && io_B_Valid_6_delay_7);
  assign PE77_valid = (io_A_Valid_7_delay_7 && io_B_Valid_7_delay_7);
  assign PE78_valid = (io_A_Valid_7_delay_8 && io_B_Valid_8_delay_7);
  assign PE79_valid = (io_A_Valid_7_delay_9 && io_B_Valid_9_delay_7);
  assign PE710_valid = (io_A_Valid_7_delay_10 && io_B_Valid_10_delay_7);
  assign PE711_valid = (io_A_Valid_7_delay_11 && io_B_Valid_11_delay_7);
  assign PE712_valid = (io_A_Valid_7_delay_12 && io_B_Valid_12_delay_7);
  assign PE713_valid = (io_A_Valid_7_delay_13 && io_B_Valid_13_delay_7);
  assign PE714_valid = (io_A_Valid_7_delay_14 && io_B_Valid_14_delay_7);
  assign PE715_valid = (io_A_Valid_7_delay_15 && io_B_Valid_15_delay_7);
  assign PE716_valid = (io_A_Valid_7_delay_16 && io_B_Valid_16_delay_7);
  assign PE717_valid = (io_A_Valid_7_delay_17 && io_B_Valid_17_delay_7);
  assign PE718_valid = (io_A_Valid_7_delay_18 && io_B_Valid_18_delay_7);
  assign PE719_valid = (io_A_Valid_7_delay_19 && io_B_Valid_19_delay_7);
  assign PE720_valid = (io_A_Valid_7_delay_20 && io_B_Valid_20_delay_7);
  assign PE721_valid = (io_A_Valid_7_delay_21 && io_B_Valid_21_delay_7);
  assign PE722_valid = (io_A_Valid_7_delay_22 && io_B_Valid_22_delay_7);
  assign PE723_valid = (io_A_Valid_7_delay_23 && io_B_Valid_23_delay_7);
  assign PE724_valid = (io_A_Valid_7_delay_24 && io_B_Valid_24_delay_7);
  assign PE725_valid = (io_A_Valid_7_delay_25 && io_B_Valid_25_delay_7);
  assign PE726_valid = (io_A_Valid_7_delay_26 && io_B_Valid_26_delay_7);
  assign PE727_valid = (io_A_Valid_7_delay_27 && io_B_Valid_27_delay_7);
  assign PE728_valid = (io_A_Valid_7_delay_28 && io_B_Valid_28_delay_7);
  assign PE729_valid = (io_A_Valid_7_delay_29 && io_B_Valid_29_delay_7);
  assign PE730_valid = (io_A_Valid_7_delay_30 && io_B_Valid_30_delay_7);
  assign PE731_valid = (io_A_Valid_7_delay_31 && io_B_Valid_31_delay_7);
  assign PE732_valid = (io_A_Valid_7_delay_32 && io_B_Valid_32_delay_7);
  assign PE733_valid = (io_A_Valid_7_delay_33 && io_B_Valid_33_delay_7);
  assign PE734_valid = (io_A_Valid_7_delay_34 && io_B_Valid_34_delay_7);
  assign PE735_valid = (io_A_Valid_7_delay_35 && io_B_Valid_35_delay_7);
  assign PE736_valid = (io_A_Valid_7_delay_36 && io_B_Valid_36_delay_7);
  assign PE737_valid = (io_A_Valid_7_delay_37 && io_B_Valid_37_delay_7);
  assign PE738_valid = (io_A_Valid_7_delay_38 && io_B_Valid_38_delay_7);
  assign PE739_valid = (io_A_Valid_7_delay_39 && io_B_Valid_39_delay_7);
  assign PE740_valid = (io_A_Valid_7_delay_40 && io_B_Valid_40_delay_7);
  assign PE741_valid = (io_A_Valid_7_delay_41 && io_B_Valid_41_delay_7);
  assign PE742_valid = (io_A_Valid_7_delay_42 && io_B_Valid_42_delay_7);
  assign PE743_valid = (io_A_Valid_7_delay_43 && io_B_Valid_43_delay_7);
  assign PE744_valid = (io_A_Valid_7_delay_44 && io_B_Valid_44_delay_7);
  assign PE745_valid = (io_A_Valid_7_delay_45 && io_B_Valid_45_delay_7);
  assign PE746_valid = (io_A_Valid_7_delay_46 && io_B_Valid_46_delay_7);
  assign PE747_valid = (io_A_Valid_7_delay_47 && io_B_Valid_47_delay_7);
  assign PE748_valid = (io_A_Valid_7_delay_48 && io_B_Valid_48_delay_7);
  assign PE749_valid = (io_A_Valid_7_delay_49 && io_B_Valid_49_delay_7);
  assign PE750_valid = (io_A_Valid_7_delay_50 && io_B_Valid_50_delay_7);
  assign PE751_valid = (io_A_Valid_7_delay_51 && io_B_Valid_51_delay_7);
  assign PE752_valid = (io_A_Valid_7_delay_52 && io_B_Valid_52_delay_7);
  assign PE753_valid = (io_A_Valid_7_delay_53 && io_B_Valid_53_delay_7);
  assign PE754_valid = (io_A_Valid_7_delay_54 && io_B_Valid_54_delay_7);
  assign PE755_valid = (io_A_Valid_7_delay_55 && io_B_Valid_55_delay_7);
  assign PE756_valid = (io_A_Valid_7_delay_56 && io_B_Valid_56_delay_7);
  assign PE757_valid = (io_A_Valid_7_delay_57 && io_B_Valid_57_delay_7);
  assign PE758_valid = (io_A_Valid_7_delay_58 && io_B_Valid_58_delay_7);
  assign PE759_valid = (io_A_Valid_7_delay_59 && io_B_Valid_59_delay_7);
  assign PE760_valid = (io_A_Valid_7_delay_60 && io_B_Valid_60_delay_7);
  assign PE761_valid = (io_A_Valid_7_delay_61 && io_B_Valid_61_delay_7);
  assign PE762_valid = (io_A_Valid_7_delay_62 && io_B_Valid_62_delay_7);
  assign PE763_valid = (io_A_Valid_7_delay_63 && io_B_Valid_63_delay_7);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      io_signCount_regNextWhen <= 16'h0;
      io_signCount_regNextWhen_1 <= 16'h0;
      io_signCount_regNextWhen_2 <= 16'h0;
      io_signCount_regNextWhen_3 <= 16'h0;
      io_signCount_regNextWhen_4 <= 16'h0;
      io_signCount_regNextWhen_5 <= 16'h0;
      io_signCount_regNextWhen_6 <= 16'h0;
      io_signCount_regNextWhen_7 <= 16'h0;
    end else begin
      if(start) begin
        io_signCount_regNextWhen <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_1 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_2 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_3 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_4 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_5 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_6 <= io_signCount;
      end
      if(start) begin
        io_signCount_regNextWhen_7 <= io_signCount;
      end
    end
  end

  always @(posedge clk) begin
    io_A_Valid_0_delay_1 <= io_A_Valid_0;
    io_A_Valid_0_delay_1_1 <= io_A_Valid_0;
    io_A_Valid_0_delay_2 <= io_A_Valid_0_delay_1_1;
    io_A_Valid_0_delay_1_2 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_1 <= io_A_Valid_0_delay_1_2;
    io_A_Valid_0_delay_3 <= io_A_Valid_0_delay_2_1;
    io_A_Valid_0_delay_1_3 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_2 <= io_A_Valid_0_delay_1_3;
    io_A_Valid_0_delay_3_1 <= io_A_Valid_0_delay_2_2;
    io_A_Valid_0_delay_4 <= io_A_Valid_0_delay_3_1;
    io_A_Valid_0_delay_1_4 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_3 <= io_A_Valid_0_delay_1_4;
    io_A_Valid_0_delay_3_2 <= io_A_Valid_0_delay_2_3;
    io_A_Valid_0_delay_4_1 <= io_A_Valid_0_delay_3_2;
    io_A_Valid_0_delay_5 <= io_A_Valid_0_delay_4_1;
    io_A_Valid_0_delay_1_5 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_4 <= io_A_Valid_0_delay_1_5;
    io_A_Valid_0_delay_3_3 <= io_A_Valid_0_delay_2_4;
    io_A_Valid_0_delay_4_2 <= io_A_Valid_0_delay_3_3;
    io_A_Valid_0_delay_5_1 <= io_A_Valid_0_delay_4_2;
    io_A_Valid_0_delay_6 <= io_A_Valid_0_delay_5_1;
    io_A_Valid_0_delay_1_6 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_5 <= io_A_Valid_0_delay_1_6;
    io_A_Valid_0_delay_3_4 <= io_A_Valid_0_delay_2_5;
    io_A_Valid_0_delay_4_3 <= io_A_Valid_0_delay_3_4;
    io_A_Valid_0_delay_5_2 <= io_A_Valid_0_delay_4_3;
    io_A_Valid_0_delay_6_1 <= io_A_Valid_0_delay_5_2;
    io_A_Valid_0_delay_7 <= io_A_Valid_0_delay_6_1;
    io_A_Valid_0_delay_1_7 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_6 <= io_A_Valid_0_delay_1_7;
    io_A_Valid_0_delay_3_5 <= io_A_Valid_0_delay_2_6;
    io_A_Valid_0_delay_4_4 <= io_A_Valid_0_delay_3_5;
    io_A_Valid_0_delay_5_3 <= io_A_Valid_0_delay_4_4;
    io_A_Valid_0_delay_6_2 <= io_A_Valid_0_delay_5_3;
    io_A_Valid_0_delay_7_1 <= io_A_Valid_0_delay_6_2;
    io_A_Valid_0_delay_8 <= io_A_Valid_0_delay_7_1;
    io_A_Valid_0_delay_1_8 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_7 <= io_A_Valid_0_delay_1_8;
    io_A_Valid_0_delay_3_6 <= io_A_Valid_0_delay_2_7;
    io_A_Valid_0_delay_4_5 <= io_A_Valid_0_delay_3_6;
    io_A_Valid_0_delay_5_4 <= io_A_Valid_0_delay_4_5;
    io_A_Valid_0_delay_6_3 <= io_A_Valid_0_delay_5_4;
    io_A_Valid_0_delay_7_2 <= io_A_Valid_0_delay_6_3;
    io_A_Valid_0_delay_8_1 <= io_A_Valid_0_delay_7_2;
    io_A_Valid_0_delay_9 <= io_A_Valid_0_delay_8_1;
    io_A_Valid_0_delay_1_9 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_8 <= io_A_Valid_0_delay_1_9;
    io_A_Valid_0_delay_3_7 <= io_A_Valid_0_delay_2_8;
    io_A_Valid_0_delay_4_6 <= io_A_Valid_0_delay_3_7;
    io_A_Valid_0_delay_5_5 <= io_A_Valid_0_delay_4_6;
    io_A_Valid_0_delay_6_4 <= io_A_Valid_0_delay_5_5;
    io_A_Valid_0_delay_7_3 <= io_A_Valid_0_delay_6_4;
    io_A_Valid_0_delay_8_2 <= io_A_Valid_0_delay_7_3;
    io_A_Valid_0_delay_9_1 <= io_A_Valid_0_delay_8_2;
    io_A_Valid_0_delay_10 <= io_A_Valid_0_delay_9_1;
    io_A_Valid_0_delay_1_10 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_9 <= io_A_Valid_0_delay_1_10;
    io_A_Valid_0_delay_3_8 <= io_A_Valid_0_delay_2_9;
    io_A_Valid_0_delay_4_7 <= io_A_Valid_0_delay_3_8;
    io_A_Valid_0_delay_5_6 <= io_A_Valid_0_delay_4_7;
    io_A_Valid_0_delay_6_5 <= io_A_Valid_0_delay_5_6;
    io_A_Valid_0_delay_7_4 <= io_A_Valid_0_delay_6_5;
    io_A_Valid_0_delay_8_3 <= io_A_Valid_0_delay_7_4;
    io_A_Valid_0_delay_9_2 <= io_A_Valid_0_delay_8_3;
    io_A_Valid_0_delay_10_1 <= io_A_Valid_0_delay_9_2;
    io_A_Valid_0_delay_11 <= io_A_Valid_0_delay_10_1;
    io_A_Valid_0_delay_1_11 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_10 <= io_A_Valid_0_delay_1_11;
    io_A_Valid_0_delay_3_9 <= io_A_Valid_0_delay_2_10;
    io_A_Valid_0_delay_4_8 <= io_A_Valid_0_delay_3_9;
    io_A_Valid_0_delay_5_7 <= io_A_Valid_0_delay_4_8;
    io_A_Valid_0_delay_6_6 <= io_A_Valid_0_delay_5_7;
    io_A_Valid_0_delay_7_5 <= io_A_Valid_0_delay_6_6;
    io_A_Valid_0_delay_8_4 <= io_A_Valid_0_delay_7_5;
    io_A_Valid_0_delay_9_3 <= io_A_Valid_0_delay_8_4;
    io_A_Valid_0_delay_10_2 <= io_A_Valid_0_delay_9_3;
    io_A_Valid_0_delay_11_1 <= io_A_Valid_0_delay_10_2;
    io_A_Valid_0_delay_12 <= io_A_Valid_0_delay_11_1;
    io_A_Valid_0_delay_1_12 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_11 <= io_A_Valid_0_delay_1_12;
    io_A_Valid_0_delay_3_10 <= io_A_Valid_0_delay_2_11;
    io_A_Valid_0_delay_4_9 <= io_A_Valid_0_delay_3_10;
    io_A_Valid_0_delay_5_8 <= io_A_Valid_0_delay_4_9;
    io_A_Valid_0_delay_6_7 <= io_A_Valid_0_delay_5_8;
    io_A_Valid_0_delay_7_6 <= io_A_Valid_0_delay_6_7;
    io_A_Valid_0_delay_8_5 <= io_A_Valid_0_delay_7_6;
    io_A_Valid_0_delay_9_4 <= io_A_Valid_0_delay_8_5;
    io_A_Valid_0_delay_10_3 <= io_A_Valid_0_delay_9_4;
    io_A_Valid_0_delay_11_2 <= io_A_Valid_0_delay_10_3;
    io_A_Valid_0_delay_12_1 <= io_A_Valid_0_delay_11_2;
    io_A_Valid_0_delay_13 <= io_A_Valid_0_delay_12_1;
    io_A_Valid_0_delay_1_13 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_12 <= io_A_Valid_0_delay_1_13;
    io_A_Valid_0_delay_3_11 <= io_A_Valid_0_delay_2_12;
    io_A_Valid_0_delay_4_10 <= io_A_Valid_0_delay_3_11;
    io_A_Valid_0_delay_5_9 <= io_A_Valid_0_delay_4_10;
    io_A_Valid_0_delay_6_8 <= io_A_Valid_0_delay_5_9;
    io_A_Valid_0_delay_7_7 <= io_A_Valid_0_delay_6_8;
    io_A_Valid_0_delay_8_6 <= io_A_Valid_0_delay_7_7;
    io_A_Valid_0_delay_9_5 <= io_A_Valid_0_delay_8_6;
    io_A_Valid_0_delay_10_4 <= io_A_Valid_0_delay_9_5;
    io_A_Valid_0_delay_11_3 <= io_A_Valid_0_delay_10_4;
    io_A_Valid_0_delay_12_2 <= io_A_Valid_0_delay_11_3;
    io_A_Valid_0_delay_13_1 <= io_A_Valid_0_delay_12_2;
    io_A_Valid_0_delay_14 <= io_A_Valid_0_delay_13_1;
    io_A_Valid_0_delay_1_14 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_13 <= io_A_Valid_0_delay_1_14;
    io_A_Valid_0_delay_3_12 <= io_A_Valid_0_delay_2_13;
    io_A_Valid_0_delay_4_11 <= io_A_Valid_0_delay_3_12;
    io_A_Valid_0_delay_5_10 <= io_A_Valid_0_delay_4_11;
    io_A_Valid_0_delay_6_9 <= io_A_Valid_0_delay_5_10;
    io_A_Valid_0_delay_7_8 <= io_A_Valid_0_delay_6_9;
    io_A_Valid_0_delay_8_7 <= io_A_Valid_0_delay_7_8;
    io_A_Valid_0_delay_9_6 <= io_A_Valid_0_delay_8_7;
    io_A_Valid_0_delay_10_5 <= io_A_Valid_0_delay_9_6;
    io_A_Valid_0_delay_11_4 <= io_A_Valid_0_delay_10_5;
    io_A_Valid_0_delay_12_3 <= io_A_Valid_0_delay_11_4;
    io_A_Valid_0_delay_13_2 <= io_A_Valid_0_delay_12_3;
    io_A_Valid_0_delay_14_1 <= io_A_Valid_0_delay_13_2;
    io_A_Valid_0_delay_15 <= io_A_Valid_0_delay_14_1;
    io_A_Valid_0_delay_1_15 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_14 <= io_A_Valid_0_delay_1_15;
    io_A_Valid_0_delay_3_13 <= io_A_Valid_0_delay_2_14;
    io_A_Valid_0_delay_4_12 <= io_A_Valid_0_delay_3_13;
    io_A_Valid_0_delay_5_11 <= io_A_Valid_0_delay_4_12;
    io_A_Valid_0_delay_6_10 <= io_A_Valid_0_delay_5_11;
    io_A_Valid_0_delay_7_9 <= io_A_Valid_0_delay_6_10;
    io_A_Valid_0_delay_8_8 <= io_A_Valid_0_delay_7_9;
    io_A_Valid_0_delay_9_7 <= io_A_Valid_0_delay_8_8;
    io_A_Valid_0_delay_10_6 <= io_A_Valid_0_delay_9_7;
    io_A_Valid_0_delay_11_5 <= io_A_Valid_0_delay_10_6;
    io_A_Valid_0_delay_12_4 <= io_A_Valid_0_delay_11_5;
    io_A_Valid_0_delay_13_3 <= io_A_Valid_0_delay_12_4;
    io_A_Valid_0_delay_14_2 <= io_A_Valid_0_delay_13_3;
    io_A_Valid_0_delay_15_1 <= io_A_Valid_0_delay_14_2;
    io_A_Valid_0_delay_16 <= io_A_Valid_0_delay_15_1;
    io_A_Valid_0_delay_1_16 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_15 <= io_A_Valid_0_delay_1_16;
    io_A_Valid_0_delay_3_14 <= io_A_Valid_0_delay_2_15;
    io_A_Valid_0_delay_4_13 <= io_A_Valid_0_delay_3_14;
    io_A_Valid_0_delay_5_12 <= io_A_Valid_0_delay_4_13;
    io_A_Valid_0_delay_6_11 <= io_A_Valid_0_delay_5_12;
    io_A_Valid_0_delay_7_10 <= io_A_Valid_0_delay_6_11;
    io_A_Valid_0_delay_8_9 <= io_A_Valid_0_delay_7_10;
    io_A_Valid_0_delay_9_8 <= io_A_Valid_0_delay_8_9;
    io_A_Valid_0_delay_10_7 <= io_A_Valid_0_delay_9_8;
    io_A_Valid_0_delay_11_6 <= io_A_Valid_0_delay_10_7;
    io_A_Valid_0_delay_12_5 <= io_A_Valid_0_delay_11_6;
    io_A_Valid_0_delay_13_4 <= io_A_Valid_0_delay_12_5;
    io_A_Valid_0_delay_14_3 <= io_A_Valid_0_delay_13_4;
    io_A_Valid_0_delay_15_2 <= io_A_Valid_0_delay_14_3;
    io_A_Valid_0_delay_16_1 <= io_A_Valid_0_delay_15_2;
    io_A_Valid_0_delay_17 <= io_A_Valid_0_delay_16_1;
    io_A_Valid_0_delay_1_17 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_16 <= io_A_Valid_0_delay_1_17;
    io_A_Valid_0_delay_3_15 <= io_A_Valid_0_delay_2_16;
    io_A_Valid_0_delay_4_14 <= io_A_Valid_0_delay_3_15;
    io_A_Valid_0_delay_5_13 <= io_A_Valid_0_delay_4_14;
    io_A_Valid_0_delay_6_12 <= io_A_Valid_0_delay_5_13;
    io_A_Valid_0_delay_7_11 <= io_A_Valid_0_delay_6_12;
    io_A_Valid_0_delay_8_10 <= io_A_Valid_0_delay_7_11;
    io_A_Valid_0_delay_9_9 <= io_A_Valid_0_delay_8_10;
    io_A_Valid_0_delay_10_8 <= io_A_Valid_0_delay_9_9;
    io_A_Valid_0_delay_11_7 <= io_A_Valid_0_delay_10_8;
    io_A_Valid_0_delay_12_6 <= io_A_Valid_0_delay_11_7;
    io_A_Valid_0_delay_13_5 <= io_A_Valid_0_delay_12_6;
    io_A_Valid_0_delay_14_4 <= io_A_Valid_0_delay_13_5;
    io_A_Valid_0_delay_15_3 <= io_A_Valid_0_delay_14_4;
    io_A_Valid_0_delay_16_2 <= io_A_Valid_0_delay_15_3;
    io_A_Valid_0_delay_17_1 <= io_A_Valid_0_delay_16_2;
    io_A_Valid_0_delay_18 <= io_A_Valid_0_delay_17_1;
    io_A_Valid_0_delay_1_18 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_17 <= io_A_Valid_0_delay_1_18;
    io_A_Valid_0_delay_3_16 <= io_A_Valid_0_delay_2_17;
    io_A_Valid_0_delay_4_15 <= io_A_Valid_0_delay_3_16;
    io_A_Valid_0_delay_5_14 <= io_A_Valid_0_delay_4_15;
    io_A_Valid_0_delay_6_13 <= io_A_Valid_0_delay_5_14;
    io_A_Valid_0_delay_7_12 <= io_A_Valid_0_delay_6_13;
    io_A_Valid_0_delay_8_11 <= io_A_Valid_0_delay_7_12;
    io_A_Valid_0_delay_9_10 <= io_A_Valid_0_delay_8_11;
    io_A_Valid_0_delay_10_9 <= io_A_Valid_0_delay_9_10;
    io_A_Valid_0_delay_11_8 <= io_A_Valid_0_delay_10_9;
    io_A_Valid_0_delay_12_7 <= io_A_Valid_0_delay_11_8;
    io_A_Valid_0_delay_13_6 <= io_A_Valid_0_delay_12_7;
    io_A_Valid_0_delay_14_5 <= io_A_Valid_0_delay_13_6;
    io_A_Valid_0_delay_15_4 <= io_A_Valid_0_delay_14_5;
    io_A_Valid_0_delay_16_3 <= io_A_Valid_0_delay_15_4;
    io_A_Valid_0_delay_17_2 <= io_A_Valid_0_delay_16_3;
    io_A_Valid_0_delay_18_1 <= io_A_Valid_0_delay_17_2;
    io_A_Valid_0_delay_19 <= io_A_Valid_0_delay_18_1;
    io_A_Valid_0_delay_1_19 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_18 <= io_A_Valid_0_delay_1_19;
    io_A_Valid_0_delay_3_17 <= io_A_Valid_0_delay_2_18;
    io_A_Valid_0_delay_4_16 <= io_A_Valid_0_delay_3_17;
    io_A_Valid_0_delay_5_15 <= io_A_Valid_0_delay_4_16;
    io_A_Valid_0_delay_6_14 <= io_A_Valid_0_delay_5_15;
    io_A_Valid_0_delay_7_13 <= io_A_Valid_0_delay_6_14;
    io_A_Valid_0_delay_8_12 <= io_A_Valid_0_delay_7_13;
    io_A_Valid_0_delay_9_11 <= io_A_Valid_0_delay_8_12;
    io_A_Valid_0_delay_10_10 <= io_A_Valid_0_delay_9_11;
    io_A_Valid_0_delay_11_9 <= io_A_Valid_0_delay_10_10;
    io_A_Valid_0_delay_12_8 <= io_A_Valid_0_delay_11_9;
    io_A_Valid_0_delay_13_7 <= io_A_Valid_0_delay_12_8;
    io_A_Valid_0_delay_14_6 <= io_A_Valid_0_delay_13_7;
    io_A_Valid_0_delay_15_5 <= io_A_Valid_0_delay_14_6;
    io_A_Valid_0_delay_16_4 <= io_A_Valid_0_delay_15_5;
    io_A_Valid_0_delay_17_3 <= io_A_Valid_0_delay_16_4;
    io_A_Valid_0_delay_18_2 <= io_A_Valid_0_delay_17_3;
    io_A_Valid_0_delay_19_1 <= io_A_Valid_0_delay_18_2;
    io_A_Valid_0_delay_20 <= io_A_Valid_0_delay_19_1;
    io_A_Valid_0_delay_1_20 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_19 <= io_A_Valid_0_delay_1_20;
    io_A_Valid_0_delay_3_18 <= io_A_Valid_0_delay_2_19;
    io_A_Valid_0_delay_4_17 <= io_A_Valid_0_delay_3_18;
    io_A_Valid_0_delay_5_16 <= io_A_Valid_0_delay_4_17;
    io_A_Valid_0_delay_6_15 <= io_A_Valid_0_delay_5_16;
    io_A_Valid_0_delay_7_14 <= io_A_Valid_0_delay_6_15;
    io_A_Valid_0_delay_8_13 <= io_A_Valid_0_delay_7_14;
    io_A_Valid_0_delay_9_12 <= io_A_Valid_0_delay_8_13;
    io_A_Valid_0_delay_10_11 <= io_A_Valid_0_delay_9_12;
    io_A_Valid_0_delay_11_10 <= io_A_Valid_0_delay_10_11;
    io_A_Valid_0_delay_12_9 <= io_A_Valid_0_delay_11_10;
    io_A_Valid_0_delay_13_8 <= io_A_Valid_0_delay_12_9;
    io_A_Valid_0_delay_14_7 <= io_A_Valid_0_delay_13_8;
    io_A_Valid_0_delay_15_6 <= io_A_Valid_0_delay_14_7;
    io_A_Valid_0_delay_16_5 <= io_A_Valid_0_delay_15_6;
    io_A_Valid_0_delay_17_4 <= io_A_Valid_0_delay_16_5;
    io_A_Valid_0_delay_18_3 <= io_A_Valid_0_delay_17_4;
    io_A_Valid_0_delay_19_2 <= io_A_Valid_0_delay_18_3;
    io_A_Valid_0_delay_20_1 <= io_A_Valid_0_delay_19_2;
    io_A_Valid_0_delay_21 <= io_A_Valid_0_delay_20_1;
    io_A_Valid_0_delay_1_21 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_20 <= io_A_Valid_0_delay_1_21;
    io_A_Valid_0_delay_3_19 <= io_A_Valid_0_delay_2_20;
    io_A_Valid_0_delay_4_18 <= io_A_Valid_0_delay_3_19;
    io_A_Valid_0_delay_5_17 <= io_A_Valid_0_delay_4_18;
    io_A_Valid_0_delay_6_16 <= io_A_Valid_0_delay_5_17;
    io_A_Valid_0_delay_7_15 <= io_A_Valid_0_delay_6_16;
    io_A_Valid_0_delay_8_14 <= io_A_Valid_0_delay_7_15;
    io_A_Valid_0_delay_9_13 <= io_A_Valid_0_delay_8_14;
    io_A_Valid_0_delay_10_12 <= io_A_Valid_0_delay_9_13;
    io_A_Valid_0_delay_11_11 <= io_A_Valid_0_delay_10_12;
    io_A_Valid_0_delay_12_10 <= io_A_Valid_0_delay_11_11;
    io_A_Valid_0_delay_13_9 <= io_A_Valid_0_delay_12_10;
    io_A_Valid_0_delay_14_8 <= io_A_Valid_0_delay_13_9;
    io_A_Valid_0_delay_15_7 <= io_A_Valid_0_delay_14_8;
    io_A_Valid_0_delay_16_6 <= io_A_Valid_0_delay_15_7;
    io_A_Valid_0_delay_17_5 <= io_A_Valid_0_delay_16_6;
    io_A_Valid_0_delay_18_4 <= io_A_Valid_0_delay_17_5;
    io_A_Valid_0_delay_19_3 <= io_A_Valid_0_delay_18_4;
    io_A_Valid_0_delay_20_2 <= io_A_Valid_0_delay_19_3;
    io_A_Valid_0_delay_21_1 <= io_A_Valid_0_delay_20_2;
    io_A_Valid_0_delay_22 <= io_A_Valid_0_delay_21_1;
    io_A_Valid_0_delay_1_22 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_21 <= io_A_Valid_0_delay_1_22;
    io_A_Valid_0_delay_3_20 <= io_A_Valid_0_delay_2_21;
    io_A_Valid_0_delay_4_19 <= io_A_Valid_0_delay_3_20;
    io_A_Valid_0_delay_5_18 <= io_A_Valid_0_delay_4_19;
    io_A_Valid_0_delay_6_17 <= io_A_Valid_0_delay_5_18;
    io_A_Valid_0_delay_7_16 <= io_A_Valid_0_delay_6_17;
    io_A_Valid_0_delay_8_15 <= io_A_Valid_0_delay_7_16;
    io_A_Valid_0_delay_9_14 <= io_A_Valid_0_delay_8_15;
    io_A_Valid_0_delay_10_13 <= io_A_Valid_0_delay_9_14;
    io_A_Valid_0_delay_11_12 <= io_A_Valid_0_delay_10_13;
    io_A_Valid_0_delay_12_11 <= io_A_Valid_0_delay_11_12;
    io_A_Valid_0_delay_13_10 <= io_A_Valid_0_delay_12_11;
    io_A_Valid_0_delay_14_9 <= io_A_Valid_0_delay_13_10;
    io_A_Valid_0_delay_15_8 <= io_A_Valid_0_delay_14_9;
    io_A_Valid_0_delay_16_7 <= io_A_Valid_0_delay_15_8;
    io_A_Valid_0_delay_17_6 <= io_A_Valid_0_delay_16_7;
    io_A_Valid_0_delay_18_5 <= io_A_Valid_0_delay_17_6;
    io_A_Valid_0_delay_19_4 <= io_A_Valid_0_delay_18_5;
    io_A_Valid_0_delay_20_3 <= io_A_Valid_0_delay_19_4;
    io_A_Valid_0_delay_21_2 <= io_A_Valid_0_delay_20_3;
    io_A_Valid_0_delay_22_1 <= io_A_Valid_0_delay_21_2;
    io_A_Valid_0_delay_23 <= io_A_Valid_0_delay_22_1;
    io_A_Valid_0_delay_1_23 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_22 <= io_A_Valid_0_delay_1_23;
    io_A_Valid_0_delay_3_21 <= io_A_Valid_0_delay_2_22;
    io_A_Valid_0_delay_4_20 <= io_A_Valid_0_delay_3_21;
    io_A_Valid_0_delay_5_19 <= io_A_Valid_0_delay_4_20;
    io_A_Valid_0_delay_6_18 <= io_A_Valid_0_delay_5_19;
    io_A_Valid_0_delay_7_17 <= io_A_Valid_0_delay_6_18;
    io_A_Valid_0_delay_8_16 <= io_A_Valid_0_delay_7_17;
    io_A_Valid_0_delay_9_15 <= io_A_Valid_0_delay_8_16;
    io_A_Valid_0_delay_10_14 <= io_A_Valid_0_delay_9_15;
    io_A_Valid_0_delay_11_13 <= io_A_Valid_0_delay_10_14;
    io_A_Valid_0_delay_12_12 <= io_A_Valid_0_delay_11_13;
    io_A_Valid_0_delay_13_11 <= io_A_Valid_0_delay_12_12;
    io_A_Valid_0_delay_14_10 <= io_A_Valid_0_delay_13_11;
    io_A_Valid_0_delay_15_9 <= io_A_Valid_0_delay_14_10;
    io_A_Valid_0_delay_16_8 <= io_A_Valid_0_delay_15_9;
    io_A_Valid_0_delay_17_7 <= io_A_Valid_0_delay_16_8;
    io_A_Valid_0_delay_18_6 <= io_A_Valid_0_delay_17_7;
    io_A_Valid_0_delay_19_5 <= io_A_Valid_0_delay_18_6;
    io_A_Valid_0_delay_20_4 <= io_A_Valid_0_delay_19_5;
    io_A_Valid_0_delay_21_3 <= io_A_Valid_0_delay_20_4;
    io_A_Valid_0_delay_22_2 <= io_A_Valid_0_delay_21_3;
    io_A_Valid_0_delay_23_1 <= io_A_Valid_0_delay_22_2;
    io_A_Valid_0_delay_24 <= io_A_Valid_0_delay_23_1;
    io_A_Valid_0_delay_1_24 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_23 <= io_A_Valid_0_delay_1_24;
    io_A_Valid_0_delay_3_22 <= io_A_Valid_0_delay_2_23;
    io_A_Valid_0_delay_4_21 <= io_A_Valid_0_delay_3_22;
    io_A_Valid_0_delay_5_20 <= io_A_Valid_0_delay_4_21;
    io_A_Valid_0_delay_6_19 <= io_A_Valid_0_delay_5_20;
    io_A_Valid_0_delay_7_18 <= io_A_Valid_0_delay_6_19;
    io_A_Valid_0_delay_8_17 <= io_A_Valid_0_delay_7_18;
    io_A_Valid_0_delay_9_16 <= io_A_Valid_0_delay_8_17;
    io_A_Valid_0_delay_10_15 <= io_A_Valid_0_delay_9_16;
    io_A_Valid_0_delay_11_14 <= io_A_Valid_0_delay_10_15;
    io_A_Valid_0_delay_12_13 <= io_A_Valid_0_delay_11_14;
    io_A_Valid_0_delay_13_12 <= io_A_Valid_0_delay_12_13;
    io_A_Valid_0_delay_14_11 <= io_A_Valid_0_delay_13_12;
    io_A_Valid_0_delay_15_10 <= io_A_Valid_0_delay_14_11;
    io_A_Valid_0_delay_16_9 <= io_A_Valid_0_delay_15_10;
    io_A_Valid_0_delay_17_8 <= io_A_Valid_0_delay_16_9;
    io_A_Valid_0_delay_18_7 <= io_A_Valid_0_delay_17_8;
    io_A_Valid_0_delay_19_6 <= io_A_Valid_0_delay_18_7;
    io_A_Valid_0_delay_20_5 <= io_A_Valid_0_delay_19_6;
    io_A_Valid_0_delay_21_4 <= io_A_Valid_0_delay_20_5;
    io_A_Valid_0_delay_22_3 <= io_A_Valid_0_delay_21_4;
    io_A_Valid_0_delay_23_2 <= io_A_Valid_0_delay_22_3;
    io_A_Valid_0_delay_24_1 <= io_A_Valid_0_delay_23_2;
    io_A_Valid_0_delay_25 <= io_A_Valid_0_delay_24_1;
    io_A_Valid_0_delay_1_25 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_24 <= io_A_Valid_0_delay_1_25;
    io_A_Valid_0_delay_3_23 <= io_A_Valid_0_delay_2_24;
    io_A_Valid_0_delay_4_22 <= io_A_Valid_0_delay_3_23;
    io_A_Valid_0_delay_5_21 <= io_A_Valid_0_delay_4_22;
    io_A_Valid_0_delay_6_20 <= io_A_Valid_0_delay_5_21;
    io_A_Valid_0_delay_7_19 <= io_A_Valid_0_delay_6_20;
    io_A_Valid_0_delay_8_18 <= io_A_Valid_0_delay_7_19;
    io_A_Valid_0_delay_9_17 <= io_A_Valid_0_delay_8_18;
    io_A_Valid_0_delay_10_16 <= io_A_Valid_0_delay_9_17;
    io_A_Valid_0_delay_11_15 <= io_A_Valid_0_delay_10_16;
    io_A_Valid_0_delay_12_14 <= io_A_Valid_0_delay_11_15;
    io_A_Valid_0_delay_13_13 <= io_A_Valid_0_delay_12_14;
    io_A_Valid_0_delay_14_12 <= io_A_Valid_0_delay_13_13;
    io_A_Valid_0_delay_15_11 <= io_A_Valid_0_delay_14_12;
    io_A_Valid_0_delay_16_10 <= io_A_Valid_0_delay_15_11;
    io_A_Valid_0_delay_17_9 <= io_A_Valid_0_delay_16_10;
    io_A_Valid_0_delay_18_8 <= io_A_Valid_0_delay_17_9;
    io_A_Valid_0_delay_19_7 <= io_A_Valid_0_delay_18_8;
    io_A_Valid_0_delay_20_6 <= io_A_Valid_0_delay_19_7;
    io_A_Valid_0_delay_21_5 <= io_A_Valid_0_delay_20_6;
    io_A_Valid_0_delay_22_4 <= io_A_Valid_0_delay_21_5;
    io_A_Valid_0_delay_23_3 <= io_A_Valid_0_delay_22_4;
    io_A_Valid_0_delay_24_2 <= io_A_Valid_0_delay_23_3;
    io_A_Valid_0_delay_25_1 <= io_A_Valid_0_delay_24_2;
    io_A_Valid_0_delay_26 <= io_A_Valid_0_delay_25_1;
    io_A_Valid_0_delay_1_26 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_25 <= io_A_Valid_0_delay_1_26;
    io_A_Valid_0_delay_3_24 <= io_A_Valid_0_delay_2_25;
    io_A_Valid_0_delay_4_23 <= io_A_Valid_0_delay_3_24;
    io_A_Valid_0_delay_5_22 <= io_A_Valid_0_delay_4_23;
    io_A_Valid_0_delay_6_21 <= io_A_Valid_0_delay_5_22;
    io_A_Valid_0_delay_7_20 <= io_A_Valid_0_delay_6_21;
    io_A_Valid_0_delay_8_19 <= io_A_Valid_0_delay_7_20;
    io_A_Valid_0_delay_9_18 <= io_A_Valid_0_delay_8_19;
    io_A_Valid_0_delay_10_17 <= io_A_Valid_0_delay_9_18;
    io_A_Valid_0_delay_11_16 <= io_A_Valid_0_delay_10_17;
    io_A_Valid_0_delay_12_15 <= io_A_Valid_0_delay_11_16;
    io_A_Valid_0_delay_13_14 <= io_A_Valid_0_delay_12_15;
    io_A_Valid_0_delay_14_13 <= io_A_Valid_0_delay_13_14;
    io_A_Valid_0_delay_15_12 <= io_A_Valid_0_delay_14_13;
    io_A_Valid_0_delay_16_11 <= io_A_Valid_0_delay_15_12;
    io_A_Valid_0_delay_17_10 <= io_A_Valid_0_delay_16_11;
    io_A_Valid_0_delay_18_9 <= io_A_Valid_0_delay_17_10;
    io_A_Valid_0_delay_19_8 <= io_A_Valid_0_delay_18_9;
    io_A_Valid_0_delay_20_7 <= io_A_Valid_0_delay_19_8;
    io_A_Valid_0_delay_21_6 <= io_A_Valid_0_delay_20_7;
    io_A_Valid_0_delay_22_5 <= io_A_Valid_0_delay_21_6;
    io_A_Valid_0_delay_23_4 <= io_A_Valid_0_delay_22_5;
    io_A_Valid_0_delay_24_3 <= io_A_Valid_0_delay_23_4;
    io_A_Valid_0_delay_25_2 <= io_A_Valid_0_delay_24_3;
    io_A_Valid_0_delay_26_1 <= io_A_Valid_0_delay_25_2;
    io_A_Valid_0_delay_27 <= io_A_Valid_0_delay_26_1;
    io_A_Valid_0_delay_1_27 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_26 <= io_A_Valid_0_delay_1_27;
    io_A_Valid_0_delay_3_25 <= io_A_Valid_0_delay_2_26;
    io_A_Valid_0_delay_4_24 <= io_A_Valid_0_delay_3_25;
    io_A_Valid_0_delay_5_23 <= io_A_Valid_0_delay_4_24;
    io_A_Valid_0_delay_6_22 <= io_A_Valid_0_delay_5_23;
    io_A_Valid_0_delay_7_21 <= io_A_Valid_0_delay_6_22;
    io_A_Valid_0_delay_8_20 <= io_A_Valid_0_delay_7_21;
    io_A_Valid_0_delay_9_19 <= io_A_Valid_0_delay_8_20;
    io_A_Valid_0_delay_10_18 <= io_A_Valid_0_delay_9_19;
    io_A_Valid_0_delay_11_17 <= io_A_Valid_0_delay_10_18;
    io_A_Valid_0_delay_12_16 <= io_A_Valid_0_delay_11_17;
    io_A_Valid_0_delay_13_15 <= io_A_Valid_0_delay_12_16;
    io_A_Valid_0_delay_14_14 <= io_A_Valid_0_delay_13_15;
    io_A_Valid_0_delay_15_13 <= io_A_Valid_0_delay_14_14;
    io_A_Valid_0_delay_16_12 <= io_A_Valid_0_delay_15_13;
    io_A_Valid_0_delay_17_11 <= io_A_Valid_0_delay_16_12;
    io_A_Valid_0_delay_18_10 <= io_A_Valid_0_delay_17_11;
    io_A_Valid_0_delay_19_9 <= io_A_Valid_0_delay_18_10;
    io_A_Valid_0_delay_20_8 <= io_A_Valid_0_delay_19_9;
    io_A_Valid_0_delay_21_7 <= io_A_Valid_0_delay_20_8;
    io_A_Valid_0_delay_22_6 <= io_A_Valid_0_delay_21_7;
    io_A_Valid_0_delay_23_5 <= io_A_Valid_0_delay_22_6;
    io_A_Valid_0_delay_24_4 <= io_A_Valid_0_delay_23_5;
    io_A_Valid_0_delay_25_3 <= io_A_Valid_0_delay_24_4;
    io_A_Valid_0_delay_26_2 <= io_A_Valid_0_delay_25_3;
    io_A_Valid_0_delay_27_1 <= io_A_Valid_0_delay_26_2;
    io_A_Valid_0_delay_28 <= io_A_Valid_0_delay_27_1;
    io_A_Valid_0_delay_1_28 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_27 <= io_A_Valid_0_delay_1_28;
    io_A_Valid_0_delay_3_26 <= io_A_Valid_0_delay_2_27;
    io_A_Valid_0_delay_4_25 <= io_A_Valid_0_delay_3_26;
    io_A_Valid_0_delay_5_24 <= io_A_Valid_0_delay_4_25;
    io_A_Valid_0_delay_6_23 <= io_A_Valid_0_delay_5_24;
    io_A_Valid_0_delay_7_22 <= io_A_Valid_0_delay_6_23;
    io_A_Valid_0_delay_8_21 <= io_A_Valid_0_delay_7_22;
    io_A_Valid_0_delay_9_20 <= io_A_Valid_0_delay_8_21;
    io_A_Valid_0_delay_10_19 <= io_A_Valid_0_delay_9_20;
    io_A_Valid_0_delay_11_18 <= io_A_Valid_0_delay_10_19;
    io_A_Valid_0_delay_12_17 <= io_A_Valid_0_delay_11_18;
    io_A_Valid_0_delay_13_16 <= io_A_Valid_0_delay_12_17;
    io_A_Valid_0_delay_14_15 <= io_A_Valid_0_delay_13_16;
    io_A_Valid_0_delay_15_14 <= io_A_Valid_0_delay_14_15;
    io_A_Valid_0_delay_16_13 <= io_A_Valid_0_delay_15_14;
    io_A_Valid_0_delay_17_12 <= io_A_Valid_0_delay_16_13;
    io_A_Valid_0_delay_18_11 <= io_A_Valid_0_delay_17_12;
    io_A_Valid_0_delay_19_10 <= io_A_Valid_0_delay_18_11;
    io_A_Valid_0_delay_20_9 <= io_A_Valid_0_delay_19_10;
    io_A_Valid_0_delay_21_8 <= io_A_Valid_0_delay_20_9;
    io_A_Valid_0_delay_22_7 <= io_A_Valid_0_delay_21_8;
    io_A_Valid_0_delay_23_6 <= io_A_Valid_0_delay_22_7;
    io_A_Valid_0_delay_24_5 <= io_A_Valid_0_delay_23_6;
    io_A_Valid_0_delay_25_4 <= io_A_Valid_0_delay_24_5;
    io_A_Valid_0_delay_26_3 <= io_A_Valid_0_delay_25_4;
    io_A_Valid_0_delay_27_2 <= io_A_Valid_0_delay_26_3;
    io_A_Valid_0_delay_28_1 <= io_A_Valid_0_delay_27_2;
    io_A_Valid_0_delay_29 <= io_A_Valid_0_delay_28_1;
    io_A_Valid_0_delay_1_29 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_28 <= io_A_Valid_0_delay_1_29;
    io_A_Valid_0_delay_3_27 <= io_A_Valid_0_delay_2_28;
    io_A_Valid_0_delay_4_26 <= io_A_Valid_0_delay_3_27;
    io_A_Valid_0_delay_5_25 <= io_A_Valid_0_delay_4_26;
    io_A_Valid_0_delay_6_24 <= io_A_Valid_0_delay_5_25;
    io_A_Valid_0_delay_7_23 <= io_A_Valid_0_delay_6_24;
    io_A_Valid_0_delay_8_22 <= io_A_Valid_0_delay_7_23;
    io_A_Valid_0_delay_9_21 <= io_A_Valid_0_delay_8_22;
    io_A_Valid_0_delay_10_20 <= io_A_Valid_0_delay_9_21;
    io_A_Valid_0_delay_11_19 <= io_A_Valid_0_delay_10_20;
    io_A_Valid_0_delay_12_18 <= io_A_Valid_0_delay_11_19;
    io_A_Valid_0_delay_13_17 <= io_A_Valid_0_delay_12_18;
    io_A_Valid_0_delay_14_16 <= io_A_Valid_0_delay_13_17;
    io_A_Valid_0_delay_15_15 <= io_A_Valid_0_delay_14_16;
    io_A_Valid_0_delay_16_14 <= io_A_Valid_0_delay_15_15;
    io_A_Valid_0_delay_17_13 <= io_A_Valid_0_delay_16_14;
    io_A_Valid_0_delay_18_12 <= io_A_Valid_0_delay_17_13;
    io_A_Valid_0_delay_19_11 <= io_A_Valid_0_delay_18_12;
    io_A_Valid_0_delay_20_10 <= io_A_Valid_0_delay_19_11;
    io_A_Valid_0_delay_21_9 <= io_A_Valid_0_delay_20_10;
    io_A_Valid_0_delay_22_8 <= io_A_Valid_0_delay_21_9;
    io_A_Valid_0_delay_23_7 <= io_A_Valid_0_delay_22_8;
    io_A_Valid_0_delay_24_6 <= io_A_Valid_0_delay_23_7;
    io_A_Valid_0_delay_25_5 <= io_A_Valid_0_delay_24_6;
    io_A_Valid_0_delay_26_4 <= io_A_Valid_0_delay_25_5;
    io_A_Valid_0_delay_27_3 <= io_A_Valid_0_delay_26_4;
    io_A_Valid_0_delay_28_2 <= io_A_Valid_0_delay_27_3;
    io_A_Valid_0_delay_29_1 <= io_A_Valid_0_delay_28_2;
    io_A_Valid_0_delay_30 <= io_A_Valid_0_delay_29_1;
    io_A_Valid_0_delay_1_30 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_29 <= io_A_Valid_0_delay_1_30;
    io_A_Valid_0_delay_3_28 <= io_A_Valid_0_delay_2_29;
    io_A_Valid_0_delay_4_27 <= io_A_Valid_0_delay_3_28;
    io_A_Valid_0_delay_5_26 <= io_A_Valid_0_delay_4_27;
    io_A_Valid_0_delay_6_25 <= io_A_Valid_0_delay_5_26;
    io_A_Valid_0_delay_7_24 <= io_A_Valid_0_delay_6_25;
    io_A_Valid_0_delay_8_23 <= io_A_Valid_0_delay_7_24;
    io_A_Valid_0_delay_9_22 <= io_A_Valid_0_delay_8_23;
    io_A_Valid_0_delay_10_21 <= io_A_Valid_0_delay_9_22;
    io_A_Valid_0_delay_11_20 <= io_A_Valid_0_delay_10_21;
    io_A_Valid_0_delay_12_19 <= io_A_Valid_0_delay_11_20;
    io_A_Valid_0_delay_13_18 <= io_A_Valid_0_delay_12_19;
    io_A_Valid_0_delay_14_17 <= io_A_Valid_0_delay_13_18;
    io_A_Valid_0_delay_15_16 <= io_A_Valid_0_delay_14_17;
    io_A_Valid_0_delay_16_15 <= io_A_Valid_0_delay_15_16;
    io_A_Valid_0_delay_17_14 <= io_A_Valid_0_delay_16_15;
    io_A_Valid_0_delay_18_13 <= io_A_Valid_0_delay_17_14;
    io_A_Valid_0_delay_19_12 <= io_A_Valid_0_delay_18_13;
    io_A_Valid_0_delay_20_11 <= io_A_Valid_0_delay_19_12;
    io_A_Valid_0_delay_21_10 <= io_A_Valid_0_delay_20_11;
    io_A_Valid_0_delay_22_9 <= io_A_Valid_0_delay_21_10;
    io_A_Valid_0_delay_23_8 <= io_A_Valid_0_delay_22_9;
    io_A_Valid_0_delay_24_7 <= io_A_Valid_0_delay_23_8;
    io_A_Valid_0_delay_25_6 <= io_A_Valid_0_delay_24_7;
    io_A_Valid_0_delay_26_5 <= io_A_Valid_0_delay_25_6;
    io_A_Valid_0_delay_27_4 <= io_A_Valid_0_delay_26_5;
    io_A_Valid_0_delay_28_3 <= io_A_Valid_0_delay_27_4;
    io_A_Valid_0_delay_29_2 <= io_A_Valid_0_delay_28_3;
    io_A_Valid_0_delay_30_1 <= io_A_Valid_0_delay_29_2;
    io_A_Valid_0_delay_31 <= io_A_Valid_0_delay_30_1;
    io_A_Valid_0_delay_1_31 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_30 <= io_A_Valid_0_delay_1_31;
    io_A_Valid_0_delay_3_29 <= io_A_Valid_0_delay_2_30;
    io_A_Valid_0_delay_4_28 <= io_A_Valid_0_delay_3_29;
    io_A_Valid_0_delay_5_27 <= io_A_Valid_0_delay_4_28;
    io_A_Valid_0_delay_6_26 <= io_A_Valid_0_delay_5_27;
    io_A_Valid_0_delay_7_25 <= io_A_Valid_0_delay_6_26;
    io_A_Valid_0_delay_8_24 <= io_A_Valid_0_delay_7_25;
    io_A_Valid_0_delay_9_23 <= io_A_Valid_0_delay_8_24;
    io_A_Valid_0_delay_10_22 <= io_A_Valid_0_delay_9_23;
    io_A_Valid_0_delay_11_21 <= io_A_Valid_0_delay_10_22;
    io_A_Valid_0_delay_12_20 <= io_A_Valid_0_delay_11_21;
    io_A_Valid_0_delay_13_19 <= io_A_Valid_0_delay_12_20;
    io_A_Valid_0_delay_14_18 <= io_A_Valid_0_delay_13_19;
    io_A_Valid_0_delay_15_17 <= io_A_Valid_0_delay_14_18;
    io_A_Valid_0_delay_16_16 <= io_A_Valid_0_delay_15_17;
    io_A_Valid_0_delay_17_15 <= io_A_Valid_0_delay_16_16;
    io_A_Valid_0_delay_18_14 <= io_A_Valid_0_delay_17_15;
    io_A_Valid_0_delay_19_13 <= io_A_Valid_0_delay_18_14;
    io_A_Valid_0_delay_20_12 <= io_A_Valid_0_delay_19_13;
    io_A_Valid_0_delay_21_11 <= io_A_Valid_0_delay_20_12;
    io_A_Valid_0_delay_22_10 <= io_A_Valid_0_delay_21_11;
    io_A_Valid_0_delay_23_9 <= io_A_Valid_0_delay_22_10;
    io_A_Valid_0_delay_24_8 <= io_A_Valid_0_delay_23_9;
    io_A_Valid_0_delay_25_7 <= io_A_Valid_0_delay_24_8;
    io_A_Valid_0_delay_26_6 <= io_A_Valid_0_delay_25_7;
    io_A_Valid_0_delay_27_5 <= io_A_Valid_0_delay_26_6;
    io_A_Valid_0_delay_28_4 <= io_A_Valid_0_delay_27_5;
    io_A_Valid_0_delay_29_3 <= io_A_Valid_0_delay_28_4;
    io_A_Valid_0_delay_30_2 <= io_A_Valid_0_delay_29_3;
    io_A_Valid_0_delay_31_1 <= io_A_Valid_0_delay_30_2;
    io_A_Valid_0_delay_32 <= io_A_Valid_0_delay_31_1;
    io_A_Valid_0_delay_1_32 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_31 <= io_A_Valid_0_delay_1_32;
    io_A_Valid_0_delay_3_30 <= io_A_Valid_0_delay_2_31;
    io_A_Valid_0_delay_4_29 <= io_A_Valid_0_delay_3_30;
    io_A_Valid_0_delay_5_28 <= io_A_Valid_0_delay_4_29;
    io_A_Valid_0_delay_6_27 <= io_A_Valid_0_delay_5_28;
    io_A_Valid_0_delay_7_26 <= io_A_Valid_0_delay_6_27;
    io_A_Valid_0_delay_8_25 <= io_A_Valid_0_delay_7_26;
    io_A_Valid_0_delay_9_24 <= io_A_Valid_0_delay_8_25;
    io_A_Valid_0_delay_10_23 <= io_A_Valid_0_delay_9_24;
    io_A_Valid_0_delay_11_22 <= io_A_Valid_0_delay_10_23;
    io_A_Valid_0_delay_12_21 <= io_A_Valid_0_delay_11_22;
    io_A_Valid_0_delay_13_20 <= io_A_Valid_0_delay_12_21;
    io_A_Valid_0_delay_14_19 <= io_A_Valid_0_delay_13_20;
    io_A_Valid_0_delay_15_18 <= io_A_Valid_0_delay_14_19;
    io_A_Valid_0_delay_16_17 <= io_A_Valid_0_delay_15_18;
    io_A_Valid_0_delay_17_16 <= io_A_Valid_0_delay_16_17;
    io_A_Valid_0_delay_18_15 <= io_A_Valid_0_delay_17_16;
    io_A_Valid_0_delay_19_14 <= io_A_Valid_0_delay_18_15;
    io_A_Valid_0_delay_20_13 <= io_A_Valid_0_delay_19_14;
    io_A_Valid_0_delay_21_12 <= io_A_Valid_0_delay_20_13;
    io_A_Valid_0_delay_22_11 <= io_A_Valid_0_delay_21_12;
    io_A_Valid_0_delay_23_10 <= io_A_Valid_0_delay_22_11;
    io_A_Valid_0_delay_24_9 <= io_A_Valid_0_delay_23_10;
    io_A_Valid_0_delay_25_8 <= io_A_Valid_0_delay_24_9;
    io_A_Valid_0_delay_26_7 <= io_A_Valid_0_delay_25_8;
    io_A_Valid_0_delay_27_6 <= io_A_Valid_0_delay_26_7;
    io_A_Valid_0_delay_28_5 <= io_A_Valid_0_delay_27_6;
    io_A_Valid_0_delay_29_4 <= io_A_Valid_0_delay_28_5;
    io_A_Valid_0_delay_30_3 <= io_A_Valid_0_delay_29_4;
    io_A_Valid_0_delay_31_2 <= io_A_Valid_0_delay_30_3;
    io_A_Valid_0_delay_32_1 <= io_A_Valid_0_delay_31_2;
    io_A_Valid_0_delay_33 <= io_A_Valid_0_delay_32_1;
    io_A_Valid_0_delay_1_33 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_32 <= io_A_Valid_0_delay_1_33;
    io_A_Valid_0_delay_3_31 <= io_A_Valid_0_delay_2_32;
    io_A_Valid_0_delay_4_30 <= io_A_Valid_0_delay_3_31;
    io_A_Valid_0_delay_5_29 <= io_A_Valid_0_delay_4_30;
    io_A_Valid_0_delay_6_28 <= io_A_Valid_0_delay_5_29;
    io_A_Valid_0_delay_7_27 <= io_A_Valid_0_delay_6_28;
    io_A_Valid_0_delay_8_26 <= io_A_Valid_0_delay_7_27;
    io_A_Valid_0_delay_9_25 <= io_A_Valid_0_delay_8_26;
    io_A_Valid_0_delay_10_24 <= io_A_Valid_0_delay_9_25;
    io_A_Valid_0_delay_11_23 <= io_A_Valid_0_delay_10_24;
    io_A_Valid_0_delay_12_22 <= io_A_Valid_0_delay_11_23;
    io_A_Valid_0_delay_13_21 <= io_A_Valid_0_delay_12_22;
    io_A_Valid_0_delay_14_20 <= io_A_Valid_0_delay_13_21;
    io_A_Valid_0_delay_15_19 <= io_A_Valid_0_delay_14_20;
    io_A_Valid_0_delay_16_18 <= io_A_Valid_0_delay_15_19;
    io_A_Valid_0_delay_17_17 <= io_A_Valid_0_delay_16_18;
    io_A_Valid_0_delay_18_16 <= io_A_Valid_0_delay_17_17;
    io_A_Valid_0_delay_19_15 <= io_A_Valid_0_delay_18_16;
    io_A_Valid_0_delay_20_14 <= io_A_Valid_0_delay_19_15;
    io_A_Valid_0_delay_21_13 <= io_A_Valid_0_delay_20_14;
    io_A_Valid_0_delay_22_12 <= io_A_Valid_0_delay_21_13;
    io_A_Valid_0_delay_23_11 <= io_A_Valid_0_delay_22_12;
    io_A_Valid_0_delay_24_10 <= io_A_Valid_0_delay_23_11;
    io_A_Valid_0_delay_25_9 <= io_A_Valid_0_delay_24_10;
    io_A_Valid_0_delay_26_8 <= io_A_Valid_0_delay_25_9;
    io_A_Valid_0_delay_27_7 <= io_A_Valid_0_delay_26_8;
    io_A_Valid_0_delay_28_6 <= io_A_Valid_0_delay_27_7;
    io_A_Valid_0_delay_29_5 <= io_A_Valid_0_delay_28_6;
    io_A_Valid_0_delay_30_4 <= io_A_Valid_0_delay_29_5;
    io_A_Valid_0_delay_31_3 <= io_A_Valid_0_delay_30_4;
    io_A_Valid_0_delay_32_2 <= io_A_Valid_0_delay_31_3;
    io_A_Valid_0_delay_33_1 <= io_A_Valid_0_delay_32_2;
    io_A_Valid_0_delay_34 <= io_A_Valid_0_delay_33_1;
    io_A_Valid_0_delay_1_34 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_33 <= io_A_Valid_0_delay_1_34;
    io_A_Valid_0_delay_3_32 <= io_A_Valid_0_delay_2_33;
    io_A_Valid_0_delay_4_31 <= io_A_Valid_0_delay_3_32;
    io_A_Valid_0_delay_5_30 <= io_A_Valid_0_delay_4_31;
    io_A_Valid_0_delay_6_29 <= io_A_Valid_0_delay_5_30;
    io_A_Valid_0_delay_7_28 <= io_A_Valid_0_delay_6_29;
    io_A_Valid_0_delay_8_27 <= io_A_Valid_0_delay_7_28;
    io_A_Valid_0_delay_9_26 <= io_A_Valid_0_delay_8_27;
    io_A_Valid_0_delay_10_25 <= io_A_Valid_0_delay_9_26;
    io_A_Valid_0_delay_11_24 <= io_A_Valid_0_delay_10_25;
    io_A_Valid_0_delay_12_23 <= io_A_Valid_0_delay_11_24;
    io_A_Valid_0_delay_13_22 <= io_A_Valid_0_delay_12_23;
    io_A_Valid_0_delay_14_21 <= io_A_Valid_0_delay_13_22;
    io_A_Valid_0_delay_15_20 <= io_A_Valid_0_delay_14_21;
    io_A_Valid_0_delay_16_19 <= io_A_Valid_0_delay_15_20;
    io_A_Valid_0_delay_17_18 <= io_A_Valid_0_delay_16_19;
    io_A_Valid_0_delay_18_17 <= io_A_Valid_0_delay_17_18;
    io_A_Valid_0_delay_19_16 <= io_A_Valid_0_delay_18_17;
    io_A_Valid_0_delay_20_15 <= io_A_Valid_0_delay_19_16;
    io_A_Valid_0_delay_21_14 <= io_A_Valid_0_delay_20_15;
    io_A_Valid_0_delay_22_13 <= io_A_Valid_0_delay_21_14;
    io_A_Valid_0_delay_23_12 <= io_A_Valid_0_delay_22_13;
    io_A_Valid_0_delay_24_11 <= io_A_Valid_0_delay_23_12;
    io_A_Valid_0_delay_25_10 <= io_A_Valid_0_delay_24_11;
    io_A_Valid_0_delay_26_9 <= io_A_Valid_0_delay_25_10;
    io_A_Valid_0_delay_27_8 <= io_A_Valid_0_delay_26_9;
    io_A_Valid_0_delay_28_7 <= io_A_Valid_0_delay_27_8;
    io_A_Valid_0_delay_29_6 <= io_A_Valid_0_delay_28_7;
    io_A_Valid_0_delay_30_5 <= io_A_Valid_0_delay_29_6;
    io_A_Valid_0_delay_31_4 <= io_A_Valid_0_delay_30_5;
    io_A_Valid_0_delay_32_3 <= io_A_Valid_0_delay_31_4;
    io_A_Valid_0_delay_33_2 <= io_A_Valid_0_delay_32_3;
    io_A_Valid_0_delay_34_1 <= io_A_Valid_0_delay_33_2;
    io_A_Valid_0_delay_35 <= io_A_Valid_0_delay_34_1;
    io_A_Valid_0_delay_1_35 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_34 <= io_A_Valid_0_delay_1_35;
    io_A_Valid_0_delay_3_33 <= io_A_Valid_0_delay_2_34;
    io_A_Valid_0_delay_4_32 <= io_A_Valid_0_delay_3_33;
    io_A_Valid_0_delay_5_31 <= io_A_Valid_0_delay_4_32;
    io_A_Valid_0_delay_6_30 <= io_A_Valid_0_delay_5_31;
    io_A_Valid_0_delay_7_29 <= io_A_Valid_0_delay_6_30;
    io_A_Valid_0_delay_8_28 <= io_A_Valid_0_delay_7_29;
    io_A_Valid_0_delay_9_27 <= io_A_Valid_0_delay_8_28;
    io_A_Valid_0_delay_10_26 <= io_A_Valid_0_delay_9_27;
    io_A_Valid_0_delay_11_25 <= io_A_Valid_0_delay_10_26;
    io_A_Valid_0_delay_12_24 <= io_A_Valid_0_delay_11_25;
    io_A_Valid_0_delay_13_23 <= io_A_Valid_0_delay_12_24;
    io_A_Valid_0_delay_14_22 <= io_A_Valid_0_delay_13_23;
    io_A_Valid_0_delay_15_21 <= io_A_Valid_0_delay_14_22;
    io_A_Valid_0_delay_16_20 <= io_A_Valid_0_delay_15_21;
    io_A_Valid_0_delay_17_19 <= io_A_Valid_0_delay_16_20;
    io_A_Valid_0_delay_18_18 <= io_A_Valid_0_delay_17_19;
    io_A_Valid_0_delay_19_17 <= io_A_Valid_0_delay_18_18;
    io_A_Valid_0_delay_20_16 <= io_A_Valid_0_delay_19_17;
    io_A_Valid_0_delay_21_15 <= io_A_Valid_0_delay_20_16;
    io_A_Valid_0_delay_22_14 <= io_A_Valid_0_delay_21_15;
    io_A_Valid_0_delay_23_13 <= io_A_Valid_0_delay_22_14;
    io_A_Valid_0_delay_24_12 <= io_A_Valid_0_delay_23_13;
    io_A_Valid_0_delay_25_11 <= io_A_Valid_0_delay_24_12;
    io_A_Valid_0_delay_26_10 <= io_A_Valid_0_delay_25_11;
    io_A_Valid_0_delay_27_9 <= io_A_Valid_0_delay_26_10;
    io_A_Valid_0_delay_28_8 <= io_A_Valid_0_delay_27_9;
    io_A_Valid_0_delay_29_7 <= io_A_Valid_0_delay_28_8;
    io_A_Valid_0_delay_30_6 <= io_A_Valid_0_delay_29_7;
    io_A_Valid_0_delay_31_5 <= io_A_Valid_0_delay_30_6;
    io_A_Valid_0_delay_32_4 <= io_A_Valid_0_delay_31_5;
    io_A_Valid_0_delay_33_3 <= io_A_Valid_0_delay_32_4;
    io_A_Valid_0_delay_34_2 <= io_A_Valid_0_delay_33_3;
    io_A_Valid_0_delay_35_1 <= io_A_Valid_0_delay_34_2;
    io_A_Valid_0_delay_36 <= io_A_Valid_0_delay_35_1;
    io_A_Valid_0_delay_1_36 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_35 <= io_A_Valid_0_delay_1_36;
    io_A_Valid_0_delay_3_34 <= io_A_Valid_0_delay_2_35;
    io_A_Valid_0_delay_4_33 <= io_A_Valid_0_delay_3_34;
    io_A_Valid_0_delay_5_32 <= io_A_Valid_0_delay_4_33;
    io_A_Valid_0_delay_6_31 <= io_A_Valid_0_delay_5_32;
    io_A_Valid_0_delay_7_30 <= io_A_Valid_0_delay_6_31;
    io_A_Valid_0_delay_8_29 <= io_A_Valid_0_delay_7_30;
    io_A_Valid_0_delay_9_28 <= io_A_Valid_0_delay_8_29;
    io_A_Valid_0_delay_10_27 <= io_A_Valid_0_delay_9_28;
    io_A_Valid_0_delay_11_26 <= io_A_Valid_0_delay_10_27;
    io_A_Valid_0_delay_12_25 <= io_A_Valid_0_delay_11_26;
    io_A_Valid_0_delay_13_24 <= io_A_Valid_0_delay_12_25;
    io_A_Valid_0_delay_14_23 <= io_A_Valid_0_delay_13_24;
    io_A_Valid_0_delay_15_22 <= io_A_Valid_0_delay_14_23;
    io_A_Valid_0_delay_16_21 <= io_A_Valid_0_delay_15_22;
    io_A_Valid_0_delay_17_20 <= io_A_Valid_0_delay_16_21;
    io_A_Valid_0_delay_18_19 <= io_A_Valid_0_delay_17_20;
    io_A_Valid_0_delay_19_18 <= io_A_Valid_0_delay_18_19;
    io_A_Valid_0_delay_20_17 <= io_A_Valid_0_delay_19_18;
    io_A_Valid_0_delay_21_16 <= io_A_Valid_0_delay_20_17;
    io_A_Valid_0_delay_22_15 <= io_A_Valid_0_delay_21_16;
    io_A_Valid_0_delay_23_14 <= io_A_Valid_0_delay_22_15;
    io_A_Valid_0_delay_24_13 <= io_A_Valid_0_delay_23_14;
    io_A_Valid_0_delay_25_12 <= io_A_Valid_0_delay_24_13;
    io_A_Valid_0_delay_26_11 <= io_A_Valid_0_delay_25_12;
    io_A_Valid_0_delay_27_10 <= io_A_Valid_0_delay_26_11;
    io_A_Valid_0_delay_28_9 <= io_A_Valid_0_delay_27_10;
    io_A_Valid_0_delay_29_8 <= io_A_Valid_0_delay_28_9;
    io_A_Valid_0_delay_30_7 <= io_A_Valid_0_delay_29_8;
    io_A_Valid_0_delay_31_6 <= io_A_Valid_0_delay_30_7;
    io_A_Valid_0_delay_32_5 <= io_A_Valid_0_delay_31_6;
    io_A_Valid_0_delay_33_4 <= io_A_Valid_0_delay_32_5;
    io_A_Valid_0_delay_34_3 <= io_A_Valid_0_delay_33_4;
    io_A_Valid_0_delay_35_2 <= io_A_Valid_0_delay_34_3;
    io_A_Valid_0_delay_36_1 <= io_A_Valid_0_delay_35_2;
    io_A_Valid_0_delay_37 <= io_A_Valid_0_delay_36_1;
    io_A_Valid_0_delay_1_37 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_36 <= io_A_Valid_0_delay_1_37;
    io_A_Valid_0_delay_3_35 <= io_A_Valid_0_delay_2_36;
    io_A_Valid_0_delay_4_34 <= io_A_Valid_0_delay_3_35;
    io_A_Valid_0_delay_5_33 <= io_A_Valid_0_delay_4_34;
    io_A_Valid_0_delay_6_32 <= io_A_Valid_0_delay_5_33;
    io_A_Valid_0_delay_7_31 <= io_A_Valid_0_delay_6_32;
    io_A_Valid_0_delay_8_30 <= io_A_Valid_0_delay_7_31;
    io_A_Valid_0_delay_9_29 <= io_A_Valid_0_delay_8_30;
    io_A_Valid_0_delay_10_28 <= io_A_Valid_0_delay_9_29;
    io_A_Valid_0_delay_11_27 <= io_A_Valid_0_delay_10_28;
    io_A_Valid_0_delay_12_26 <= io_A_Valid_0_delay_11_27;
    io_A_Valid_0_delay_13_25 <= io_A_Valid_0_delay_12_26;
    io_A_Valid_0_delay_14_24 <= io_A_Valid_0_delay_13_25;
    io_A_Valid_0_delay_15_23 <= io_A_Valid_0_delay_14_24;
    io_A_Valid_0_delay_16_22 <= io_A_Valid_0_delay_15_23;
    io_A_Valid_0_delay_17_21 <= io_A_Valid_0_delay_16_22;
    io_A_Valid_0_delay_18_20 <= io_A_Valid_0_delay_17_21;
    io_A_Valid_0_delay_19_19 <= io_A_Valid_0_delay_18_20;
    io_A_Valid_0_delay_20_18 <= io_A_Valid_0_delay_19_19;
    io_A_Valid_0_delay_21_17 <= io_A_Valid_0_delay_20_18;
    io_A_Valid_0_delay_22_16 <= io_A_Valid_0_delay_21_17;
    io_A_Valid_0_delay_23_15 <= io_A_Valid_0_delay_22_16;
    io_A_Valid_0_delay_24_14 <= io_A_Valid_0_delay_23_15;
    io_A_Valid_0_delay_25_13 <= io_A_Valid_0_delay_24_14;
    io_A_Valid_0_delay_26_12 <= io_A_Valid_0_delay_25_13;
    io_A_Valid_0_delay_27_11 <= io_A_Valid_0_delay_26_12;
    io_A_Valid_0_delay_28_10 <= io_A_Valid_0_delay_27_11;
    io_A_Valid_0_delay_29_9 <= io_A_Valid_0_delay_28_10;
    io_A_Valid_0_delay_30_8 <= io_A_Valid_0_delay_29_9;
    io_A_Valid_0_delay_31_7 <= io_A_Valid_0_delay_30_8;
    io_A_Valid_0_delay_32_6 <= io_A_Valid_0_delay_31_7;
    io_A_Valid_0_delay_33_5 <= io_A_Valid_0_delay_32_6;
    io_A_Valid_0_delay_34_4 <= io_A_Valid_0_delay_33_5;
    io_A_Valid_0_delay_35_3 <= io_A_Valid_0_delay_34_4;
    io_A_Valid_0_delay_36_2 <= io_A_Valid_0_delay_35_3;
    io_A_Valid_0_delay_37_1 <= io_A_Valid_0_delay_36_2;
    io_A_Valid_0_delay_38 <= io_A_Valid_0_delay_37_1;
    io_A_Valid_0_delay_1_38 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_37 <= io_A_Valid_0_delay_1_38;
    io_A_Valid_0_delay_3_36 <= io_A_Valid_0_delay_2_37;
    io_A_Valid_0_delay_4_35 <= io_A_Valid_0_delay_3_36;
    io_A_Valid_0_delay_5_34 <= io_A_Valid_0_delay_4_35;
    io_A_Valid_0_delay_6_33 <= io_A_Valid_0_delay_5_34;
    io_A_Valid_0_delay_7_32 <= io_A_Valid_0_delay_6_33;
    io_A_Valid_0_delay_8_31 <= io_A_Valid_0_delay_7_32;
    io_A_Valid_0_delay_9_30 <= io_A_Valid_0_delay_8_31;
    io_A_Valid_0_delay_10_29 <= io_A_Valid_0_delay_9_30;
    io_A_Valid_0_delay_11_28 <= io_A_Valid_0_delay_10_29;
    io_A_Valid_0_delay_12_27 <= io_A_Valid_0_delay_11_28;
    io_A_Valid_0_delay_13_26 <= io_A_Valid_0_delay_12_27;
    io_A_Valid_0_delay_14_25 <= io_A_Valid_0_delay_13_26;
    io_A_Valid_0_delay_15_24 <= io_A_Valid_0_delay_14_25;
    io_A_Valid_0_delay_16_23 <= io_A_Valid_0_delay_15_24;
    io_A_Valid_0_delay_17_22 <= io_A_Valid_0_delay_16_23;
    io_A_Valid_0_delay_18_21 <= io_A_Valid_0_delay_17_22;
    io_A_Valid_0_delay_19_20 <= io_A_Valid_0_delay_18_21;
    io_A_Valid_0_delay_20_19 <= io_A_Valid_0_delay_19_20;
    io_A_Valid_0_delay_21_18 <= io_A_Valid_0_delay_20_19;
    io_A_Valid_0_delay_22_17 <= io_A_Valid_0_delay_21_18;
    io_A_Valid_0_delay_23_16 <= io_A_Valid_0_delay_22_17;
    io_A_Valid_0_delay_24_15 <= io_A_Valid_0_delay_23_16;
    io_A_Valid_0_delay_25_14 <= io_A_Valid_0_delay_24_15;
    io_A_Valid_0_delay_26_13 <= io_A_Valid_0_delay_25_14;
    io_A_Valid_0_delay_27_12 <= io_A_Valid_0_delay_26_13;
    io_A_Valid_0_delay_28_11 <= io_A_Valid_0_delay_27_12;
    io_A_Valid_0_delay_29_10 <= io_A_Valid_0_delay_28_11;
    io_A_Valid_0_delay_30_9 <= io_A_Valid_0_delay_29_10;
    io_A_Valid_0_delay_31_8 <= io_A_Valid_0_delay_30_9;
    io_A_Valid_0_delay_32_7 <= io_A_Valid_0_delay_31_8;
    io_A_Valid_0_delay_33_6 <= io_A_Valid_0_delay_32_7;
    io_A_Valid_0_delay_34_5 <= io_A_Valid_0_delay_33_6;
    io_A_Valid_0_delay_35_4 <= io_A_Valid_0_delay_34_5;
    io_A_Valid_0_delay_36_3 <= io_A_Valid_0_delay_35_4;
    io_A_Valid_0_delay_37_2 <= io_A_Valid_0_delay_36_3;
    io_A_Valid_0_delay_38_1 <= io_A_Valid_0_delay_37_2;
    io_A_Valid_0_delay_39 <= io_A_Valid_0_delay_38_1;
    io_A_Valid_0_delay_1_39 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_38 <= io_A_Valid_0_delay_1_39;
    io_A_Valid_0_delay_3_37 <= io_A_Valid_0_delay_2_38;
    io_A_Valid_0_delay_4_36 <= io_A_Valid_0_delay_3_37;
    io_A_Valid_0_delay_5_35 <= io_A_Valid_0_delay_4_36;
    io_A_Valid_0_delay_6_34 <= io_A_Valid_0_delay_5_35;
    io_A_Valid_0_delay_7_33 <= io_A_Valid_0_delay_6_34;
    io_A_Valid_0_delay_8_32 <= io_A_Valid_0_delay_7_33;
    io_A_Valid_0_delay_9_31 <= io_A_Valid_0_delay_8_32;
    io_A_Valid_0_delay_10_30 <= io_A_Valid_0_delay_9_31;
    io_A_Valid_0_delay_11_29 <= io_A_Valid_0_delay_10_30;
    io_A_Valid_0_delay_12_28 <= io_A_Valid_0_delay_11_29;
    io_A_Valid_0_delay_13_27 <= io_A_Valid_0_delay_12_28;
    io_A_Valid_0_delay_14_26 <= io_A_Valid_0_delay_13_27;
    io_A_Valid_0_delay_15_25 <= io_A_Valid_0_delay_14_26;
    io_A_Valid_0_delay_16_24 <= io_A_Valid_0_delay_15_25;
    io_A_Valid_0_delay_17_23 <= io_A_Valid_0_delay_16_24;
    io_A_Valid_0_delay_18_22 <= io_A_Valid_0_delay_17_23;
    io_A_Valid_0_delay_19_21 <= io_A_Valid_0_delay_18_22;
    io_A_Valid_0_delay_20_20 <= io_A_Valid_0_delay_19_21;
    io_A_Valid_0_delay_21_19 <= io_A_Valid_0_delay_20_20;
    io_A_Valid_0_delay_22_18 <= io_A_Valid_0_delay_21_19;
    io_A_Valid_0_delay_23_17 <= io_A_Valid_0_delay_22_18;
    io_A_Valid_0_delay_24_16 <= io_A_Valid_0_delay_23_17;
    io_A_Valid_0_delay_25_15 <= io_A_Valid_0_delay_24_16;
    io_A_Valid_0_delay_26_14 <= io_A_Valid_0_delay_25_15;
    io_A_Valid_0_delay_27_13 <= io_A_Valid_0_delay_26_14;
    io_A_Valid_0_delay_28_12 <= io_A_Valid_0_delay_27_13;
    io_A_Valid_0_delay_29_11 <= io_A_Valid_0_delay_28_12;
    io_A_Valid_0_delay_30_10 <= io_A_Valid_0_delay_29_11;
    io_A_Valid_0_delay_31_9 <= io_A_Valid_0_delay_30_10;
    io_A_Valid_0_delay_32_8 <= io_A_Valid_0_delay_31_9;
    io_A_Valid_0_delay_33_7 <= io_A_Valid_0_delay_32_8;
    io_A_Valid_0_delay_34_6 <= io_A_Valid_0_delay_33_7;
    io_A_Valid_0_delay_35_5 <= io_A_Valid_0_delay_34_6;
    io_A_Valid_0_delay_36_4 <= io_A_Valid_0_delay_35_5;
    io_A_Valid_0_delay_37_3 <= io_A_Valid_0_delay_36_4;
    io_A_Valid_0_delay_38_2 <= io_A_Valid_0_delay_37_3;
    io_A_Valid_0_delay_39_1 <= io_A_Valid_0_delay_38_2;
    io_A_Valid_0_delay_40 <= io_A_Valid_0_delay_39_1;
    io_A_Valid_0_delay_1_40 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_39 <= io_A_Valid_0_delay_1_40;
    io_A_Valid_0_delay_3_38 <= io_A_Valid_0_delay_2_39;
    io_A_Valid_0_delay_4_37 <= io_A_Valid_0_delay_3_38;
    io_A_Valid_0_delay_5_36 <= io_A_Valid_0_delay_4_37;
    io_A_Valid_0_delay_6_35 <= io_A_Valid_0_delay_5_36;
    io_A_Valid_0_delay_7_34 <= io_A_Valid_0_delay_6_35;
    io_A_Valid_0_delay_8_33 <= io_A_Valid_0_delay_7_34;
    io_A_Valid_0_delay_9_32 <= io_A_Valid_0_delay_8_33;
    io_A_Valid_0_delay_10_31 <= io_A_Valid_0_delay_9_32;
    io_A_Valid_0_delay_11_30 <= io_A_Valid_0_delay_10_31;
    io_A_Valid_0_delay_12_29 <= io_A_Valid_0_delay_11_30;
    io_A_Valid_0_delay_13_28 <= io_A_Valid_0_delay_12_29;
    io_A_Valid_0_delay_14_27 <= io_A_Valid_0_delay_13_28;
    io_A_Valid_0_delay_15_26 <= io_A_Valid_0_delay_14_27;
    io_A_Valid_0_delay_16_25 <= io_A_Valid_0_delay_15_26;
    io_A_Valid_0_delay_17_24 <= io_A_Valid_0_delay_16_25;
    io_A_Valid_0_delay_18_23 <= io_A_Valid_0_delay_17_24;
    io_A_Valid_0_delay_19_22 <= io_A_Valid_0_delay_18_23;
    io_A_Valid_0_delay_20_21 <= io_A_Valid_0_delay_19_22;
    io_A_Valid_0_delay_21_20 <= io_A_Valid_0_delay_20_21;
    io_A_Valid_0_delay_22_19 <= io_A_Valid_0_delay_21_20;
    io_A_Valid_0_delay_23_18 <= io_A_Valid_0_delay_22_19;
    io_A_Valid_0_delay_24_17 <= io_A_Valid_0_delay_23_18;
    io_A_Valid_0_delay_25_16 <= io_A_Valid_0_delay_24_17;
    io_A_Valid_0_delay_26_15 <= io_A_Valid_0_delay_25_16;
    io_A_Valid_0_delay_27_14 <= io_A_Valid_0_delay_26_15;
    io_A_Valid_0_delay_28_13 <= io_A_Valid_0_delay_27_14;
    io_A_Valid_0_delay_29_12 <= io_A_Valid_0_delay_28_13;
    io_A_Valid_0_delay_30_11 <= io_A_Valid_0_delay_29_12;
    io_A_Valid_0_delay_31_10 <= io_A_Valid_0_delay_30_11;
    io_A_Valid_0_delay_32_9 <= io_A_Valid_0_delay_31_10;
    io_A_Valid_0_delay_33_8 <= io_A_Valid_0_delay_32_9;
    io_A_Valid_0_delay_34_7 <= io_A_Valid_0_delay_33_8;
    io_A_Valid_0_delay_35_6 <= io_A_Valid_0_delay_34_7;
    io_A_Valid_0_delay_36_5 <= io_A_Valid_0_delay_35_6;
    io_A_Valid_0_delay_37_4 <= io_A_Valid_0_delay_36_5;
    io_A_Valid_0_delay_38_3 <= io_A_Valid_0_delay_37_4;
    io_A_Valid_0_delay_39_2 <= io_A_Valid_0_delay_38_3;
    io_A_Valid_0_delay_40_1 <= io_A_Valid_0_delay_39_2;
    io_A_Valid_0_delay_41 <= io_A_Valid_0_delay_40_1;
    io_A_Valid_0_delay_1_41 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_40 <= io_A_Valid_0_delay_1_41;
    io_A_Valid_0_delay_3_39 <= io_A_Valid_0_delay_2_40;
    io_A_Valid_0_delay_4_38 <= io_A_Valid_0_delay_3_39;
    io_A_Valid_0_delay_5_37 <= io_A_Valid_0_delay_4_38;
    io_A_Valid_0_delay_6_36 <= io_A_Valid_0_delay_5_37;
    io_A_Valid_0_delay_7_35 <= io_A_Valid_0_delay_6_36;
    io_A_Valid_0_delay_8_34 <= io_A_Valid_0_delay_7_35;
    io_A_Valid_0_delay_9_33 <= io_A_Valid_0_delay_8_34;
    io_A_Valid_0_delay_10_32 <= io_A_Valid_0_delay_9_33;
    io_A_Valid_0_delay_11_31 <= io_A_Valid_0_delay_10_32;
    io_A_Valid_0_delay_12_30 <= io_A_Valid_0_delay_11_31;
    io_A_Valid_0_delay_13_29 <= io_A_Valid_0_delay_12_30;
    io_A_Valid_0_delay_14_28 <= io_A_Valid_0_delay_13_29;
    io_A_Valid_0_delay_15_27 <= io_A_Valid_0_delay_14_28;
    io_A_Valid_0_delay_16_26 <= io_A_Valid_0_delay_15_27;
    io_A_Valid_0_delay_17_25 <= io_A_Valid_0_delay_16_26;
    io_A_Valid_0_delay_18_24 <= io_A_Valid_0_delay_17_25;
    io_A_Valid_0_delay_19_23 <= io_A_Valid_0_delay_18_24;
    io_A_Valid_0_delay_20_22 <= io_A_Valid_0_delay_19_23;
    io_A_Valid_0_delay_21_21 <= io_A_Valid_0_delay_20_22;
    io_A_Valid_0_delay_22_20 <= io_A_Valid_0_delay_21_21;
    io_A_Valid_0_delay_23_19 <= io_A_Valid_0_delay_22_20;
    io_A_Valid_0_delay_24_18 <= io_A_Valid_0_delay_23_19;
    io_A_Valid_0_delay_25_17 <= io_A_Valid_0_delay_24_18;
    io_A_Valid_0_delay_26_16 <= io_A_Valid_0_delay_25_17;
    io_A_Valid_0_delay_27_15 <= io_A_Valid_0_delay_26_16;
    io_A_Valid_0_delay_28_14 <= io_A_Valid_0_delay_27_15;
    io_A_Valid_0_delay_29_13 <= io_A_Valid_0_delay_28_14;
    io_A_Valid_0_delay_30_12 <= io_A_Valid_0_delay_29_13;
    io_A_Valid_0_delay_31_11 <= io_A_Valid_0_delay_30_12;
    io_A_Valid_0_delay_32_10 <= io_A_Valid_0_delay_31_11;
    io_A_Valid_0_delay_33_9 <= io_A_Valid_0_delay_32_10;
    io_A_Valid_0_delay_34_8 <= io_A_Valid_0_delay_33_9;
    io_A_Valid_0_delay_35_7 <= io_A_Valid_0_delay_34_8;
    io_A_Valid_0_delay_36_6 <= io_A_Valid_0_delay_35_7;
    io_A_Valid_0_delay_37_5 <= io_A_Valid_0_delay_36_6;
    io_A_Valid_0_delay_38_4 <= io_A_Valid_0_delay_37_5;
    io_A_Valid_0_delay_39_3 <= io_A_Valid_0_delay_38_4;
    io_A_Valid_0_delay_40_2 <= io_A_Valid_0_delay_39_3;
    io_A_Valid_0_delay_41_1 <= io_A_Valid_0_delay_40_2;
    io_A_Valid_0_delay_42 <= io_A_Valid_0_delay_41_1;
    io_A_Valid_0_delay_1_42 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_41 <= io_A_Valid_0_delay_1_42;
    io_A_Valid_0_delay_3_40 <= io_A_Valid_0_delay_2_41;
    io_A_Valid_0_delay_4_39 <= io_A_Valid_0_delay_3_40;
    io_A_Valid_0_delay_5_38 <= io_A_Valid_0_delay_4_39;
    io_A_Valid_0_delay_6_37 <= io_A_Valid_0_delay_5_38;
    io_A_Valid_0_delay_7_36 <= io_A_Valid_0_delay_6_37;
    io_A_Valid_0_delay_8_35 <= io_A_Valid_0_delay_7_36;
    io_A_Valid_0_delay_9_34 <= io_A_Valid_0_delay_8_35;
    io_A_Valid_0_delay_10_33 <= io_A_Valid_0_delay_9_34;
    io_A_Valid_0_delay_11_32 <= io_A_Valid_0_delay_10_33;
    io_A_Valid_0_delay_12_31 <= io_A_Valid_0_delay_11_32;
    io_A_Valid_0_delay_13_30 <= io_A_Valid_0_delay_12_31;
    io_A_Valid_0_delay_14_29 <= io_A_Valid_0_delay_13_30;
    io_A_Valid_0_delay_15_28 <= io_A_Valid_0_delay_14_29;
    io_A_Valid_0_delay_16_27 <= io_A_Valid_0_delay_15_28;
    io_A_Valid_0_delay_17_26 <= io_A_Valid_0_delay_16_27;
    io_A_Valid_0_delay_18_25 <= io_A_Valid_0_delay_17_26;
    io_A_Valid_0_delay_19_24 <= io_A_Valid_0_delay_18_25;
    io_A_Valid_0_delay_20_23 <= io_A_Valid_0_delay_19_24;
    io_A_Valid_0_delay_21_22 <= io_A_Valid_0_delay_20_23;
    io_A_Valid_0_delay_22_21 <= io_A_Valid_0_delay_21_22;
    io_A_Valid_0_delay_23_20 <= io_A_Valid_0_delay_22_21;
    io_A_Valid_0_delay_24_19 <= io_A_Valid_0_delay_23_20;
    io_A_Valid_0_delay_25_18 <= io_A_Valid_0_delay_24_19;
    io_A_Valid_0_delay_26_17 <= io_A_Valid_0_delay_25_18;
    io_A_Valid_0_delay_27_16 <= io_A_Valid_0_delay_26_17;
    io_A_Valid_0_delay_28_15 <= io_A_Valid_0_delay_27_16;
    io_A_Valid_0_delay_29_14 <= io_A_Valid_0_delay_28_15;
    io_A_Valid_0_delay_30_13 <= io_A_Valid_0_delay_29_14;
    io_A_Valid_0_delay_31_12 <= io_A_Valid_0_delay_30_13;
    io_A_Valid_0_delay_32_11 <= io_A_Valid_0_delay_31_12;
    io_A_Valid_0_delay_33_10 <= io_A_Valid_0_delay_32_11;
    io_A_Valid_0_delay_34_9 <= io_A_Valid_0_delay_33_10;
    io_A_Valid_0_delay_35_8 <= io_A_Valid_0_delay_34_9;
    io_A_Valid_0_delay_36_7 <= io_A_Valid_0_delay_35_8;
    io_A_Valid_0_delay_37_6 <= io_A_Valid_0_delay_36_7;
    io_A_Valid_0_delay_38_5 <= io_A_Valid_0_delay_37_6;
    io_A_Valid_0_delay_39_4 <= io_A_Valid_0_delay_38_5;
    io_A_Valid_0_delay_40_3 <= io_A_Valid_0_delay_39_4;
    io_A_Valid_0_delay_41_2 <= io_A_Valid_0_delay_40_3;
    io_A_Valid_0_delay_42_1 <= io_A_Valid_0_delay_41_2;
    io_A_Valid_0_delay_43 <= io_A_Valid_0_delay_42_1;
    io_A_Valid_0_delay_1_43 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_42 <= io_A_Valid_0_delay_1_43;
    io_A_Valid_0_delay_3_41 <= io_A_Valid_0_delay_2_42;
    io_A_Valid_0_delay_4_40 <= io_A_Valid_0_delay_3_41;
    io_A_Valid_0_delay_5_39 <= io_A_Valid_0_delay_4_40;
    io_A_Valid_0_delay_6_38 <= io_A_Valid_0_delay_5_39;
    io_A_Valid_0_delay_7_37 <= io_A_Valid_0_delay_6_38;
    io_A_Valid_0_delay_8_36 <= io_A_Valid_0_delay_7_37;
    io_A_Valid_0_delay_9_35 <= io_A_Valid_0_delay_8_36;
    io_A_Valid_0_delay_10_34 <= io_A_Valid_0_delay_9_35;
    io_A_Valid_0_delay_11_33 <= io_A_Valid_0_delay_10_34;
    io_A_Valid_0_delay_12_32 <= io_A_Valid_0_delay_11_33;
    io_A_Valid_0_delay_13_31 <= io_A_Valid_0_delay_12_32;
    io_A_Valid_0_delay_14_30 <= io_A_Valid_0_delay_13_31;
    io_A_Valid_0_delay_15_29 <= io_A_Valid_0_delay_14_30;
    io_A_Valid_0_delay_16_28 <= io_A_Valid_0_delay_15_29;
    io_A_Valid_0_delay_17_27 <= io_A_Valid_0_delay_16_28;
    io_A_Valid_0_delay_18_26 <= io_A_Valid_0_delay_17_27;
    io_A_Valid_0_delay_19_25 <= io_A_Valid_0_delay_18_26;
    io_A_Valid_0_delay_20_24 <= io_A_Valid_0_delay_19_25;
    io_A_Valid_0_delay_21_23 <= io_A_Valid_0_delay_20_24;
    io_A_Valid_0_delay_22_22 <= io_A_Valid_0_delay_21_23;
    io_A_Valid_0_delay_23_21 <= io_A_Valid_0_delay_22_22;
    io_A_Valid_0_delay_24_20 <= io_A_Valid_0_delay_23_21;
    io_A_Valid_0_delay_25_19 <= io_A_Valid_0_delay_24_20;
    io_A_Valid_0_delay_26_18 <= io_A_Valid_0_delay_25_19;
    io_A_Valid_0_delay_27_17 <= io_A_Valid_0_delay_26_18;
    io_A_Valid_0_delay_28_16 <= io_A_Valid_0_delay_27_17;
    io_A_Valid_0_delay_29_15 <= io_A_Valid_0_delay_28_16;
    io_A_Valid_0_delay_30_14 <= io_A_Valid_0_delay_29_15;
    io_A_Valid_0_delay_31_13 <= io_A_Valid_0_delay_30_14;
    io_A_Valid_0_delay_32_12 <= io_A_Valid_0_delay_31_13;
    io_A_Valid_0_delay_33_11 <= io_A_Valid_0_delay_32_12;
    io_A_Valid_0_delay_34_10 <= io_A_Valid_0_delay_33_11;
    io_A_Valid_0_delay_35_9 <= io_A_Valid_0_delay_34_10;
    io_A_Valid_0_delay_36_8 <= io_A_Valid_0_delay_35_9;
    io_A_Valid_0_delay_37_7 <= io_A_Valid_0_delay_36_8;
    io_A_Valid_0_delay_38_6 <= io_A_Valid_0_delay_37_7;
    io_A_Valid_0_delay_39_5 <= io_A_Valid_0_delay_38_6;
    io_A_Valid_0_delay_40_4 <= io_A_Valid_0_delay_39_5;
    io_A_Valid_0_delay_41_3 <= io_A_Valid_0_delay_40_4;
    io_A_Valid_0_delay_42_2 <= io_A_Valid_0_delay_41_3;
    io_A_Valid_0_delay_43_1 <= io_A_Valid_0_delay_42_2;
    io_A_Valid_0_delay_44 <= io_A_Valid_0_delay_43_1;
    io_A_Valid_0_delay_1_44 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_43 <= io_A_Valid_0_delay_1_44;
    io_A_Valid_0_delay_3_42 <= io_A_Valid_0_delay_2_43;
    io_A_Valid_0_delay_4_41 <= io_A_Valid_0_delay_3_42;
    io_A_Valid_0_delay_5_40 <= io_A_Valid_0_delay_4_41;
    io_A_Valid_0_delay_6_39 <= io_A_Valid_0_delay_5_40;
    io_A_Valid_0_delay_7_38 <= io_A_Valid_0_delay_6_39;
    io_A_Valid_0_delay_8_37 <= io_A_Valid_0_delay_7_38;
    io_A_Valid_0_delay_9_36 <= io_A_Valid_0_delay_8_37;
    io_A_Valid_0_delay_10_35 <= io_A_Valid_0_delay_9_36;
    io_A_Valid_0_delay_11_34 <= io_A_Valid_0_delay_10_35;
    io_A_Valid_0_delay_12_33 <= io_A_Valid_0_delay_11_34;
    io_A_Valid_0_delay_13_32 <= io_A_Valid_0_delay_12_33;
    io_A_Valid_0_delay_14_31 <= io_A_Valid_0_delay_13_32;
    io_A_Valid_0_delay_15_30 <= io_A_Valid_0_delay_14_31;
    io_A_Valid_0_delay_16_29 <= io_A_Valid_0_delay_15_30;
    io_A_Valid_0_delay_17_28 <= io_A_Valid_0_delay_16_29;
    io_A_Valid_0_delay_18_27 <= io_A_Valid_0_delay_17_28;
    io_A_Valid_0_delay_19_26 <= io_A_Valid_0_delay_18_27;
    io_A_Valid_0_delay_20_25 <= io_A_Valid_0_delay_19_26;
    io_A_Valid_0_delay_21_24 <= io_A_Valid_0_delay_20_25;
    io_A_Valid_0_delay_22_23 <= io_A_Valid_0_delay_21_24;
    io_A_Valid_0_delay_23_22 <= io_A_Valid_0_delay_22_23;
    io_A_Valid_0_delay_24_21 <= io_A_Valid_0_delay_23_22;
    io_A_Valid_0_delay_25_20 <= io_A_Valid_0_delay_24_21;
    io_A_Valid_0_delay_26_19 <= io_A_Valid_0_delay_25_20;
    io_A_Valid_0_delay_27_18 <= io_A_Valid_0_delay_26_19;
    io_A_Valid_0_delay_28_17 <= io_A_Valid_0_delay_27_18;
    io_A_Valid_0_delay_29_16 <= io_A_Valid_0_delay_28_17;
    io_A_Valid_0_delay_30_15 <= io_A_Valid_0_delay_29_16;
    io_A_Valid_0_delay_31_14 <= io_A_Valid_0_delay_30_15;
    io_A_Valid_0_delay_32_13 <= io_A_Valid_0_delay_31_14;
    io_A_Valid_0_delay_33_12 <= io_A_Valid_0_delay_32_13;
    io_A_Valid_0_delay_34_11 <= io_A_Valid_0_delay_33_12;
    io_A_Valid_0_delay_35_10 <= io_A_Valid_0_delay_34_11;
    io_A_Valid_0_delay_36_9 <= io_A_Valid_0_delay_35_10;
    io_A_Valid_0_delay_37_8 <= io_A_Valid_0_delay_36_9;
    io_A_Valid_0_delay_38_7 <= io_A_Valid_0_delay_37_8;
    io_A_Valid_0_delay_39_6 <= io_A_Valid_0_delay_38_7;
    io_A_Valid_0_delay_40_5 <= io_A_Valid_0_delay_39_6;
    io_A_Valid_0_delay_41_4 <= io_A_Valid_0_delay_40_5;
    io_A_Valid_0_delay_42_3 <= io_A_Valid_0_delay_41_4;
    io_A_Valid_0_delay_43_2 <= io_A_Valid_0_delay_42_3;
    io_A_Valid_0_delay_44_1 <= io_A_Valid_0_delay_43_2;
    io_A_Valid_0_delay_45 <= io_A_Valid_0_delay_44_1;
    io_A_Valid_0_delay_1_45 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_44 <= io_A_Valid_0_delay_1_45;
    io_A_Valid_0_delay_3_43 <= io_A_Valid_0_delay_2_44;
    io_A_Valid_0_delay_4_42 <= io_A_Valid_0_delay_3_43;
    io_A_Valid_0_delay_5_41 <= io_A_Valid_0_delay_4_42;
    io_A_Valid_0_delay_6_40 <= io_A_Valid_0_delay_5_41;
    io_A_Valid_0_delay_7_39 <= io_A_Valid_0_delay_6_40;
    io_A_Valid_0_delay_8_38 <= io_A_Valid_0_delay_7_39;
    io_A_Valid_0_delay_9_37 <= io_A_Valid_0_delay_8_38;
    io_A_Valid_0_delay_10_36 <= io_A_Valid_0_delay_9_37;
    io_A_Valid_0_delay_11_35 <= io_A_Valid_0_delay_10_36;
    io_A_Valid_0_delay_12_34 <= io_A_Valid_0_delay_11_35;
    io_A_Valid_0_delay_13_33 <= io_A_Valid_0_delay_12_34;
    io_A_Valid_0_delay_14_32 <= io_A_Valid_0_delay_13_33;
    io_A_Valid_0_delay_15_31 <= io_A_Valid_0_delay_14_32;
    io_A_Valid_0_delay_16_30 <= io_A_Valid_0_delay_15_31;
    io_A_Valid_0_delay_17_29 <= io_A_Valid_0_delay_16_30;
    io_A_Valid_0_delay_18_28 <= io_A_Valid_0_delay_17_29;
    io_A_Valid_0_delay_19_27 <= io_A_Valid_0_delay_18_28;
    io_A_Valid_0_delay_20_26 <= io_A_Valid_0_delay_19_27;
    io_A_Valid_0_delay_21_25 <= io_A_Valid_0_delay_20_26;
    io_A_Valid_0_delay_22_24 <= io_A_Valid_0_delay_21_25;
    io_A_Valid_0_delay_23_23 <= io_A_Valid_0_delay_22_24;
    io_A_Valid_0_delay_24_22 <= io_A_Valid_0_delay_23_23;
    io_A_Valid_0_delay_25_21 <= io_A_Valid_0_delay_24_22;
    io_A_Valid_0_delay_26_20 <= io_A_Valid_0_delay_25_21;
    io_A_Valid_0_delay_27_19 <= io_A_Valid_0_delay_26_20;
    io_A_Valid_0_delay_28_18 <= io_A_Valid_0_delay_27_19;
    io_A_Valid_0_delay_29_17 <= io_A_Valid_0_delay_28_18;
    io_A_Valid_0_delay_30_16 <= io_A_Valid_0_delay_29_17;
    io_A_Valid_0_delay_31_15 <= io_A_Valid_0_delay_30_16;
    io_A_Valid_0_delay_32_14 <= io_A_Valid_0_delay_31_15;
    io_A_Valid_0_delay_33_13 <= io_A_Valid_0_delay_32_14;
    io_A_Valid_0_delay_34_12 <= io_A_Valid_0_delay_33_13;
    io_A_Valid_0_delay_35_11 <= io_A_Valid_0_delay_34_12;
    io_A_Valid_0_delay_36_10 <= io_A_Valid_0_delay_35_11;
    io_A_Valid_0_delay_37_9 <= io_A_Valid_0_delay_36_10;
    io_A_Valid_0_delay_38_8 <= io_A_Valid_0_delay_37_9;
    io_A_Valid_0_delay_39_7 <= io_A_Valid_0_delay_38_8;
    io_A_Valid_0_delay_40_6 <= io_A_Valid_0_delay_39_7;
    io_A_Valid_0_delay_41_5 <= io_A_Valid_0_delay_40_6;
    io_A_Valid_0_delay_42_4 <= io_A_Valid_0_delay_41_5;
    io_A_Valid_0_delay_43_3 <= io_A_Valid_0_delay_42_4;
    io_A_Valid_0_delay_44_2 <= io_A_Valid_0_delay_43_3;
    io_A_Valid_0_delay_45_1 <= io_A_Valid_0_delay_44_2;
    io_A_Valid_0_delay_46 <= io_A_Valid_0_delay_45_1;
    io_A_Valid_0_delay_1_46 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_45 <= io_A_Valid_0_delay_1_46;
    io_A_Valid_0_delay_3_44 <= io_A_Valid_0_delay_2_45;
    io_A_Valid_0_delay_4_43 <= io_A_Valid_0_delay_3_44;
    io_A_Valid_0_delay_5_42 <= io_A_Valid_0_delay_4_43;
    io_A_Valid_0_delay_6_41 <= io_A_Valid_0_delay_5_42;
    io_A_Valid_0_delay_7_40 <= io_A_Valid_0_delay_6_41;
    io_A_Valid_0_delay_8_39 <= io_A_Valid_0_delay_7_40;
    io_A_Valid_0_delay_9_38 <= io_A_Valid_0_delay_8_39;
    io_A_Valid_0_delay_10_37 <= io_A_Valid_0_delay_9_38;
    io_A_Valid_0_delay_11_36 <= io_A_Valid_0_delay_10_37;
    io_A_Valid_0_delay_12_35 <= io_A_Valid_0_delay_11_36;
    io_A_Valid_0_delay_13_34 <= io_A_Valid_0_delay_12_35;
    io_A_Valid_0_delay_14_33 <= io_A_Valid_0_delay_13_34;
    io_A_Valid_0_delay_15_32 <= io_A_Valid_0_delay_14_33;
    io_A_Valid_0_delay_16_31 <= io_A_Valid_0_delay_15_32;
    io_A_Valid_0_delay_17_30 <= io_A_Valid_0_delay_16_31;
    io_A_Valid_0_delay_18_29 <= io_A_Valid_0_delay_17_30;
    io_A_Valid_0_delay_19_28 <= io_A_Valid_0_delay_18_29;
    io_A_Valid_0_delay_20_27 <= io_A_Valid_0_delay_19_28;
    io_A_Valid_0_delay_21_26 <= io_A_Valid_0_delay_20_27;
    io_A_Valid_0_delay_22_25 <= io_A_Valid_0_delay_21_26;
    io_A_Valid_0_delay_23_24 <= io_A_Valid_0_delay_22_25;
    io_A_Valid_0_delay_24_23 <= io_A_Valid_0_delay_23_24;
    io_A_Valid_0_delay_25_22 <= io_A_Valid_0_delay_24_23;
    io_A_Valid_0_delay_26_21 <= io_A_Valid_0_delay_25_22;
    io_A_Valid_0_delay_27_20 <= io_A_Valid_0_delay_26_21;
    io_A_Valid_0_delay_28_19 <= io_A_Valid_0_delay_27_20;
    io_A_Valid_0_delay_29_18 <= io_A_Valid_0_delay_28_19;
    io_A_Valid_0_delay_30_17 <= io_A_Valid_0_delay_29_18;
    io_A_Valid_0_delay_31_16 <= io_A_Valid_0_delay_30_17;
    io_A_Valid_0_delay_32_15 <= io_A_Valid_0_delay_31_16;
    io_A_Valid_0_delay_33_14 <= io_A_Valid_0_delay_32_15;
    io_A_Valid_0_delay_34_13 <= io_A_Valid_0_delay_33_14;
    io_A_Valid_0_delay_35_12 <= io_A_Valid_0_delay_34_13;
    io_A_Valid_0_delay_36_11 <= io_A_Valid_0_delay_35_12;
    io_A_Valid_0_delay_37_10 <= io_A_Valid_0_delay_36_11;
    io_A_Valid_0_delay_38_9 <= io_A_Valid_0_delay_37_10;
    io_A_Valid_0_delay_39_8 <= io_A_Valid_0_delay_38_9;
    io_A_Valid_0_delay_40_7 <= io_A_Valid_0_delay_39_8;
    io_A_Valid_0_delay_41_6 <= io_A_Valid_0_delay_40_7;
    io_A_Valid_0_delay_42_5 <= io_A_Valid_0_delay_41_6;
    io_A_Valid_0_delay_43_4 <= io_A_Valid_0_delay_42_5;
    io_A_Valid_0_delay_44_3 <= io_A_Valid_0_delay_43_4;
    io_A_Valid_0_delay_45_2 <= io_A_Valid_0_delay_44_3;
    io_A_Valid_0_delay_46_1 <= io_A_Valid_0_delay_45_2;
    io_A_Valid_0_delay_47 <= io_A_Valid_0_delay_46_1;
    io_A_Valid_0_delay_1_47 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_46 <= io_A_Valid_0_delay_1_47;
    io_A_Valid_0_delay_3_45 <= io_A_Valid_0_delay_2_46;
    io_A_Valid_0_delay_4_44 <= io_A_Valid_0_delay_3_45;
    io_A_Valid_0_delay_5_43 <= io_A_Valid_0_delay_4_44;
    io_A_Valid_0_delay_6_42 <= io_A_Valid_0_delay_5_43;
    io_A_Valid_0_delay_7_41 <= io_A_Valid_0_delay_6_42;
    io_A_Valid_0_delay_8_40 <= io_A_Valid_0_delay_7_41;
    io_A_Valid_0_delay_9_39 <= io_A_Valid_0_delay_8_40;
    io_A_Valid_0_delay_10_38 <= io_A_Valid_0_delay_9_39;
    io_A_Valid_0_delay_11_37 <= io_A_Valid_0_delay_10_38;
    io_A_Valid_0_delay_12_36 <= io_A_Valid_0_delay_11_37;
    io_A_Valid_0_delay_13_35 <= io_A_Valid_0_delay_12_36;
    io_A_Valid_0_delay_14_34 <= io_A_Valid_0_delay_13_35;
    io_A_Valid_0_delay_15_33 <= io_A_Valid_0_delay_14_34;
    io_A_Valid_0_delay_16_32 <= io_A_Valid_0_delay_15_33;
    io_A_Valid_0_delay_17_31 <= io_A_Valid_0_delay_16_32;
    io_A_Valid_0_delay_18_30 <= io_A_Valid_0_delay_17_31;
    io_A_Valid_0_delay_19_29 <= io_A_Valid_0_delay_18_30;
    io_A_Valid_0_delay_20_28 <= io_A_Valid_0_delay_19_29;
    io_A_Valid_0_delay_21_27 <= io_A_Valid_0_delay_20_28;
    io_A_Valid_0_delay_22_26 <= io_A_Valid_0_delay_21_27;
    io_A_Valid_0_delay_23_25 <= io_A_Valid_0_delay_22_26;
    io_A_Valid_0_delay_24_24 <= io_A_Valid_0_delay_23_25;
    io_A_Valid_0_delay_25_23 <= io_A_Valid_0_delay_24_24;
    io_A_Valid_0_delay_26_22 <= io_A_Valid_0_delay_25_23;
    io_A_Valid_0_delay_27_21 <= io_A_Valid_0_delay_26_22;
    io_A_Valid_0_delay_28_20 <= io_A_Valid_0_delay_27_21;
    io_A_Valid_0_delay_29_19 <= io_A_Valid_0_delay_28_20;
    io_A_Valid_0_delay_30_18 <= io_A_Valid_0_delay_29_19;
    io_A_Valid_0_delay_31_17 <= io_A_Valid_0_delay_30_18;
    io_A_Valid_0_delay_32_16 <= io_A_Valid_0_delay_31_17;
    io_A_Valid_0_delay_33_15 <= io_A_Valid_0_delay_32_16;
    io_A_Valid_0_delay_34_14 <= io_A_Valid_0_delay_33_15;
    io_A_Valid_0_delay_35_13 <= io_A_Valid_0_delay_34_14;
    io_A_Valid_0_delay_36_12 <= io_A_Valid_0_delay_35_13;
    io_A_Valid_0_delay_37_11 <= io_A_Valid_0_delay_36_12;
    io_A_Valid_0_delay_38_10 <= io_A_Valid_0_delay_37_11;
    io_A_Valid_0_delay_39_9 <= io_A_Valid_0_delay_38_10;
    io_A_Valid_0_delay_40_8 <= io_A_Valid_0_delay_39_9;
    io_A_Valid_0_delay_41_7 <= io_A_Valid_0_delay_40_8;
    io_A_Valid_0_delay_42_6 <= io_A_Valid_0_delay_41_7;
    io_A_Valid_0_delay_43_5 <= io_A_Valid_0_delay_42_6;
    io_A_Valid_0_delay_44_4 <= io_A_Valid_0_delay_43_5;
    io_A_Valid_0_delay_45_3 <= io_A_Valid_0_delay_44_4;
    io_A_Valid_0_delay_46_2 <= io_A_Valid_0_delay_45_3;
    io_A_Valid_0_delay_47_1 <= io_A_Valid_0_delay_46_2;
    io_A_Valid_0_delay_48 <= io_A_Valid_0_delay_47_1;
    io_A_Valid_0_delay_1_48 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_47 <= io_A_Valid_0_delay_1_48;
    io_A_Valid_0_delay_3_46 <= io_A_Valid_0_delay_2_47;
    io_A_Valid_0_delay_4_45 <= io_A_Valid_0_delay_3_46;
    io_A_Valid_0_delay_5_44 <= io_A_Valid_0_delay_4_45;
    io_A_Valid_0_delay_6_43 <= io_A_Valid_0_delay_5_44;
    io_A_Valid_0_delay_7_42 <= io_A_Valid_0_delay_6_43;
    io_A_Valid_0_delay_8_41 <= io_A_Valid_0_delay_7_42;
    io_A_Valid_0_delay_9_40 <= io_A_Valid_0_delay_8_41;
    io_A_Valid_0_delay_10_39 <= io_A_Valid_0_delay_9_40;
    io_A_Valid_0_delay_11_38 <= io_A_Valid_0_delay_10_39;
    io_A_Valid_0_delay_12_37 <= io_A_Valid_0_delay_11_38;
    io_A_Valid_0_delay_13_36 <= io_A_Valid_0_delay_12_37;
    io_A_Valid_0_delay_14_35 <= io_A_Valid_0_delay_13_36;
    io_A_Valid_0_delay_15_34 <= io_A_Valid_0_delay_14_35;
    io_A_Valid_0_delay_16_33 <= io_A_Valid_0_delay_15_34;
    io_A_Valid_0_delay_17_32 <= io_A_Valid_0_delay_16_33;
    io_A_Valid_0_delay_18_31 <= io_A_Valid_0_delay_17_32;
    io_A_Valid_0_delay_19_30 <= io_A_Valid_0_delay_18_31;
    io_A_Valid_0_delay_20_29 <= io_A_Valid_0_delay_19_30;
    io_A_Valid_0_delay_21_28 <= io_A_Valid_0_delay_20_29;
    io_A_Valid_0_delay_22_27 <= io_A_Valid_0_delay_21_28;
    io_A_Valid_0_delay_23_26 <= io_A_Valid_0_delay_22_27;
    io_A_Valid_0_delay_24_25 <= io_A_Valid_0_delay_23_26;
    io_A_Valid_0_delay_25_24 <= io_A_Valid_0_delay_24_25;
    io_A_Valid_0_delay_26_23 <= io_A_Valid_0_delay_25_24;
    io_A_Valid_0_delay_27_22 <= io_A_Valid_0_delay_26_23;
    io_A_Valid_0_delay_28_21 <= io_A_Valid_0_delay_27_22;
    io_A_Valid_0_delay_29_20 <= io_A_Valid_0_delay_28_21;
    io_A_Valid_0_delay_30_19 <= io_A_Valid_0_delay_29_20;
    io_A_Valid_0_delay_31_18 <= io_A_Valid_0_delay_30_19;
    io_A_Valid_0_delay_32_17 <= io_A_Valid_0_delay_31_18;
    io_A_Valid_0_delay_33_16 <= io_A_Valid_0_delay_32_17;
    io_A_Valid_0_delay_34_15 <= io_A_Valid_0_delay_33_16;
    io_A_Valid_0_delay_35_14 <= io_A_Valid_0_delay_34_15;
    io_A_Valid_0_delay_36_13 <= io_A_Valid_0_delay_35_14;
    io_A_Valid_0_delay_37_12 <= io_A_Valid_0_delay_36_13;
    io_A_Valid_0_delay_38_11 <= io_A_Valid_0_delay_37_12;
    io_A_Valid_0_delay_39_10 <= io_A_Valid_0_delay_38_11;
    io_A_Valid_0_delay_40_9 <= io_A_Valid_0_delay_39_10;
    io_A_Valid_0_delay_41_8 <= io_A_Valid_0_delay_40_9;
    io_A_Valid_0_delay_42_7 <= io_A_Valid_0_delay_41_8;
    io_A_Valid_0_delay_43_6 <= io_A_Valid_0_delay_42_7;
    io_A_Valid_0_delay_44_5 <= io_A_Valid_0_delay_43_6;
    io_A_Valid_0_delay_45_4 <= io_A_Valid_0_delay_44_5;
    io_A_Valid_0_delay_46_3 <= io_A_Valid_0_delay_45_4;
    io_A_Valid_0_delay_47_2 <= io_A_Valid_0_delay_46_3;
    io_A_Valid_0_delay_48_1 <= io_A_Valid_0_delay_47_2;
    io_A_Valid_0_delay_49 <= io_A_Valid_0_delay_48_1;
    io_A_Valid_0_delay_1_49 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_48 <= io_A_Valid_0_delay_1_49;
    io_A_Valid_0_delay_3_47 <= io_A_Valid_0_delay_2_48;
    io_A_Valid_0_delay_4_46 <= io_A_Valid_0_delay_3_47;
    io_A_Valid_0_delay_5_45 <= io_A_Valid_0_delay_4_46;
    io_A_Valid_0_delay_6_44 <= io_A_Valid_0_delay_5_45;
    io_A_Valid_0_delay_7_43 <= io_A_Valid_0_delay_6_44;
    io_A_Valid_0_delay_8_42 <= io_A_Valid_0_delay_7_43;
    io_A_Valid_0_delay_9_41 <= io_A_Valid_0_delay_8_42;
    io_A_Valid_0_delay_10_40 <= io_A_Valid_0_delay_9_41;
    io_A_Valid_0_delay_11_39 <= io_A_Valid_0_delay_10_40;
    io_A_Valid_0_delay_12_38 <= io_A_Valid_0_delay_11_39;
    io_A_Valid_0_delay_13_37 <= io_A_Valid_0_delay_12_38;
    io_A_Valid_0_delay_14_36 <= io_A_Valid_0_delay_13_37;
    io_A_Valid_0_delay_15_35 <= io_A_Valid_0_delay_14_36;
    io_A_Valid_0_delay_16_34 <= io_A_Valid_0_delay_15_35;
    io_A_Valid_0_delay_17_33 <= io_A_Valid_0_delay_16_34;
    io_A_Valid_0_delay_18_32 <= io_A_Valid_0_delay_17_33;
    io_A_Valid_0_delay_19_31 <= io_A_Valid_0_delay_18_32;
    io_A_Valid_0_delay_20_30 <= io_A_Valid_0_delay_19_31;
    io_A_Valid_0_delay_21_29 <= io_A_Valid_0_delay_20_30;
    io_A_Valid_0_delay_22_28 <= io_A_Valid_0_delay_21_29;
    io_A_Valid_0_delay_23_27 <= io_A_Valid_0_delay_22_28;
    io_A_Valid_0_delay_24_26 <= io_A_Valid_0_delay_23_27;
    io_A_Valid_0_delay_25_25 <= io_A_Valid_0_delay_24_26;
    io_A_Valid_0_delay_26_24 <= io_A_Valid_0_delay_25_25;
    io_A_Valid_0_delay_27_23 <= io_A_Valid_0_delay_26_24;
    io_A_Valid_0_delay_28_22 <= io_A_Valid_0_delay_27_23;
    io_A_Valid_0_delay_29_21 <= io_A_Valid_0_delay_28_22;
    io_A_Valid_0_delay_30_20 <= io_A_Valid_0_delay_29_21;
    io_A_Valid_0_delay_31_19 <= io_A_Valid_0_delay_30_20;
    io_A_Valid_0_delay_32_18 <= io_A_Valid_0_delay_31_19;
    io_A_Valid_0_delay_33_17 <= io_A_Valid_0_delay_32_18;
    io_A_Valid_0_delay_34_16 <= io_A_Valid_0_delay_33_17;
    io_A_Valid_0_delay_35_15 <= io_A_Valid_0_delay_34_16;
    io_A_Valid_0_delay_36_14 <= io_A_Valid_0_delay_35_15;
    io_A_Valid_0_delay_37_13 <= io_A_Valid_0_delay_36_14;
    io_A_Valid_0_delay_38_12 <= io_A_Valid_0_delay_37_13;
    io_A_Valid_0_delay_39_11 <= io_A_Valid_0_delay_38_12;
    io_A_Valid_0_delay_40_10 <= io_A_Valid_0_delay_39_11;
    io_A_Valid_0_delay_41_9 <= io_A_Valid_0_delay_40_10;
    io_A_Valid_0_delay_42_8 <= io_A_Valid_0_delay_41_9;
    io_A_Valid_0_delay_43_7 <= io_A_Valid_0_delay_42_8;
    io_A_Valid_0_delay_44_6 <= io_A_Valid_0_delay_43_7;
    io_A_Valid_0_delay_45_5 <= io_A_Valid_0_delay_44_6;
    io_A_Valid_0_delay_46_4 <= io_A_Valid_0_delay_45_5;
    io_A_Valid_0_delay_47_3 <= io_A_Valid_0_delay_46_4;
    io_A_Valid_0_delay_48_2 <= io_A_Valid_0_delay_47_3;
    io_A_Valid_0_delay_49_1 <= io_A_Valid_0_delay_48_2;
    io_A_Valid_0_delay_50 <= io_A_Valid_0_delay_49_1;
    io_A_Valid_0_delay_1_50 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_49 <= io_A_Valid_0_delay_1_50;
    io_A_Valid_0_delay_3_48 <= io_A_Valid_0_delay_2_49;
    io_A_Valid_0_delay_4_47 <= io_A_Valid_0_delay_3_48;
    io_A_Valid_0_delay_5_46 <= io_A_Valid_0_delay_4_47;
    io_A_Valid_0_delay_6_45 <= io_A_Valid_0_delay_5_46;
    io_A_Valid_0_delay_7_44 <= io_A_Valid_0_delay_6_45;
    io_A_Valid_0_delay_8_43 <= io_A_Valid_0_delay_7_44;
    io_A_Valid_0_delay_9_42 <= io_A_Valid_0_delay_8_43;
    io_A_Valid_0_delay_10_41 <= io_A_Valid_0_delay_9_42;
    io_A_Valid_0_delay_11_40 <= io_A_Valid_0_delay_10_41;
    io_A_Valid_0_delay_12_39 <= io_A_Valid_0_delay_11_40;
    io_A_Valid_0_delay_13_38 <= io_A_Valid_0_delay_12_39;
    io_A_Valid_0_delay_14_37 <= io_A_Valid_0_delay_13_38;
    io_A_Valid_0_delay_15_36 <= io_A_Valid_0_delay_14_37;
    io_A_Valid_0_delay_16_35 <= io_A_Valid_0_delay_15_36;
    io_A_Valid_0_delay_17_34 <= io_A_Valid_0_delay_16_35;
    io_A_Valid_0_delay_18_33 <= io_A_Valid_0_delay_17_34;
    io_A_Valid_0_delay_19_32 <= io_A_Valid_0_delay_18_33;
    io_A_Valid_0_delay_20_31 <= io_A_Valid_0_delay_19_32;
    io_A_Valid_0_delay_21_30 <= io_A_Valid_0_delay_20_31;
    io_A_Valid_0_delay_22_29 <= io_A_Valid_0_delay_21_30;
    io_A_Valid_0_delay_23_28 <= io_A_Valid_0_delay_22_29;
    io_A_Valid_0_delay_24_27 <= io_A_Valid_0_delay_23_28;
    io_A_Valid_0_delay_25_26 <= io_A_Valid_0_delay_24_27;
    io_A_Valid_0_delay_26_25 <= io_A_Valid_0_delay_25_26;
    io_A_Valid_0_delay_27_24 <= io_A_Valid_0_delay_26_25;
    io_A_Valid_0_delay_28_23 <= io_A_Valid_0_delay_27_24;
    io_A_Valid_0_delay_29_22 <= io_A_Valid_0_delay_28_23;
    io_A_Valid_0_delay_30_21 <= io_A_Valid_0_delay_29_22;
    io_A_Valid_0_delay_31_20 <= io_A_Valid_0_delay_30_21;
    io_A_Valid_0_delay_32_19 <= io_A_Valid_0_delay_31_20;
    io_A_Valid_0_delay_33_18 <= io_A_Valid_0_delay_32_19;
    io_A_Valid_0_delay_34_17 <= io_A_Valid_0_delay_33_18;
    io_A_Valid_0_delay_35_16 <= io_A_Valid_0_delay_34_17;
    io_A_Valid_0_delay_36_15 <= io_A_Valid_0_delay_35_16;
    io_A_Valid_0_delay_37_14 <= io_A_Valid_0_delay_36_15;
    io_A_Valid_0_delay_38_13 <= io_A_Valid_0_delay_37_14;
    io_A_Valid_0_delay_39_12 <= io_A_Valid_0_delay_38_13;
    io_A_Valid_0_delay_40_11 <= io_A_Valid_0_delay_39_12;
    io_A_Valid_0_delay_41_10 <= io_A_Valid_0_delay_40_11;
    io_A_Valid_0_delay_42_9 <= io_A_Valid_0_delay_41_10;
    io_A_Valid_0_delay_43_8 <= io_A_Valid_0_delay_42_9;
    io_A_Valid_0_delay_44_7 <= io_A_Valid_0_delay_43_8;
    io_A_Valid_0_delay_45_6 <= io_A_Valid_0_delay_44_7;
    io_A_Valid_0_delay_46_5 <= io_A_Valid_0_delay_45_6;
    io_A_Valid_0_delay_47_4 <= io_A_Valid_0_delay_46_5;
    io_A_Valid_0_delay_48_3 <= io_A_Valid_0_delay_47_4;
    io_A_Valid_0_delay_49_2 <= io_A_Valid_0_delay_48_3;
    io_A_Valid_0_delay_50_1 <= io_A_Valid_0_delay_49_2;
    io_A_Valid_0_delay_51 <= io_A_Valid_0_delay_50_1;
    io_A_Valid_0_delay_1_51 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_50 <= io_A_Valid_0_delay_1_51;
    io_A_Valid_0_delay_3_49 <= io_A_Valid_0_delay_2_50;
    io_A_Valid_0_delay_4_48 <= io_A_Valid_0_delay_3_49;
    io_A_Valid_0_delay_5_47 <= io_A_Valid_0_delay_4_48;
    io_A_Valid_0_delay_6_46 <= io_A_Valid_0_delay_5_47;
    io_A_Valid_0_delay_7_45 <= io_A_Valid_0_delay_6_46;
    io_A_Valid_0_delay_8_44 <= io_A_Valid_0_delay_7_45;
    io_A_Valid_0_delay_9_43 <= io_A_Valid_0_delay_8_44;
    io_A_Valid_0_delay_10_42 <= io_A_Valid_0_delay_9_43;
    io_A_Valid_0_delay_11_41 <= io_A_Valid_0_delay_10_42;
    io_A_Valid_0_delay_12_40 <= io_A_Valid_0_delay_11_41;
    io_A_Valid_0_delay_13_39 <= io_A_Valid_0_delay_12_40;
    io_A_Valid_0_delay_14_38 <= io_A_Valid_0_delay_13_39;
    io_A_Valid_0_delay_15_37 <= io_A_Valid_0_delay_14_38;
    io_A_Valid_0_delay_16_36 <= io_A_Valid_0_delay_15_37;
    io_A_Valid_0_delay_17_35 <= io_A_Valid_0_delay_16_36;
    io_A_Valid_0_delay_18_34 <= io_A_Valid_0_delay_17_35;
    io_A_Valid_0_delay_19_33 <= io_A_Valid_0_delay_18_34;
    io_A_Valid_0_delay_20_32 <= io_A_Valid_0_delay_19_33;
    io_A_Valid_0_delay_21_31 <= io_A_Valid_0_delay_20_32;
    io_A_Valid_0_delay_22_30 <= io_A_Valid_0_delay_21_31;
    io_A_Valid_0_delay_23_29 <= io_A_Valid_0_delay_22_30;
    io_A_Valid_0_delay_24_28 <= io_A_Valid_0_delay_23_29;
    io_A_Valid_0_delay_25_27 <= io_A_Valid_0_delay_24_28;
    io_A_Valid_0_delay_26_26 <= io_A_Valid_0_delay_25_27;
    io_A_Valid_0_delay_27_25 <= io_A_Valid_0_delay_26_26;
    io_A_Valid_0_delay_28_24 <= io_A_Valid_0_delay_27_25;
    io_A_Valid_0_delay_29_23 <= io_A_Valid_0_delay_28_24;
    io_A_Valid_0_delay_30_22 <= io_A_Valid_0_delay_29_23;
    io_A_Valid_0_delay_31_21 <= io_A_Valid_0_delay_30_22;
    io_A_Valid_0_delay_32_20 <= io_A_Valid_0_delay_31_21;
    io_A_Valid_0_delay_33_19 <= io_A_Valid_0_delay_32_20;
    io_A_Valid_0_delay_34_18 <= io_A_Valid_0_delay_33_19;
    io_A_Valid_0_delay_35_17 <= io_A_Valid_0_delay_34_18;
    io_A_Valid_0_delay_36_16 <= io_A_Valid_0_delay_35_17;
    io_A_Valid_0_delay_37_15 <= io_A_Valid_0_delay_36_16;
    io_A_Valid_0_delay_38_14 <= io_A_Valid_0_delay_37_15;
    io_A_Valid_0_delay_39_13 <= io_A_Valid_0_delay_38_14;
    io_A_Valid_0_delay_40_12 <= io_A_Valid_0_delay_39_13;
    io_A_Valid_0_delay_41_11 <= io_A_Valid_0_delay_40_12;
    io_A_Valid_0_delay_42_10 <= io_A_Valid_0_delay_41_11;
    io_A_Valid_0_delay_43_9 <= io_A_Valid_0_delay_42_10;
    io_A_Valid_0_delay_44_8 <= io_A_Valid_0_delay_43_9;
    io_A_Valid_0_delay_45_7 <= io_A_Valid_0_delay_44_8;
    io_A_Valid_0_delay_46_6 <= io_A_Valid_0_delay_45_7;
    io_A_Valid_0_delay_47_5 <= io_A_Valid_0_delay_46_6;
    io_A_Valid_0_delay_48_4 <= io_A_Valid_0_delay_47_5;
    io_A_Valid_0_delay_49_3 <= io_A_Valid_0_delay_48_4;
    io_A_Valid_0_delay_50_2 <= io_A_Valid_0_delay_49_3;
    io_A_Valid_0_delay_51_1 <= io_A_Valid_0_delay_50_2;
    io_A_Valid_0_delay_52 <= io_A_Valid_0_delay_51_1;
    io_A_Valid_0_delay_1_52 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_51 <= io_A_Valid_0_delay_1_52;
    io_A_Valid_0_delay_3_50 <= io_A_Valid_0_delay_2_51;
    io_A_Valid_0_delay_4_49 <= io_A_Valid_0_delay_3_50;
    io_A_Valid_0_delay_5_48 <= io_A_Valid_0_delay_4_49;
    io_A_Valid_0_delay_6_47 <= io_A_Valid_0_delay_5_48;
    io_A_Valid_0_delay_7_46 <= io_A_Valid_0_delay_6_47;
    io_A_Valid_0_delay_8_45 <= io_A_Valid_0_delay_7_46;
    io_A_Valid_0_delay_9_44 <= io_A_Valid_0_delay_8_45;
    io_A_Valid_0_delay_10_43 <= io_A_Valid_0_delay_9_44;
    io_A_Valid_0_delay_11_42 <= io_A_Valid_0_delay_10_43;
    io_A_Valid_0_delay_12_41 <= io_A_Valid_0_delay_11_42;
    io_A_Valid_0_delay_13_40 <= io_A_Valid_0_delay_12_41;
    io_A_Valid_0_delay_14_39 <= io_A_Valid_0_delay_13_40;
    io_A_Valid_0_delay_15_38 <= io_A_Valid_0_delay_14_39;
    io_A_Valid_0_delay_16_37 <= io_A_Valid_0_delay_15_38;
    io_A_Valid_0_delay_17_36 <= io_A_Valid_0_delay_16_37;
    io_A_Valid_0_delay_18_35 <= io_A_Valid_0_delay_17_36;
    io_A_Valid_0_delay_19_34 <= io_A_Valid_0_delay_18_35;
    io_A_Valid_0_delay_20_33 <= io_A_Valid_0_delay_19_34;
    io_A_Valid_0_delay_21_32 <= io_A_Valid_0_delay_20_33;
    io_A_Valid_0_delay_22_31 <= io_A_Valid_0_delay_21_32;
    io_A_Valid_0_delay_23_30 <= io_A_Valid_0_delay_22_31;
    io_A_Valid_0_delay_24_29 <= io_A_Valid_0_delay_23_30;
    io_A_Valid_0_delay_25_28 <= io_A_Valid_0_delay_24_29;
    io_A_Valid_0_delay_26_27 <= io_A_Valid_0_delay_25_28;
    io_A_Valid_0_delay_27_26 <= io_A_Valid_0_delay_26_27;
    io_A_Valid_0_delay_28_25 <= io_A_Valid_0_delay_27_26;
    io_A_Valid_0_delay_29_24 <= io_A_Valid_0_delay_28_25;
    io_A_Valid_0_delay_30_23 <= io_A_Valid_0_delay_29_24;
    io_A_Valid_0_delay_31_22 <= io_A_Valid_0_delay_30_23;
    io_A_Valid_0_delay_32_21 <= io_A_Valid_0_delay_31_22;
    io_A_Valid_0_delay_33_20 <= io_A_Valid_0_delay_32_21;
    io_A_Valid_0_delay_34_19 <= io_A_Valid_0_delay_33_20;
    io_A_Valid_0_delay_35_18 <= io_A_Valid_0_delay_34_19;
    io_A_Valid_0_delay_36_17 <= io_A_Valid_0_delay_35_18;
    io_A_Valid_0_delay_37_16 <= io_A_Valid_0_delay_36_17;
    io_A_Valid_0_delay_38_15 <= io_A_Valid_0_delay_37_16;
    io_A_Valid_0_delay_39_14 <= io_A_Valid_0_delay_38_15;
    io_A_Valid_0_delay_40_13 <= io_A_Valid_0_delay_39_14;
    io_A_Valid_0_delay_41_12 <= io_A_Valid_0_delay_40_13;
    io_A_Valid_0_delay_42_11 <= io_A_Valid_0_delay_41_12;
    io_A_Valid_0_delay_43_10 <= io_A_Valid_0_delay_42_11;
    io_A_Valid_0_delay_44_9 <= io_A_Valid_0_delay_43_10;
    io_A_Valid_0_delay_45_8 <= io_A_Valid_0_delay_44_9;
    io_A_Valid_0_delay_46_7 <= io_A_Valid_0_delay_45_8;
    io_A_Valid_0_delay_47_6 <= io_A_Valid_0_delay_46_7;
    io_A_Valid_0_delay_48_5 <= io_A_Valid_0_delay_47_6;
    io_A_Valid_0_delay_49_4 <= io_A_Valid_0_delay_48_5;
    io_A_Valid_0_delay_50_3 <= io_A_Valid_0_delay_49_4;
    io_A_Valid_0_delay_51_2 <= io_A_Valid_0_delay_50_3;
    io_A_Valid_0_delay_52_1 <= io_A_Valid_0_delay_51_2;
    io_A_Valid_0_delay_53 <= io_A_Valid_0_delay_52_1;
    io_A_Valid_0_delay_1_53 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_52 <= io_A_Valid_0_delay_1_53;
    io_A_Valid_0_delay_3_51 <= io_A_Valid_0_delay_2_52;
    io_A_Valid_0_delay_4_50 <= io_A_Valid_0_delay_3_51;
    io_A_Valid_0_delay_5_49 <= io_A_Valid_0_delay_4_50;
    io_A_Valid_0_delay_6_48 <= io_A_Valid_0_delay_5_49;
    io_A_Valid_0_delay_7_47 <= io_A_Valid_0_delay_6_48;
    io_A_Valid_0_delay_8_46 <= io_A_Valid_0_delay_7_47;
    io_A_Valid_0_delay_9_45 <= io_A_Valid_0_delay_8_46;
    io_A_Valid_0_delay_10_44 <= io_A_Valid_0_delay_9_45;
    io_A_Valid_0_delay_11_43 <= io_A_Valid_0_delay_10_44;
    io_A_Valid_0_delay_12_42 <= io_A_Valid_0_delay_11_43;
    io_A_Valid_0_delay_13_41 <= io_A_Valid_0_delay_12_42;
    io_A_Valid_0_delay_14_40 <= io_A_Valid_0_delay_13_41;
    io_A_Valid_0_delay_15_39 <= io_A_Valid_0_delay_14_40;
    io_A_Valid_0_delay_16_38 <= io_A_Valid_0_delay_15_39;
    io_A_Valid_0_delay_17_37 <= io_A_Valid_0_delay_16_38;
    io_A_Valid_0_delay_18_36 <= io_A_Valid_0_delay_17_37;
    io_A_Valid_0_delay_19_35 <= io_A_Valid_0_delay_18_36;
    io_A_Valid_0_delay_20_34 <= io_A_Valid_0_delay_19_35;
    io_A_Valid_0_delay_21_33 <= io_A_Valid_0_delay_20_34;
    io_A_Valid_0_delay_22_32 <= io_A_Valid_0_delay_21_33;
    io_A_Valid_0_delay_23_31 <= io_A_Valid_0_delay_22_32;
    io_A_Valid_0_delay_24_30 <= io_A_Valid_0_delay_23_31;
    io_A_Valid_0_delay_25_29 <= io_A_Valid_0_delay_24_30;
    io_A_Valid_0_delay_26_28 <= io_A_Valid_0_delay_25_29;
    io_A_Valid_0_delay_27_27 <= io_A_Valid_0_delay_26_28;
    io_A_Valid_0_delay_28_26 <= io_A_Valid_0_delay_27_27;
    io_A_Valid_0_delay_29_25 <= io_A_Valid_0_delay_28_26;
    io_A_Valid_0_delay_30_24 <= io_A_Valid_0_delay_29_25;
    io_A_Valid_0_delay_31_23 <= io_A_Valid_0_delay_30_24;
    io_A_Valid_0_delay_32_22 <= io_A_Valid_0_delay_31_23;
    io_A_Valid_0_delay_33_21 <= io_A_Valid_0_delay_32_22;
    io_A_Valid_0_delay_34_20 <= io_A_Valid_0_delay_33_21;
    io_A_Valid_0_delay_35_19 <= io_A_Valid_0_delay_34_20;
    io_A_Valid_0_delay_36_18 <= io_A_Valid_0_delay_35_19;
    io_A_Valid_0_delay_37_17 <= io_A_Valid_0_delay_36_18;
    io_A_Valid_0_delay_38_16 <= io_A_Valid_0_delay_37_17;
    io_A_Valid_0_delay_39_15 <= io_A_Valid_0_delay_38_16;
    io_A_Valid_0_delay_40_14 <= io_A_Valid_0_delay_39_15;
    io_A_Valid_0_delay_41_13 <= io_A_Valid_0_delay_40_14;
    io_A_Valid_0_delay_42_12 <= io_A_Valid_0_delay_41_13;
    io_A_Valid_0_delay_43_11 <= io_A_Valid_0_delay_42_12;
    io_A_Valid_0_delay_44_10 <= io_A_Valid_0_delay_43_11;
    io_A_Valid_0_delay_45_9 <= io_A_Valid_0_delay_44_10;
    io_A_Valid_0_delay_46_8 <= io_A_Valid_0_delay_45_9;
    io_A_Valid_0_delay_47_7 <= io_A_Valid_0_delay_46_8;
    io_A_Valid_0_delay_48_6 <= io_A_Valid_0_delay_47_7;
    io_A_Valid_0_delay_49_5 <= io_A_Valid_0_delay_48_6;
    io_A_Valid_0_delay_50_4 <= io_A_Valid_0_delay_49_5;
    io_A_Valid_0_delay_51_3 <= io_A_Valid_0_delay_50_4;
    io_A_Valid_0_delay_52_2 <= io_A_Valid_0_delay_51_3;
    io_A_Valid_0_delay_53_1 <= io_A_Valid_0_delay_52_2;
    io_A_Valid_0_delay_54 <= io_A_Valid_0_delay_53_1;
    io_A_Valid_0_delay_1_54 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_53 <= io_A_Valid_0_delay_1_54;
    io_A_Valid_0_delay_3_52 <= io_A_Valid_0_delay_2_53;
    io_A_Valid_0_delay_4_51 <= io_A_Valid_0_delay_3_52;
    io_A_Valid_0_delay_5_50 <= io_A_Valid_0_delay_4_51;
    io_A_Valid_0_delay_6_49 <= io_A_Valid_0_delay_5_50;
    io_A_Valid_0_delay_7_48 <= io_A_Valid_0_delay_6_49;
    io_A_Valid_0_delay_8_47 <= io_A_Valid_0_delay_7_48;
    io_A_Valid_0_delay_9_46 <= io_A_Valid_0_delay_8_47;
    io_A_Valid_0_delay_10_45 <= io_A_Valid_0_delay_9_46;
    io_A_Valid_0_delay_11_44 <= io_A_Valid_0_delay_10_45;
    io_A_Valid_0_delay_12_43 <= io_A_Valid_0_delay_11_44;
    io_A_Valid_0_delay_13_42 <= io_A_Valid_0_delay_12_43;
    io_A_Valid_0_delay_14_41 <= io_A_Valid_0_delay_13_42;
    io_A_Valid_0_delay_15_40 <= io_A_Valid_0_delay_14_41;
    io_A_Valid_0_delay_16_39 <= io_A_Valid_0_delay_15_40;
    io_A_Valid_0_delay_17_38 <= io_A_Valid_0_delay_16_39;
    io_A_Valid_0_delay_18_37 <= io_A_Valid_0_delay_17_38;
    io_A_Valid_0_delay_19_36 <= io_A_Valid_0_delay_18_37;
    io_A_Valid_0_delay_20_35 <= io_A_Valid_0_delay_19_36;
    io_A_Valid_0_delay_21_34 <= io_A_Valid_0_delay_20_35;
    io_A_Valid_0_delay_22_33 <= io_A_Valid_0_delay_21_34;
    io_A_Valid_0_delay_23_32 <= io_A_Valid_0_delay_22_33;
    io_A_Valid_0_delay_24_31 <= io_A_Valid_0_delay_23_32;
    io_A_Valid_0_delay_25_30 <= io_A_Valid_0_delay_24_31;
    io_A_Valid_0_delay_26_29 <= io_A_Valid_0_delay_25_30;
    io_A_Valid_0_delay_27_28 <= io_A_Valid_0_delay_26_29;
    io_A_Valid_0_delay_28_27 <= io_A_Valid_0_delay_27_28;
    io_A_Valid_0_delay_29_26 <= io_A_Valid_0_delay_28_27;
    io_A_Valid_0_delay_30_25 <= io_A_Valid_0_delay_29_26;
    io_A_Valid_0_delay_31_24 <= io_A_Valid_0_delay_30_25;
    io_A_Valid_0_delay_32_23 <= io_A_Valid_0_delay_31_24;
    io_A_Valid_0_delay_33_22 <= io_A_Valid_0_delay_32_23;
    io_A_Valid_0_delay_34_21 <= io_A_Valid_0_delay_33_22;
    io_A_Valid_0_delay_35_20 <= io_A_Valid_0_delay_34_21;
    io_A_Valid_0_delay_36_19 <= io_A_Valid_0_delay_35_20;
    io_A_Valid_0_delay_37_18 <= io_A_Valid_0_delay_36_19;
    io_A_Valid_0_delay_38_17 <= io_A_Valid_0_delay_37_18;
    io_A_Valid_0_delay_39_16 <= io_A_Valid_0_delay_38_17;
    io_A_Valid_0_delay_40_15 <= io_A_Valid_0_delay_39_16;
    io_A_Valid_0_delay_41_14 <= io_A_Valid_0_delay_40_15;
    io_A_Valid_0_delay_42_13 <= io_A_Valid_0_delay_41_14;
    io_A_Valid_0_delay_43_12 <= io_A_Valid_0_delay_42_13;
    io_A_Valid_0_delay_44_11 <= io_A_Valid_0_delay_43_12;
    io_A_Valid_0_delay_45_10 <= io_A_Valid_0_delay_44_11;
    io_A_Valid_0_delay_46_9 <= io_A_Valid_0_delay_45_10;
    io_A_Valid_0_delay_47_8 <= io_A_Valid_0_delay_46_9;
    io_A_Valid_0_delay_48_7 <= io_A_Valid_0_delay_47_8;
    io_A_Valid_0_delay_49_6 <= io_A_Valid_0_delay_48_7;
    io_A_Valid_0_delay_50_5 <= io_A_Valid_0_delay_49_6;
    io_A_Valid_0_delay_51_4 <= io_A_Valid_0_delay_50_5;
    io_A_Valid_0_delay_52_3 <= io_A_Valid_0_delay_51_4;
    io_A_Valid_0_delay_53_2 <= io_A_Valid_0_delay_52_3;
    io_A_Valid_0_delay_54_1 <= io_A_Valid_0_delay_53_2;
    io_A_Valid_0_delay_55 <= io_A_Valid_0_delay_54_1;
    io_A_Valid_0_delay_1_55 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_54 <= io_A_Valid_0_delay_1_55;
    io_A_Valid_0_delay_3_53 <= io_A_Valid_0_delay_2_54;
    io_A_Valid_0_delay_4_52 <= io_A_Valid_0_delay_3_53;
    io_A_Valid_0_delay_5_51 <= io_A_Valid_0_delay_4_52;
    io_A_Valid_0_delay_6_50 <= io_A_Valid_0_delay_5_51;
    io_A_Valid_0_delay_7_49 <= io_A_Valid_0_delay_6_50;
    io_A_Valid_0_delay_8_48 <= io_A_Valid_0_delay_7_49;
    io_A_Valid_0_delay_9_47 <= io_A_Valid_0_delay_8_48;
    io_A_Valid_0_delay_10_46 <= io_A_Valid_0_delay_9_47;
    io_A_Valid_0_delay_11_45 <= io_A_Valid_0_delay_10_46;
    io_A_Valid_0_delay_12_44 <= io_A_Valid_0_delay_11_45;
    io_A_Valid_0_delay_13_43 <= io_A_Valid_0_delay_12_44;
    io_A_Valid_0_delay_14_42 <= io_A_Valid_0_delay_13_43;
    io_A_Valid_0_delay_15_41 <= io_A_Valid_0_delay_14_42;
    io_A_Valid_0_delay_16_40 <= io_A_Valid_0_delay_15_41;
    io_A_Valid_0_delay_17_39 <= io_A_Valid_0_delay_16_40;
    io_A_Valid_0_delay_18_38 <= io_A_Valid_0_delay_17_39;
    io_A_Valid_0_delay_19_37 <= io_A_Valid_0_delay_18_38;
    io_A_Valid_0_delay_20_36 <= io_A_Valid_0_delay_19_37;
    io_A_Valid_0_delay_21_35 <= io_A_Valid_0_delay_20_36;
    io_A_Valid_0_delay_22_34 <= io_A_Valid_0_delay_21_35;
    io_A_Valid_0_delay_23_33 <= io_A_Valid_0_delay_22_34;
    io_A_Valid_0_delay_24_32 <= io_A_Valid_0_delay_23_33;
    io_A_Valid_0_delay_25_31 <= io_A_Valid_0_delay_24_32;
    io_A_Valid_0_delay_26_30 <= io_A_Valid_0_delay_25_31;
    io_A_Valid_0_delay_27_29 <= io_A_Valid_0_delay_26_30;
    io_A_Valid_0_delay_28_28 <= io_A_Valid_0_delay_27_29;
    io_A_Valid_0_delay_29_27 <= io_A_Valid_0_delay_28_28;
    io_A_Valid_0_delay_30_26 <= io_A_Valid_0_delay_29_27;
    io_A_Valid_0_delay_31_25 <= io_A_Valid_0_delay_30_26;
    io_A_Valid_0_delay_32_24 <= io_A_Valid_0_delay_31_25;
    io_A_Valid_0_delay_33_23 <= io_A_Valid_0_delay_32_24;
    io_A_Valid_0_delay_34_22 <= io_A_Valid_0_delay_33_23;
    io_A_Valid_0_delay_35_21 <= io_A_Valid_0_delay_34_22;
    io_A_Valid_0_delay_36_20 <= io_A_Valid_0_delay_35_21;
    io_A_Valid_0_delay_37_19 <= io_A_Valid_0_delay_36_20;
    io_A_Valid_0_delay_38_18 <= io_A_Valid_0_delay_37_19;
    io_A_Valid_0_delay_39_17 <= io_A_Valid_0_delay_38_18;
    io_A_Valid_0_delay_40_16 <= io_A_Valid_0_delay_39_17;
    io_A_Valid_0_delay_41_15 <= io_A_Valid_0_delay_40_16;
    io_A_Valid_0_delay_42_14 <= io_A_Valid_0_delay_41_15;
    io_A_Valid_0_delay_43_13 <= io_A_Valid_0_delay_42_14;
    io_A_Valid_0_delay_44_12 <= io_A_Valid_0_delay_43_13;
    io_A_Valid_0_delay_45_11 <= io_A_Valid_0_delay_44_12;
    io_A_Valid_0_delay_46_10 <= io_A_Valid_0_delay_45_11;
    io_A_Valid_0_delay_47_9 <= io_A_Valid_0_delay_46_10;
    io_A_Valid_0_delay_48_8 <= io_A_Valid_0_delay_47_9;
    io_A_Valid_0_delay_49_7 <= io_A_Valid_0_delay_48_8;
    io_A_Valid_0_delay_50_6 <= io_A_Valid_0_delay_49_7;
    io_A_Valid_0_delay_51_5 <= io_A_Valid_0_delay_50_6;
    io_A_Valid_0_delay_52_4 <= io_A_Valid_0_delay_51_5;
    io_A_Valid_0_delay_53_3 <= io_A_Valid_0_delay_52_4;
    io_A_Valid_0_delay_54_2 <= io_A_Valid_0_delay_53_3;
    io_A_Valid_0_delay_55_1 <= io_A_Valid_0_delay_54_2;
    io_A_Valid_0_delay_56 <= io_A_Valid_0_delay_55_1;
    io_A_Valid_0_delay_1_56 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_55 <= io_A_Valid_0_delay_1_56;
    io_A_Valid_0_delay_3_54 <= io_A_Valid_0_delay_2_55;
    io_A_Valid_0_delay_4_53 <= io_A_Valid_0_delay_3_54;
    io_A_Valid_0_delay_5_52 <= io_A_Valid_0_delay_4_53;
    io_A_Valid_0_delay_6_51 <= io_A_Valid_0_delay_5_52;
    io_A_Valid_0_delay_7_50 <= io_A_Valid_0_delay_6_51;
    io_A_Valid_0_delay_8_49 <= io_A_Valid_0_delay_7_50;
    io_A_Valid_0_delay_9_48 <= io_A_Valid_0_delay_8_49;
    io_A_Valid_0_delay_10_47 <= io_A_Valid_0_delay_9_48;
    io_A_Valid_0_delay_11_46 <= io_A_Valid_0_delay_10_47;
    io_A_Valid_0_delay_12_45 <= io_A_Valid_0_delay_11_46;
    io_A_Valid_0_delay_13_44 <= io_A_Valid_0_delay_12_45;
    io_A_Valid_0_delay_14_43 <= io_A_Valid_0_delay_13_44;
    io_A_Valid_0_delay_15_42 <= io_A_Valid_0_delay_14_43;
    io_A_Valid_0_delay_16_41 <= io_A_Valid_0_delay_15_42;
    io_A_Valid_0_delay_17_40 <= io_A_Valid_0_delay_16_41;
    io_A_Valid_0_delay_18_39 <= io_A_Valid_0_delay_17_40;
    io_A_Valid_0_delay_19_38 <= io_A_Valid_0_delay_18_39;
    io_A_Valid_0_delay_20_37 <= io_A_Valid_0_delay_19_38;
    io_A_Valid_0_delay_21_36 <= io_A_Valid_0_delay_20_37;
    io_A_Valid_0_delay_22_35 <= io_A_Valid_0_delay_21_36;
    io_A_Valid_0_delay_23_34 <= io_A_Valid_0_delay_22_35;
    io_A_Valid_0_delay_24_33 <= io_A_Valid_0_delay_23_34;
    io_A_Valid_0_delay_25_32 <= io_A_Valid_0_delay_24_33;
    io_A_Valid_0_delay_26_31 <= io_A_Valid_0_delay_25_32;
    io_A_Valid_0_delay_27_30 <= io_A_Valid_0_delay_26_31;
    io_A_Valid_0_delay_28_29 <= io_A_Valid_0_delay_27_30;
    io_A_Valid_0_delay_29_28 <= io_A_Valid_0_delay_28_29;
    io_A_Valid_0_delay_30_27 <= io_A_Valid_0_delay_29_28;
    io_A_Valid_0_delay_31_26 <= io_A_Valid_0_delay_30_27;
    io_A_Valid_0_delay_32_25 <= io_A_Valid_0_delay_31_26;
    io_A_Valid_0_delay_33_24 <= io_A_Valid_0_delay_32_25;
    io_A_Valid_0_delay_34_23 <= io_A_Valid_0_delay_33_24;
    io_A_Valid_0_delay_35_22 <= io_A_Valid_0_delay_34_23;
    io_A_Valid_0_delay_36_21 <= io_A_Valid_0_delay_35_22;
    io_A_Valid_0_delay_37_20 <= io_A_Valid_0_delay_36_21;
    io_A_Valid_0_delay_38_19 <= io_A_Valid_0_delay_37_20;
    io_A_Valid_0_delay_39_18 <= io_A_Valid_0_delay_38_19;
    io_A_Valid_0_delay_40_17 <= io_A_Valid_0_delay_39_18;
    io_A_Valid_0_delay_41_16 <= io_A_Valid_0_delay_40_17;
    io_A_Valid_0_delay_42_15 <= io_A_Valid_0_delay_41_16;
    io_A_Valid_0_delay_43_14 <= io_A_Valid_0_delay_42_15;
    io_A_Valid_0_delay_44_13 <= io_A_Valid_0_delay_43_14;
    io_A_Valid_0_delay_45_12 <= io_A_Valid_0_delay_44_13;
    io_A_Valid_0_delay_46_11 <= io_A_Valid_0_delay_45_12;
    io_A_Valid_0_delay_47_10 <= io_A_Valid_0_delay_46_11;
    io_A_Valid_0_delay_48_9 <= io_A_Valid_0_delay_47_10;
    io_A_Valid_0_delay_49_8 <= io_A_Valid_0_delay_48_9;
    io_A_Valid_0_delay_50_7 <= io_A_Valid_0_delay_49_8;
    io_A_Valid_0_delay_51_6 <= io_A_Valid_0_delay_50_7;
    io_A_Valid_0_delay_52_5 <= io_A_Valid_0_delay_51_6;
    io_A_Valid_0_delay_53_4 <= io_A_Valid_0_delay_52_5;
    io_A_Valid_0_delay_54_3 <= io_A_Valid_0_delay_53_4;
    io_A_Valid_0_delay_55_2 <= io_A_Valid_0_delay_54_3;
    io_A_Valid_0_delay_56_1 <= io_A_Valid_0_delay_55_2;
    io_A_Valid_0_delay_57 <= io_A_Valid_0_delay_56_1;
    io_A_Valid_0_delay_1_57 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_56 <= io_A_Valid_0_delay_1_57;
    io_A_Valid_0_delay_3_55 <= io_A_Valid_0_delay_2_56;
    io_A_Valid_0_delay_4_54 <= io_A_Valid_0_delay_3_55;
    io_A_Valid_0_delay_5_53 <= io_A_Valid_0_delay_4_54;
    io_A_Valid_0_delay_6_52 <= io_A_Valid_0_delay_5_53;
    io_A_Valid_0_delay_7_51 <= io_A_Valid_0_delay_6_52;
    io_A_Valid_0_delay_8_50 <= io_A_Valid_0_delay_7_51;
    io_A_Valid_0_delay_9_49 <= io_A_Valid_0_delay_8_50;
    io_A_Valid_0_delay_10_48 <= io_A_Valid_0_delay_9_49;
    io_A_Valid_0_delay_11_47 <= io_A_Valid_0_delay_10_48;
    io_A_Valid_0_delay_12_46 <= io_A_Valid_0_delay_11_47;
    io_A_Valid_0_delay_13_45 <= io_A_Valid_0_delay_12_46;
    io_A_Valid_0_delay_14_44 <= io_A_Valid_0_delay_13_45;
    io_A_Valid_0_delay_15_43 <= io_A_Valid_0_delay_14_44;
    io_A_Valid_0_delay_16_42 <= io_A_Valid_0_delay_15_43;
    io_A_Valid_0_delay_17_41 <= io_A_Valid_0_delay_16_42;
    io_A_Valid_0_delay_18_40 <= io_A_Valid_0_delay_17_41;
    io_A_Valid_0_delay_19_39 <= io_A_Valid_0_delay_18_40;
    io_A_Valid_0_delay_20_38 <= io_A_Valid_0_delay_19_39;
    io_A_Valid_0_delay_21_37 <= io_A_Valid_0_delay_20_38;
    io_A_Valid_0_delay_22_36 <= io_A_Valid_0_delay_21_37;
    io_A_Valid_0_delay_23_35 <= io_A_Valid_0_delay_22_36;
    io_A_Valid_0_delay_24_34 <= io_A_Valid_0_delay_23_35;
    io_A_Valid_0_delay_25_33 <= io_A_Valid_0_delay_24_34;
    io_A_Valid_0_delay_26_32 <= io_A_Valid_0_delay_25_33;
    io_A_Valid_0_delay_27_31 <= io_A_Valid_0_delay_26_32;
    io_A_Valid_0_delay_28_30 <= io_A_Valid_0_delay_27_31;
    io_A_Valid_0_delay_29_29 <= io_A_Valid_0_delay_28_30;
    io_A_Valid_0_delay_30_28 <= io_A_Valid_0_delay_29_29;
    io_A_Valid_0_delay_31_27 <= io_A_Valid_0_delay_30_28;
    io_A_Valid_0_delay_32_26 <= io_A_Valid_0_delay_31_27;
    io_A_Valid_0_delay_33_25 <= io_A_Valid_0_delay_32_26;
    io_A_Valid_0_delay_34_24 <= io_A_Valid_0_delay_33_25;
    io_A_Valid_0_delay_35_23 <= io_A_Valid_0_delay_34_24;
    io_A_Valid_0_delay_36_22 <= io_A_Valid_0_delay_35_23;
    io_A_Valid_0_delay_37_21 <= io_A_Valid_0_delay_36_22;
    io_A_Valid_0_delay_38_20 <= io_A_Valid_0_delay_37_21;
    io_A_Valid_0_delay_39_19 <= io_A_Valid_0_delay_38_20;
    io_A_Valid_0_delay_40_18 <= io_A_Valid_0_delay_39_19;
    io_A_Valid_0_delay_41_17 <= io_A_Valid_0_delay_40_18;
    io_A_Valid_0_delay_42_16 <= io_A_Valid_0_delay_41_17;
    io_A_Valid_0_delay_43_15 <= io_A_Valid_0_delay_42_16;
    io_A_Valid_0_delay_44_14 <= io_A_Valid_0_delay_43_15;
    io_A_Valid_0_delay_45_13 <= io_A_Valid_0_delay_44_14;
    io_A_Valid_0_delay_46_12 <= io_A_Valid_0_delay_45_13;
    io_A_Valid_0_delay_47_11 <= io_A_Valid_0_delay_46_12;
    io_A_Valid_0_delay_48_10 <= io_A_Valid_0_delay_47_11;
    io_A_Valid_0_delay_49_9 <= io_A_Valid_0_delay_48_10;
    io_A_Valid_0_delay_50_8 <= io_A_Valid_0_delay_49_9;
    io_A_Valid_0_delay_51_7 <= io_A_Valid_0_delay_50_8;
    io_A_Valid_0_delay_52_6 <= io_A_Valid_0_delay_51_7;
    io_A_Valid_0_delay_53_5 <= io_A_Valid_0_delay_52_6;
    io_A_Valid_0_delay_54_4 <= io_A_Valid_0_delay_53_5;
    io_A_Valid_0_delay_55_3 <= io_A_Valid_0_delay_54_4;
    io_A_Valid_0_delay_56_2 <= io_A_Valid_0_delay_55_3;
    io_A_Valid_0_delay_57_1 <= io_A_Valid_0_delay_56_2;
    io_A_Valid_0_delay_58 <= io_A_Valid_0_delay_57_1;
    io_A_Valid_0_delay_1_58 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_57 <= io_A_Valid_0_delay_1_58;
    io_A_Valid_0_delay_3_56 <= io_A_Valid_0_delay_2_57;
    io_A_Valid_0_delay_4_55 <= io_A_Valid_0_delay_3_56;
    io_A_Valid_0_delay_5_54 <= io_A_Valid_0_delay_4_55;
    io_A_Valid_0_delay_6_53 <= io_A_Valid_0_delay_5_54;
    io_A_Valid_0_delay_7_52 <= io_A_Valid_0_delay_6_53;
    io_A_Valid_0_delay_8_51 <= io_A_Valid_0_delay_7_52;
    io_A_Valid_0_delay_9_50 <= io_A_Valid_0_delay_8_51;
    io_A_Valid_0_delay_10_49 <= io_A_Valid_0_delay_9_50;
    io_A_Valid_0_delay_11_48 <= io_A_Valid_0_delay_10_49;
    io_A_Valid_0_delay_12_47 <= io_A_Valid_0_delay_11_48;
    io_A_Valid_0_delay_13_46 <= io_A_Valid_0_delay_12_47;
    io_A_Valid_0_delay_14_45 <= io_A_Valid_0_delay_13_46;
    io_A_Valid_0_delay_15_44 <= io_A_Valid_0_delay_14_45;
    io_A_Valid_0_delay_16_43 <= io_A_Valid_0_delay_15_44;
    io_A_Valid_0_delay_17_42 <= io_A_Valid_0_delay_16_43;
    io_A_Valid_0_delay_18_41 <= io_A_Valid_0_delay_17_42;
    io_A_Valid_0_delay_19_40 <= io_A_Valid_0_delay_18_41;
    io_A_Valid_0_delay_20_39 <= io_A_Valid_0_delay_19_40;
    io_A_Valid_0_delay_21_38 <= io_A_Valid_0_delay_20_39;
    io_A_Valid_0_delay_22_37 <= io_A_Valid_0_delay_21_38;
    io_A_Valid_0_delay_23_36 <= io_A_Valid_0_delay_22_37;
    io_A_Valid_0_delay_24_35 <= io_A_Valid_0_delay_23_36;
    io_A_Valid_0_delay_25_34 <= io_A_Valid_0_delay_24_35;
    io_A_Valid_0_delay_26_33 <= io_A_Valid_0_delay_25_34;
    io_A_Valid_0_delay_27_32 <= io_A_Valid_0_delay_26_33;
    io_A_Valid_0_delay_28_31 <= io_A_Valid_0_delay_27_32;
    io_A_Valid_0_delay_29_30 <= io_A_Valid_0_delay_28_31;
    io_A_Valid_0_delay_30_29 <= io_A_Valid_0_delay_29_30;
    io_A_Valid_0_delay_31_28 <= io_A_Valid_0_delay_30_29;
    io_A_Valid_0_delay_32_27 <= io_A_Valid_0_delay_31_28;
    io_A_Valid_0_delay_33_26 <= io_A_Valid_0_delay_32_27;
    io_A_Valid_0_delay_34_25 <= io_A_Valid_0_delay_33_26;
    io_A_Valid_0_delay_35_24 <= io_A_Valid_0_delay_34_25;
    io_A_Valid_0_delay_36_23 <= io_A_Valid_0_delay_35_24;
    io_A_Valid_0_delay_37_22 <= io_A_Valid_0_delay_36_23;
    io_A_Valid_0_delay_38_21 <= io_A_Valid_0_delay_37_22;
    io_A_Valid_0_delay_39_20 <= io_A_Valid_0_delay_38_21;
    io_A_Valid_0_delay_40_19 <= io_A_Valid_0_delay_39_20;
    io_A_Valid_0_delay_41_18 <= io_A_Valid_0_delay_40_19;
    io_A_Valid_0_delay_42_17 <= io_A_Valid_0_delay_41_18;
    io_A_Valid_0_delay_43_16 <= io_A_Valid_0_delay_42_17;
    io_A_Valid_0_delay_44_15 <= io_A_Valid_0_delay_43_16;
    io_A_Valid_0_delay_45_14 <= io_A_Valid_0_delay_44_15;
    io_A_Valid_0_delay_46_13 <= io_A_Valid_0_delay_45_14;
    io_A_Valid_0_delay_47_12 <= io_A_Valid_0_delay_46_13;
    io_A_Valid_0_delay_48_11 <= io_A_Valid_0_delay_47_12;
    io_A_Valid_0_delay_49_10 <= io_A_Valid_0_delay_48_11;
    io_A_Valid_0_delay_50_9 <= io_A_Valid_0_delay_49_10;
    io_A_Valid_0_delay_51_8 <= io_A_Valid_0_delay_50_9;
    io_A_Valid_0_delay_52_7 <= io_A_Valid_0_delay_51_8;
    io_A_Valid_0_delay_53_6 <= io_A_Valid_0_delay_52_7;
    io_A_Valid_0_delay_54_5 <= io_A_Valid_0_delay_53_6;
    io_A_Valid_0_delay_55_4 <= io_A_Valid_0_delay_54_5;
    io_A_Valid_0_delay_56_3 <= io_A_Valid_0_delay_55_4;
    io_A_Valid_0_delay_57_2 <= io_A_Valid_0_delay_56_3;
    io_A_Valid_0_delay_58_1 <= io_A_Valid_0_delay_57_2;
    io_A_Valid_0_delay_59 <= io_A_Valid_0_delay_58_1;
    io_A_Valid_0_delay_1_59 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_58 <= io_A_Valid_0_delay_1_59;
    io_A_Valid_0_delay_3_57 <= io_A_Valid_0_delay_2_58;
    io_A_Valid_0_delay_4_56 <= io_A_Valid_0_delay_3_57;
    io_A_Valid_0_delay_5_55 <= io_A_Valid_0_delay_4_56;
    io_A_Valid_0_delay_6_54 <= io_A_Valid_0_delay_5_55;
    io_A_Valid_0_delay_7_53 <= io_A_Valid_0_delay_6_54;
    io_A_Valid_0_delay_8_52 <= io_A_Valid_0_delay_7_53;
    io_A_Valid_0_delay_9_51 <= io_A_Valid_0_delay_8_52;
    io_A_Valid_0_delay_10_50 <= io_A_Valid_0_delay_9_51;
    io_A_Valid_0_delay_11_49 <= io_A_Valid_0_delay_10_50;
    io_A_Valid_0_delay_12_48 <= io_A_Valid_0_delay_11_49;
    io_A_Valid_0_delay_13_47 <= io_A_Valid_0_delay_12_48;
    io_A_Valid_0_delay_14_46 <= io_A_Valid_0_delay_13_47;
    io_A_Valid_0_delay_15_45 <= io_A_Valid_0_delay_14_46;
    io_A_Valid_0_delay_16_44 <= io_A_Valid_0_delay_15_45;
    io_A_Valid_0_delay_17_43 <= io_A_Valid_0_delay_16_44;
    io_A_Valid_0_delay_18_42 <= io_A_Valid_0_delay_17_43;
    io_A_Valid_0_delay_19_41 <= io_A_Valid_0_delay_18_42;
    io_A_Valid_0_delay_20_40 <= io_A_Valid_0_delay_19_41;
    io_A_Valid_0_delay_21_39 <= io_A_Valid_0_delay_20_40;
    io_A_Valid_0_delay_22_38 <= io_A_Valid_0_delay_21_39;
    io_A_Valid_0_delay_23_37 <= io_A_Valid_0_delay_22_38;
    io_A_Valid_0_delay_24_36 <= io_A_Valid_0_delay_23_37;
    io_A_Valid_0_delay_25_35 <= io_A_Valid_0_delay_24_36;
    io_A_Valid_0_delay_26_34 <= io_A_Valid_0_delay_25_35;
    io_A_Valid_0_delay_27_33 <= io_A_Valid_0_delay_26_34;
    io_A_Valid_0_delay_28_32 <= io_A_Valid_0_delay_27_33;
    io_A_Valid_0_delay_29_31 <= io_A_Valid_0_delay_28_32;
    io_A_Valid_0_delay_30_30 <= io_A_Valid_0_delay_29_31;
    io_A_Valid_0_delay_31_29 <= io_A_Valid_0_delay_30_30;
    io_A_Valid_0_delay_32_28 <= io_A_Valid_0_delay_31_29;
    io_A_Valid_0_delay_33_27 <= io_A_Valid_0_delay_32_28;
    io_A_Valid_0_delay_34_26 <= io_A_Valid_0_delay_33_27;
    io_A_Valid_0_delay_35_25 <= io_A_Valid_0_delay_34_26;
    io_A_Valid_0_delay_36_24 <= io_A_Valid_0_delay_35_25;
    io_A_Valid_0_delay_37_23 <= io_A_Valid_0_delay_36_24;
    io_A_Valid_0_delay_38_22 <= io_A_Valid_0_delay_37_23;
    io_A_Valid_0_delay_39_21 <= io_A_Valid_0_delay_38_22;
    io_A_Valid_0_delay_40_20 <= io_A_Valid_0_delay_39_21;
    io_A_Valid_0_delay_41_19 <= io_A_Valid_0_delay_40_20;
    io_A_Valid_0_delay_42_18 <= io_A_Valid_0_delay_41_19;
    io_A_Valid_0_delay_43_17 <= io_A_Valid_0_delay_42_18;
    io_A_Valid_0_delay_44_16 <= io_A_Valid_0_delay_43_17;
    io_A_Valid_0_delay_45_15 <= io_A_Valid_0_delay_44_16;
    io_A_Valid_0_delay_46_14 <= io_A_Valid_0_delay_45_15;
    io_A_Valid_0_delay_47_13 <= io_A_Valid_0_delay_46_14;
    io_A_Valid_0_delay_48_12 <= io_A_Valid_0_delay_47_13;
    io_A_Valid_0_delay_49_11 <= io_A_Valid_0_delay_48_12;
    io_A_Valid_0_delay_50_10 <= io_A_Valid_0_delay_49_11;
    io_A_Valid_0_delay_51_9 <= io_A_Valid_0_delay_50_10;
    io_A_Valid_0_delay_52_8 <= io_A_Valid_0_delay_51_9;
    io_A_Valid_0_delay_53_7 <= io_A_Valid_0_delay_52_8;
    io_A_Valid_0_delay_54_6 <= io_A_Valid_0_delay_53_7;
    io_A_Valid_0_delay_55_5 <= io_A_Valid_0_delay_54_6;
    io_A_Valid_0_delay_56_4 <= io_A_Valid_0_delay_55_5;
    io_A_Valid_0_delay_57_3 <= io_A_Valid_0_delay_56_4;
    io_A_Valid_0_delay_58_2 <= io_A_Valid_0_delay_57_3;
    io_A_Valid_0_delay_59_1 <= io_A_Valid_0_delay_58_2;
    io_A_Valid_0_delay_60 <= io_A_Valid_0_delay_59_1;
    io_A_Valid_0_delay_1_60 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_59 <= io_A_Valid_0_delay_1_60;
    io_A_Valid_0_delay_3_58 <= io_A_Valid_0_delay_2_59;
    io_A_Valid_0_delay_4_57 <= io_A_Valid_0_delay_3_58;
    io_A_Valid_0_delay_5_56 <= io_A_Valid_0_delay_4_57;
    io_A_Valid_0_delay_6_55 <= io_A_Valid_0_delay_5_56;
    io_A_Valid_0_delay_7_54 <= io_A_Valid_0_delay_6_55;
    io_A_Valid_0_delay_8_53 <= io_A_Valid_0_delay_7_54;
    io_A_Valid_0_delay_9_52 <= io_A_Valid_0_delay_8_53;
    io_A_Valid_0_delay_10_51 <= io_A_Valid_0_delay_9_52;
    io_A_Valid_0_delay_11_50 <= io_A_Valid_0_delay_10_51;
    io_A_Valid_0_delay_12_49 <= io_A_Valid_0_delay_11_50;
    io_A_Valid_0_delay_13_48 <= io_A_Valid_0_delay_12_49;
    io_A_Valid_0_delay_14_47 <= io_A_Valid_0_delay_13_48;
    io_A_Valid_0_delay_15_46 <= io_A_Valid_0_delay_14_47;
    io_A_Valid_0_delay_16_45 <= io_A_Valid_0_delay_15_46;
    io_A_Valid_0_delay_17_44 <= io_A_Valid_0_delay_16_45;
    io_A_Valid_0_delay_18_43 <= io_A_Valid_0_delay_17_44;
    io_A_Valid_0_delay_19_42 <= io_A_Valid_0_delay_18_43;
    io_A_Valid_0_delay_20_41 <= io_A_Valid_0_delay_19_42;
    io_A_Valid_0_delay_21_40 <= io_A_Valid_0_delay_20_41;
    io_A_Valid_0_delay_22_39 <= io_A_Valid_0_delay_21_40;
    io_A_Valid_0_delay_23_38 <= io_A_Valid_0_delay_22_39;
    io_A_Valid_0_delay_24_37 <= io_A_Valid_0_delay_23_38;
    io_A_Valid_0_delay_25_36 <= io_A_Valid_0_delay_24_37;
    io_A_Valid_0_delay_26_35 <= io_A_Valid_0_delay_25_36;
    io_A_Valid_0_delay_27_34 <= io_A_Valid_0_delay_26_35;
    io_A_Valid_0_delay_28_33 <= io_A_Valid_0_delay_27_34;
    io_A_Valid_0_delay_29_32 <= io_A_Valid_0_delay_28_33;
    io_A_Valid_0_delay_30_31 <= io_A_Valid_0_delay_29_32;
    io_A_Valid_0_delay_31_30 <= io_A_Valid_0_delay_30_31;
    io_A_Valid_0_delay_32_29 <= io_A_Valid_0_delay_31_30;
    io_A_Valid_0_delay_33_28 <= io_A_Valid_0_delay_32_29;
    io_A_Valid_0_delay_34_27 <= io_A_Valid_0_delay_33_28;
    io_A_Valid_0_delay_35_26 <= io_A_Valid_0_delay_34_27;
    io_A_Valid_0_delay_36_25 <= io_A_Valid_0_delay_35_26;
    io_A_Valid_0_delay_37_24 <= io_A_Valid_0_delay_36_25;
    io_A_Valid_0_delay_38_23 <= io_A_Valid_0_delay_37_24;
    io_A_Valid_0_delay_39_22 <= io_A_Valid_0_delay_38_23;
    io_A_Valid_0_delay_40_21 <= io_A_Valid_0_delay_39_22;
    io_A_Valid_0_delay_41_20 <= io_A_Valid_0_delay_40_21;
    io_A_Valid_0_delay_42_19 <= io_A_Valid_0_delay_41_20;
    io_A_Valid_0_delay_43_18 <= io_A_Valid_0_delay_42_19;
    io_A_Valid_0_delay_44_17 <= io_A_Valid_0_delay_43_18;
    io_A_Valid_0_delay_45_16 <= io_A_Valid_0_delay_44_17;
    io_A_Valid_0_delay_46_15 <= io_A_Valid_0_delay_45_16;
    io_A_Valid_0_delay_47_14 <= io_A_Valid_0_delay_46_15;
    io_A_Valid_0_delay_48_13 <= io_A_Valid_0_delay_47_14;
    io_A_Valid_0_delay_49_12 <= io_A_Valid_0_delay_48_13;
    io_A_Valid_0_delay_50_11 <= io_A_Valid_0_delay_49_12;
    io_A_Valid_0_delay_51_10 <= io_A_Valid_0_delay_50_11;
    io_A_Valid_0_delay_52_9 <= io_A_Valid_0_delay_51_10;
    io_A_Valid_0_delay_53_8 <= io_A_Valid_0_delay_52_9;
    io_A_Valid_0_delay_54_7 <= io_A_Valid_0_delay_53_8;
    io_A_Valid_0_delay_55_6 <= io_A_Valid_0_delay_54_7;
    io_A_Valid_0_delay_56_5 <= io_A_Valid_0_delay_55_6;
    io_A_Valid_0_delay_57_4 <= io_A_Valid_0_delay_56_5;
    io_A_Valid_0_delay_58_3 <= io_A_Valid_0_delay_57_4;
    io_A_Valid_0_delay_59_2 <= io_A_Valid_0_delay_58_3;
    io_A_Valid_0_delay_60_1 <= io_A_Valid_0_delay_59_2;
    io_A_Valid_0_delay_61 <= io_A_Valid_0_delay_60_1;
    io_A_Valid_0_delay_1_61 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_60 <= io_A_Valid_0_delay_1_61;
    io_A_Valid_0_delay_3_59 <= io_A_Valid_0_delay_2_60;
    io_A_Valid_0_delay_4_58 <= io_A_Valid_0_delay_3_59;
    io_A_Valid_0_delay_5_57 <= io_A_Valid_0_delay_4_58;
    io_A_Valid_0_delay_6_56 <= io_A_Valid_0_delay_5_57;
    io_A_Valid_0_delay_7_55 <= io_A_Valid_0_delay_6_56;
    io_A_Valid_0_delay_8_54 <= io_A_Valid_0_delay_7_55;
    io_A_Valid_0_delay_9_53 <= io_A_Valid_0_delay_8_54;
    io_A_Valid_0_delay_10_52 <= io_A_Valid_0_delay_9_53;
    io_A_Valid_0_delay_11_51 <= io_A_Valid_0_delay_10_52;
    io_A_Valid_0_delay_12_50 <= io_A_Valid_0_delay_11_51;
    io_A_Valid_0_delay_13_49 <= io_A_Valid_0_delay_12_50;
    io_A_Valid_0_delay_14_48 <= io_A_Valid_0_delay_13_49;
    io_A_Valid_0_delay_15_47 <= io_A_Valid_0_delay_14_48;
    io_A_Valid_0_delay_16_46 <= io_A_Valid_0_delay_15_47;
    io_A_Valid_0_delay_17_45 <= io_A_Valid_0_delay_16_46;
    io_A_Valid_0_delay_18_44 <= io_A_Valid_0_delay_17_45;
    io_A_Valid_0_delay_19_43 <= io_A_Valid_0_delay_18_44;
    io_A_Valid_0_delay_20_42 <= io_A_Valid_0_delay_19_43;
    io_A_Valid_0_delay_21_41 <= io_A_Valid_0_delay_20_42;
    io_A_Valid_0_delay_22_40 <= io_A_Valid_0_delay_21_41;
    io_A_Valid_0_delay_23_39 <= io_A_Valid_0_delay_22_40;
    io_A_Valid_0_delay_24_38 <= io_A_Valid_0_delay_23_39;
    io_A_Valid_0_delay_25_37 <= io_A_Valid_0_delay_24_38;
    io_A_Valid_0_delay_26_36 <= io_A_Valid_0_delay_25_37;
    io_A_Valid_0_delay_27_35 <= io_A_Valid_0_delay_26_36;
    io_A_Valid_0_delay_28_34 <= io_A_Valid_0_delay_27_35;
    io_A_Valid_0_delay_29_33 <= io_A_Valid_0_delay_28_34;
    io_A_Valid_0_delay_30_32 <= io_A_Valid_0_delay_29_33;
    io_A_Valid_0_delay_31_31 <= io_A_Valid_0_delay_30_32;
    io_A_Valid_0_delay_32_30 <= io_A_Valid_0_delay_31_31;
    io_A_Valid_0_delay_33_29 <= io_A_Valid_0_delay_32_30;
    io_A_Valid_0_delay_34_28 <= io_A_Valid_0_delay_33_29;
    io_A_Valid_0_delay_35_27 <= io_A_Valid_0_delay_34_28;
    io_A_Valid_0_delay_36_26 <= io_A_Valid_0_delay_35_27;
    io_A_Valid_0_delay_37_25 <= io_A_Valid_0_delay_36_26;
    io_A_Valid_0_delay_38_24 <= io_A_Valid_0_delay_37_25;
    io_A_Valid_0_delay_39_23 <= io_A_Valid_0_delay_38_24;
    io_A_Valid_0_delay_40_22 <= io_A_Valid_0_delay_39_23;
    io_A_Valid_0_delay_41_21 <= io_A_Valid_0_delay_40_22;
    io_A_Valid_0_delay_42_20 <= io_A_Valid_0_delay_41_21;
    io_A_Valid_0_delay_43_19 <= io_A_Valid_0_delay_42_20;
    io_A_Valid_0_delay_44_18 <= io_A_Valid_0_delay_43_19;
    io_A_Valid_0_delay_45_17 <= io_A_Valid_0_delay_44_18;
    io_A_Valid_0_delay_46_16 <= io_A_Valid_0_delay_45_17;
    io_A_Valid_0_delay_47_15 <= io_A_Valid_0_delay_46_16;
    io_A_Valid_0_delay_48_14 <= io_A_Valid_0_delay_47_15;
    io_A_Valid_0_delay_49_13 <= io_A_Valid_0_delay_48_14;
    io_A_Valid_0_delay_50_12 <= io_A_Valid_0_delay_49_13;
    io_A_Valid_0_delay_51_11 <= io_A_Valid_0_delay_50_12;
    io_A_Valid_0_delay_52_10 <= io_A_Valid_0_delay_51_11;
    io_A_Valid_0_delay_53_9 <= io_A_Valid_0_delay_52_10;
    io_A_Valid_0_delay_54_8 <= io_A_Valid_0_delay_53_9;
    io_A_Valid_0_delay_55_7 <= io_A_Valid_0_delay_54_8;
    io_A_Valid_0_delay_56_6 <= io_A_Valid_0_delay_55_7;
    io_A_Valid_0_delay_57_5 <= io_A_Valid_0_delay_56_6;
    io_A_Valid_0_delay_58_4 <= io_A_Valid_0_delay_57_5;
    io_A_Valid_0_delay_59_3 <= io_A_Valid_0_delay_58_4;
    io_A_Valid_0_delay_60_2 <= io_A_Valid_0_delay_59_3;
    io_A_Valid_0_delay_61_1 <= io_A_Valid_0_delay_60_2;
    io_A_Valid_0_delay_62 <= io_A_Valid_0_delay_61_1;
    io_A_Valid_0_delay_1_62 <= io_A_Valid_0;
    io_A_Valid_0_delay_2_61 <= io_A_Valid_0_delay_1_62;
    io_A_Valid_0_delay_3_60 <= io_A_Valid_0_delay_2_61;
    io_A_Valid_0_delay_4_59 <= io_A_Valid_0_delay_3_60;
    io_A_Valid_0_delay_5_58 <= io_A_Valid_0_delay_4_59;
    io_A_Valid_0_delay_6_57 <= io_A_Valid_0_delay_5_58;
    io_A_Valid_0_delay_7_56 <= io_A_Valid_0_delay_6_57;
    io_A_Valid_0_delay_8_55 <= io_A_Valid_0_delay_7_56;
    io_A_Valid_0_delay_9_54 <= io_A_Valid_0_delay_8_55;
    io_A_Valid_0_delay_10_53 <= io_A_Valid_0_delay_9_54;
    io_A_Valid_0_delay_11_52 <= io_A_Valid_0_delay_10_53;
    io_A_Valid_0_delay_12_51 <= io_A_Valid_0_delay_11_52;
    io_A_Valid_0_delay_13_50 <= io_A_Valid_0_delay_12_51;
    io_A_Valid_0_delay_14_49 <= io_A_Valid_0_delay_13_50;
    io_A_Valid_0_delay_15_48 <= io_A_Valid_0_delay_14_49;
    io_A_Valid_0_delay_16_47 <= io_A_Valid_0_delay_15_48;
    io_A_Valid_0_delay_17_46 <= io_A_Valid_0_delay_16_47;
    io_A_Valid_0_delay_18_45 <= io_A_Valid_0_delay_17_46;
    io_A_Valid_0_delay_19_44 <= io_A_Valid_0_delay_18_45;
    io_A_Valid_0_delay_20_43 <= io_A_Valid_0_delay_19_44;
    io_A_Valid_0_delay_21_42 <= io_A_Valid_0_delay_20_43;
    io_A_Valid_0_delay_22_41 <= io_A_Valid_0_delay_21_42;
    io_A_Valid_0_delay_23_40 <= io_A_Valid_0_delay_22_41;
    io_A_Valid_0_delay_24_39 <= io_A_Valid_0_delay_23_40;
    io_A_Valid_0_delay_25_38 <= io_A_Valid_0_delay_24_39;
    io_A_Valid_0_delay_26_37 <= io_A_Valid_0_delay_25_38;
    io_A_Valid_0_delay_27_36 <= io_A_Valid_0_delay_26_37;
    io_A_Valid_0_delay_28_35 <= io_A_Valid_0_delay_27_36;
    io_A_Valid_0_delay_29_34 <= io_A_Valid_0_delay_28_35;
    io_A_Valid_0_delay_30_33 <= io_A_Valid_0_delay_29_34;
    io_A_Valid_0_delay_31_32 <= io_A_Valid_0_delay_30_33;
    io_A_Valid_0_delay_32_31 <= io_A_Valid_0_delay_31_32;
    io_A_Valid_0_delay_33_30 <= io_A_Valid_0_delay_32_31;
    io_A_Valid_0_delay_34_29 <= io_A_Valid_0_delay_33_30;
    io_A_Valid_0_delay_35_28 <= io_A_Valid_0_delay_34_29;
    io_A_Valid_0_delay_36_27 <= io_A_Valid_0_delay_35_28;
    io_A_Valid_0_delay_37_26 <= io_A_Valid_0_delay_36_27;
    io_A_Valid_0_delay_38_25 <= io_A_Valid_0_delay_37_26;
    io_A_Valid_0_delay_39_24 <= io_A_Valid_0_delay_38_25;
    io_A_Valid_0_delay_40_23 <= io_A_Valid_0_delay_39_24;
    io_A_Valid_0_delay_41_22 <= io_A_Valid_0_delay_40_23;
    io_A_Valid_0_delay_42_21 <= io_A_Valid_0_delay_41_22;
    io_A_Valid_0_delay_43_20 <= io_A_Valid_0_delay_42_21;
    io_A_Valid_0_delay_44_19 <= io_A_Valid_0_delay_43_20;
    io_A_Valid_0_delay_45_18 <= io_A_Valid_0_delay_44_19;
    io_A_Valid_0_delay_46_17 <= io_A_Valid_0_delay_45_18;
    io_A_Valid_0_delay_47_16 <= io_A_Valid_0_delay_46_17;
    io_A_Valid_0_delay_48_15 <= io_A_Valid_0_delay_47_16;
    io_A_Valid_0_delay_49_14 <= io_A_Valid_0_delay_48_15;
    io_A_Valid_0_delay_50_13 <= io_A_Valid_0_delay_49_14;
    io_A_Valid_0_delay_51_12 <= io_A_Valid_0_delay_50_13;
    io_A_Valid_0_delay_52_11 <= io_A_Valid_0_delay_51_12;
    io_A_Valid_0_delay_53_10 <= io_A_Valid_0_delay_52_11;
    io_A_Valid_0_delay_54_9 <= io_A_Valid_0_delay_53_10;
    io_A_Valid_0_delay_55_8 <= io_A_Valid_0_delay_54_9;
    io_A_Valid_0_delay_56_7 <= io_A_Valid_0_delay_55_8;
    io_A_Valid_0_delay_57_6 <= io_A_Valid_0_delay_56_7;
    io_A_Valid_0_delay_58_5 <= io_A_Valid_0_delay_57_6;
    io_A_Valid_0_delay_59_4 <= io_A_Valid_0_delay_58_5;
    io_A_Valid_0_delay_60_3 <= io_A_Valid_0_delay_59_4;
    io_A_Valid_0_delay_61_2 <= io_A_Valid_0_delay_60_3;
    io_A_Valid_0_delay_62_1 <= io_A_Valid_0_delay_61_2;
    io_A_Valid_0_delay_63 <= io_A_Valid_0_delay_62_1;
    io_B_Valid_0_delay_1 <= io_B_Valid_0;
    io_A_Valid_1_delay_1 <= io_A_Valid_1;
    io_B_Valid_1_delay_1 <= io_B_Valid_1;
    io_A_Valid_1_delay_1_1 <= io_A_Valid_1;
    io_A_Valid_1_delay_2 <= io_A_Valid_1_delay_1_1;
    io_B_Valid_2_delay_1 <= io_B_Valid_2;
    io_A_Valid_1_delay_1_2 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_1 <= io_A_Valid_1_delay_1_2;
    io_A_Valid_1_delay_3 <= io_A_Valid_1_delay_2_1;
    io_B_Valid_3_delay_1 <= io_B_Valid_3;
    io_A_Valid_1_delay_1_3 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_2 <= io_A_Valid_1_delay_1_3;
    io_A_Valid_1_delay_3_1 <= io_A_Valid_1_delay_2_2;
    io_A_Valid_1_delay_4 <= io_A_Valid_1_delay_3_1;
    io_B_Valid_4_delay_1 <= io_B_Valid_4;
    io_A_Valid_1_delay_1_4 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_3 <= io_A_Valid_1_delay_1_4;
    io_A_Valid_1_delay_3_2 <= io_A_Valid_1_delay_2_3;
    io_A_Valid_1_delay_4_1 <= io_A_Valid_1_delay_3_2;
    io_A_Valid_1_delay_5 <= io_A_Valid_1_delay_4_1;
    io_B_Valid_5_delay_1 <= io_B_Valid_5;
    io_A_Valid_1_delay_1_5 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_4 <= io_A_Valid_1_delay_1_5;
    io_A_Valid_1_delay_3_3 <= io_A_Valid_1_delay_2_4;
    io_A_Valid_1_delay_4_2 <= io_A_Valid_1_delay_3_3;
    io_A_Valid_1_delay_5_1 <= io_A_Valid_1_delay_4_2;
    io_A_Valid_1_delay_6 <= io_A_Valid_1_delay_5_1;
    io_B_Valid_6_delay_1 <= io_B_Valid_6;
    io_A_Valid_1_delay_1_6 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_5 <= io_A_Valid_1_delay_1_6;
    io_A_Valid_1_delay_3_4 <= io_A_Valid_1_delay_2_5;
    io_A_Valid_1_delay_4_3 <= io_A_Valid_1_delay_3_4;
    io_A_Valid_1_delay_5_2 <= io_A_Valid_1_delay_4_3;
    io_A_Valid_1_delay_6_1 <= io_A_Valid_1_delay_5_2;
    io_A_Valid_1_delay_7 <= io_A_Valid_1_delay_6_1;
    io_B_Valid_7_delay_1 <= io_B_Valid_7;
    io_A_Valid_1_delay_1_7 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_6 <= io_A_Valid_1_delay_1_7;
    io_A_Valid_1_delay_3_5 <= io_A_Valid_1_delay_2_6;
    io_A_Valid_1_delay_4_4 <= io_A_Valid_1_delay_3_5;
    io_A_Valid_1_delay_5_3 <= io_A_Valid_1_delay_4_4;
    io_A_Valid_1_delay_6_2 <= io_A_Valid_1_delay_5_3;
    io_A_Valid_1_delay_7_1 <= io_A_Valid_1_delay_6_2;
    io_A_Valid_1_delay_8 <= io_A_Valid_1_delay_7_1;
    io_B_Valid_8_delay_1 <= io_B_Valid_8;
    io_A_Valid_1_delay_1_8 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_7 <= io_A_Valid_1_delay_1_8;
    io_A_Valid_1_delay_3_6 <= io_A_Valid_1_delay_2_7;
    io_A_Valid_1_delay_4_5 <= io_A_Valid_1_delay_3_6;
    io_A_Valid_1_delay_5_4 <= io_A_Valid_1_delay_4_5;
    io_A_Valid_1_delay_6_3 <= io_A_Valid_1_delay_5_4;
    io_A_Valid_1_delay_7_2 <= io_A_Valid_1_delay_6_3;
    io_A_Valid_1_delay_8_1 <= io_A_Valid_1_delay_7_2;
    io_A_Valid_1_delay_9 <= io_A_Valid_1_delay_8_1;
    io_B_Valid_9_delay_1 <= io_B_Valid_9;
    io_A_Valid_1_delay_1_9 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_8 <= io_A_Valid_1_delay_1_9;
    io_A_Valid_1_delay_3_7 <= io_A_Valid_1_delay_2_8;
    io_A_Valid_1_delay_4_6 <= io_A_Valid_1_delay_3_7;
    io_A_Valid_1_delay_5_5 <= io_A_Valid_1_delay_4_6;
    io_A_Valid_1_delay_6_4 <= io_A_Valid_1_delay_5_5;
    io_A_Valid_1_delay_7_3 <= io_A_Valid_1_delay_6_4;
    io_A_Valid_1_delay_8_2 <= io_A_Valid_1_delay_7_3;
    io_A_Valid_1_delay_9_1 <= io_A_Valid_1_delay_8_2;
    io_A_Valid_1_delay_10 <= io_A_Valid_1_delay_9_1;
    io_B_Valid_10_delay_1 <= io_B_Valid_10;
    io_A_Valid_1_delay_1_10 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_9 <= io_A_Valid_1_delay_1_10;
    io_A_Valid_1_delay_3_8 <= io_A_Valid_1_delay_2_9;
    io_A_Valid_1_delay_4_7 <= io_A_Valid_1_delay_3_8;
    io_A_Valid_1_delay_5_6 <= io_A_Valid_1_delay_4_7;
    io_A_Valid_1_delay_6_5 <= io_A_Valid_1_delay_5_6;
    io_A_Valid_1_delay_7_4 <= io_A_Valid_1_delay_6_5;
    io_A_Valid_1_delay_8_3 <= io_A_Valid_1_delay_7_4;
    io_A_Valid_1_delay_9_2 <= io_A_Valid_1_delay_8_3;
    io_A_Valid_1_delay_10_1 <= io_A_Valid_1_delay_9_2;
    io_A_Valid_1_delay_11 <= io_A_Valid_1_delay_10_1;
    io_B_Valid_11_delay_1 <= io_B_Valid_11;
    io_A_Valid_1_delay_1_11 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_10 <= io_A_Valid_1_delay_1_11;
    io_A_Valid_1_delay_3_9 <= io_A_Valid_1_delay_2_10;
    io_A_Valid_1_delay_4_8 <= io_A_Valid_1_delay_3_9;
    io_A_Valid_1_delay_5_7 <= io_A_Valid_1_delay_4_8;
    io_A_Valid_1_delay_6_6 <= io_A_Valid_1_delay_5_7;
    io_A_Valid_1_delay_7_5 <= io_A_Valid_1_delay_6_6;
    io_A_Valid_1_delay_8_4 <= io_A_Valid_1_delay_7_5;
    io_A_Valid_1_delay_9_3 <= io_A_Valid_1_delay_8_4;
    io_A_Valid_1_delay_10_2 <= io_A_Valid_1_delay_9_3;
    io_A_Valid_1_delay_11_1 <= io_A_Valid_1_delay_10_2;
    io_A_Valid_1_delay_12 <= io_A_Valid_1_delay_11_1;
    io_B_Valid_12_delay_1 <= io_B_Valid_12;
    io_A_Valid_1_delay_1_12 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_11 <= io_A_Valid_1_delay_1_12;
    io_A_Valid_1_delay_3_10 <= io_A_Valid_1_delay_2_11;
    io_A_Valid_1_delay_4_9 <= io_A_Valid_1_delay_3_10;
    io_A_Valid_1_delay_5_8 <= io_A_Valid_1_delay_4_9;
    io_A_Valid_1_delay_6_7 <= io_A_Valid_1_delay_5_8;
    io_A_Valid_1_delay_7_6 <= io_A_Valid_1_delay_6_7;
    io_A_Valid_1_delay_8_5 <= io_A_Valid_1_delay_7_6;
    io_A_Valid_1_delay_9_4 <= io_A_Valid_1_delay_8_5;
    io_A_Valid_1_delay_10_3 <= io_A_Valid_1_delay_9_4;
    io_A_Valid_1_delay_11_2 <= io_A_Valid_1_delay_10_3;
    io_A_Valid_1_delay_12_1 <= io_A_Valid_1_delay_11_2;
    io_A_Valid_1_delay_13 <= io_A_Valid_1_delay_12_1;
    io_B_Valid_13_delay_1 <= io_B_Valid_13;
    io_A_Valid_1_delay_1_13 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_12 <= io_A_Valid_1_delay_1_13;
    io_A_Valid_1_delay_3_11 <= io_A_Valid_1_delay_2_12;
    io_A_Valid_1_delay_4_10 <= io_A_Valid_1_delay_3_11;
    io_A_Valid_1_delay_5_9 <= io_A_Valid_1_delay_4_10;
    io_A_Valid_1_delay_6_8 <= io_A_Valid_1_delay_5_9;
    io_A_Valid_1_delay_7_7 <= io_A_Valid_1_delay_6_8;
    io_A_Valid_1_delay_8_6 <= io_A_Valid_1_delay_7_7;
    io_A_Valid_1_delay_9_5 <= io_A_Valid_1_delay_8_6;
    io_A_Valid_1_delay_10_4 <= io_A_Valid_1_delay_9_5;
    io_A_Valid_1_delay_11_3 <= io_A_Valid_1_delay_10_4;
    io_A_Valid_1_delay_12_2 <= io_A_Valid_1_delay_11_3;
    io_A_Valid_1_delay_13_1 <= io_A_Valid_1_delay_12_2;
    io_A_Valid_1_delay_14 <= io_A_Valid_1_delay_13_1;
    io_B_Valid_14_delay_1 <= io_B_Valid_14;
    io_A_Valid_1_delay_1_14 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_13 <= io_A_Valid_1_delay_1_14;
    io_A_Valid_1_delay_3_12 <= io_A_Valid_1_delay_2_13;
    io_A_Valid_1_delay_4_11 <= io_A_Valid_1_delay_3_12;
    io_A_Valid_1_delay_5_10 <= io_A_Valid_1_delay_4_11;
    io_A_Valid_1_delay_6_9 <= io_A_Valid_1_delay_5_10;
    io_A_Valid_1_delay_7_8 <= io_A_Valid_1_delay_6_9;
    io_A_Valid_1_delay_8_7 <= io_A_Valid_1_delay_7_8;
    io_A_Valid_1_delay_9_6 <= io_A_Valid_1_delay_8_7;
    io_A_Valid_1_delay_10_5 <= io_A_Valid_1_delay_9_6;
    io_A_Valid_1_delay_11_4 <= io_A_Valid_1_delay_10_5;
    io_A_Valid_1_delay_12_3 <= io_A_Valid_1_delay_11_4;
    io_A_Valid_1_delay_13_2 <= io_A_Valid_1_delay_12_3;
    io_A_Valid_1_delay_14_1 <= io_A_Valid_1_delay_13_2;
    io_A_Valid_1_delay_15 <= io_A_Valid_1_delay_14_1;
    io_B_Valid_15_delay_1 <= io_B_Valid_15;
    io_A_Valid_1_delay_1_15 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_14 <= io_A_Valid_1_delay_1_15;
    io_A_Valid_1_delay_3_13 <= io_A_Valid_1_delay_2_14;
    io_A_Valid_1_delay_4_12 <= io_A_Valid_1_delay_3_13;
    io_A_Valid_1_delay_5_11 <= io_A_Valid_1_delay_4_12;
    io_A_Valid_1_delay_6_10 <= io_A_Valid_1_delay_5_11;
    io_A_Valid_1_delay_7_9 <= io_A_Valid_1_delay_6_10;
    io_A_Valid_1_delay_8_8 <= io_A_Valid_1_delay_7_9;
    io_A_Valid_1_delay_9_7 <= io_A_Valid_1_delay_8_8;
    io_A_Valid_1_delay_10_6 <= io_A_Valid_1_delay_9_7;
    io_A_Valid_1_delay_11_5 <= io_A_Valid_1_delay_10_6;
    io_A_Valid_1_delay_12_4 <= io_A_Valid_1_delay_11_5;
    io_A_Valid_1_delay_13_3 <= io_A_Valid_1_delay_12_4;
    io_A_Valid_1_delay_14_2 <= io_A_Valid_1_delay_13_3;
    io_A_Valid_1_delay_15_1 <= io_A_Valid_1_delay_14_2;
    io_A_Valid_1_delay_16 <= io_A_Valid_1_delay_15_1;
    io_B_Valid_16_delay_1 <= io_B_Valid_16;
    io_A_Valid_1_delay_1_16 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_15 <= io_A_Valid_1_delay_1_16;
    io_A_Valid_1_delay_3_14 <= io_A_Valid_1_delay_2_15;
    io_A_Valid_1_delay_4_13 <= io_A_Valid_1_delay_3_14;
    io_A_Valid_1_delay_5_12 <= io_A_Valid_1_delay_4_13;
    io_A_Valid_1_delay_6_11 <= io_A_Valid_1_delay_5_12;
    io_A_Valid_1_delay_7_10 <= io_A_Valid_1_delay_6_11;
    io_A_Valid_1_delay_8_9 <= io_A_Valid_1_delay_7_10;
    io_A_Valid_1_delay_9_8 <= io_A_Valid_1_delay_8_9;
    io_A_Valid_1_delay_10_7 <= io_A_Valid_1_delay_9_8;
    io_A_Valid_1_delay_11_6 <= io_A_Valid_1_delay_10_7;
    io_A_Valid_1_delay_12_5 <= io_A_Valid_1_delay_11_6;
    io_A_Valid_1_delay_13_4 <= io_A_Valid_1_delay_12_5;
    io_A_Valid_1_delay_14_3 <= io_A_Valid_1_delay_13_4;
    io_A_Valid_1_delay_15_2 <= io_A_Valid_1_delay_14_3;
    io_A_Valid_1_delay_16_1 <= io_A_Valid_1_delay_15_2;
    io_A_Valid_1_delay_17 <= io_A_Valid_1_delay_16_1;
    io_B_Valid_17_delay_1 <= io_B_Valid_17;
    io_A_Valid_1_delay_1_17 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_16 <= io_A_Valid_1_delay_1_17;
    io_A_Valid_1_delay_3_15 <= io_A_Valid_1_delay_2_16;
    io_A_Valid_1_delay_4_14 <= io_A_Valid_1_delay_3_15;
    io_A_Valid_1_delay_5_13 <= io_A_Valid_1_delay_4_14;
    io_A_Valid_1_delay_6_12 <= io_A_Valid_1_delay_5_13;
    io_A_Valid_1_delay_7_11 <= io_A_Valid_1_delay_6_12;
    io_A_Valid_1_delay_8_10 <= io_A_Valid_1_delay_7_11;
    io_A_Valid_1_delay_9_9 <= io_A_Valid_1_delay_8_10;
    io_A_Valid_1_delay_10_8 <= io_A_Valid_1_delay_9_9;
    io_A_Valid_1_delay_11_7 <= io_A_Valid_1_delay_10_8;
    io_A_Valid_1_delay_12_6 <= io_A_Valid_1_delay_11_7;
    io_A_Valid_1_delay_13_5 <= io_A_Valid_1_delay_12_6;
    io_A_Valid_1_delay_14_4 <= io_A_Valid_1_delay_13_5;
    io_A_Valid_1_delay_15_3 <= io_A_Valid_1_delay_14_4;
    io_A_Valid_1_delay_16_2 <= io_A_Valid_1_delay_15_3;
    io_A_Valid_1_delay_17_1 <= io_A_Valid_1_delay_16_2;
    io_A_Valid_1_delay_18 <= io_A_Valid_1_delay_17_1;
    io_B_Valid_18_delay_1 <= io_B_Valid_18;
    io_A_Valid_1_delay_1_18 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_17 <= io_A_Valid_1_delay_1_18;
    io_A_Valid_1_delay_3_16 <= io_A_Valid_1_delay_2_17;
    io_A_Valid_1_delay_4_15 <= io_A_Valid_1_delay_3_16;
    io_A_Valid_1_delay_5_14 <= io_A_Valid_1_delay_4_15;
    io_A_Valid_1_delay_6_13 <= io_A_Valid_1_delay_5_14;
    io_A_Valid_1_delay_7_12 <= io_A_Valid_1_delay_6_13;
    io_A_Valid_1_delay_8_11 <= io_A_Valid_1_delay_7_12;
    io_A_Valid_1_delay_9_10 <= io_A_Valid_1_delay_8_11;
    io_A_Valid_1_delay_10_9 <= io_A_Valid_1_delay_9_10;
    io_A_Valid_1_delay_11_8 <= io_A_Valid_1_delay_10_9;
    io_A_Valid_1_delay_12_7 <= io_A_Valid_1_delay_11_8;
    io_A_Valid_1_delay_13_6 <= io_A_Valid_1_delay_12_7;
    io_A_Valid_1_delay_14_5 <= io_A_Valid_1_delay_13_6;
    io_A_Valid_1_delay_15_4 <= io_A_Valid_1_delay_14_5;
    io_A_Valid_1_delay_16_3 <= io_A_Valid_1_delay_15_4;
    io_A_Valid_1_delay_17_2 <= io_A_Valid_1_delay_16_3;
    io_A_Valid_1_delay_18_1 <= io_A_Valid_1_delay_17_2;
    io_A_Valid_1_delay_19 <= io_A_Valid_1_delay_18_1;
    io_B_Valid_19_delay_1 <= io_B_Valid_19;
    io_A_Valid_1_delay_1_19 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_18 <= io_A_Valid_1_delay_1_19;
    io_A_Valid_1_delay_3_17 <= io_A_Valid_1_delay_2_18;
    io_A_Valid_1_delay_4_16 <= io_A_Valid_1_delay_3_17;
    io_A_Valid_1_delay_5_15 <= io_A_Valid_1_delay_4_16;
    io_A_Valid_1_delay_6_14 <= io_A_Valid_1_delay_5_15;
    io_A_Valid_1_delay_7_13 <= io_A_Valid_1_delay_6_14;
    io_A_Valid_1_delay_8_12 <= io_A_Valid_1_delay_7_13;
    io_A_Valid_1_delay_9_11 <= io_A_Valid_1_delay_8_12;
    io_A_Valid_1_delay_10_10 <= io_A_Valid_1_delay_9_11;
    io_A_Valid_1_delay_11_9 <= io_A_Valid_1_delay_10_10;
    io_A_Valid_1_delay_12_8 <= io_A_Valid_1_delay_11_9;
    io_A_Valid_1_delay_13_7 <= io_A_Valid_1_delay_12_8;
    io_A_Valid_1_delay_14_6 <= io_A_Valid_1_delay_13_7;
    io_A_Valid_1_delay_15_5 <= io_A_Valid_1_delay_14_6;
    io_A_Valid_1_delay_16_4 <= io_A_Valid_1_delay_15_5;
    io_A_Valid_1_delay_17_3 <= io_A_Valid_1_delay_16_4;
    io_A_Valid_1_delay_18_2 <= io_A_Valid_1_delay_17_3;
    io_A_Valid_1_delay_19_1 <= io_A_Valid_1_delay_18_2;
    io_A_Valid_1_delay_20 <= io_A_Valid_1_delay_19_1;
    io_B_Valid_20_delay_1 <= io_B_Valid_20;
    io_A_Valid_1_delay_1_20 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_19 <= io_A_Valid_1_delay_1_20;
    io_A_Valid_1_delay_3_18 <= io_A_Valid_1_delay_2_19;
    io_A_Valid_1_delay_4_17 <= io_A_Valid_1_delay_3_18;
    io_A_Valid_1_delay_5_16 <= io_A_Valid_1_delay_4_17;
    io_A_Valid_1_delay_6_15 <= io_A_Valid_1_delay_5_16;
    io_A_Valid_1_delay_7_14 <= io_A_Valid_1_delay_6_15;
    io_A_Valid_1_delay_8_13 <= io_A_Valid_1_delay_7_14;
    io_A_Valid_1_delay_9_12 <= io_A_Valid_1_delay_8_13;
    io_A_Valid_1_delay_10_11 <= io_A_Valid_1_delay_9_12;
    io_A_Valid_1_delay_11_10 <= io_A_Valid_1_delay_10_11;
    io_A_Valid_1_delay_12_9 <= io_A_Valid_1_delay_11_10;
    io_A_Valid_1_delay_13_8 <= io_A_Valid_1_delay_12_9;
    io_A_Valid_1_delay_14_7 <= io_A_Valid_1_delay_13_8;
    io_A_Valid_1_delay_15_6 <= io_A_Valid_1_delay_14_7;
    io_A_Valid_1_delay_16_5 <= io_A_Valid_1_delay_15_6;
    io_A_Valid_1_delay_17_4 <= io_A_Valid_1_delay_16_5;
    io_A_Valid_1_delay_18_3 <= io_A_Valid_1_delay_17_4;
    io_A_Valid_1_delay_19_2 <= io_A_Valid_1_delay_18_3;
    io_A_Valid_1_delay_20_1 <= io_A_Valid_1_delay_19_2;
    io_A_Valid_1_delay_21 <= io_A_Valid_1_delay_20_1;
    io_B_Valid_21_delay_1 <= io_B_Valid_21;
    io_A_Valid_1_delay_1_21 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_20 <= io_A_Valid_1_delay_1_21;
    io_A_Valid_1_delay_3_19 <= io_A_Valid_1_delay_2_20;
    io_A_Valid_1_delay_4_18 <= io_A_Valid_1_delay_3_19;
    io_A_Valid_1_delay_5_17 <= io_A_Valid_1_delay_4_18;
    io_A_Valid_1_delay_6_16 <= io_A_Valid_1_delay_5_17;
    io_A_Valid_1_delay_7_15 <= io_A_Valid_1_delay_6_16;
    io_A_Valid_1_delay_8_14 <= io_A_Valid_1_delay_7_15;
    io_A_Valid_1_delay_9_13 <= io_A_Valid_1_delay_8_14;
    io_A_Valid_1_delay_10_12 <= io_A_Valid_1_delay_9_13;
    io_A_Valid_1_delay_11_11 <= io_A_Valid_1_delay_10_12;
    io_A_Valid_1_delay_12_10 <= io_A_Valid_1_delay_11_11;
    io_A_Valid_1_delay_13_9 <= io_A_Valid_1_delay_12_10;
    io_A_Valid_1_delay_14_8 <= io_A_Valid_1_delay_13_9;
    io_A_Valid_1_delay_15_7 <= io_A_Valid_1_delay_14_8;
    io_A_Valid_1_delay_16_6 <= io_A_Valid_1_delay_15_7;
    io_A_Valid_1_delay_17_5 <= io_A_Valid_1_delay_16_6;
    io_A_Valid_1_delay_18_4 <= io_A_Valid_1_delay_17_5;
    io_A_Valid_1_delay_19_3 <= io_A_Valid_1_delay_18_4;
    io_A_Valid_1_delay_20_2 <= io_A_Valid_1_delay_19_3;
    io_A_Valid_1_delay_21_1 <= io_A_Valid_1_delay_20_2;
    io_A_Valid_1_delay_22 <= io_A_Valid_1_delay_21_1;
    io_B_Valid_22_delay_1 <= io_B_Valid_22;
    io_A_Valid_1_delay_1_22 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_21 <= io_A_Valid_1_delay_1_22;
    io_A_Valid_1_delay_3_20 <= io_A_Valid_1_delay_2_21;
    io_A_Valid_1_delay_4_19 <= io_A_Valid_1_delay_3_20;
    io_A_Valid_1_delay_5_18 <= io_A_Valid_1_delay_4_19;
    io_A_Valid_1_delay_6_17 <= io_A_Valid_1_delay_5_18;
    io_A_Valid_1_delay_7_16 <= io_A_Valid_1_delay_6_17;
    io_A_Valid_1_delay_8_15 <= io_A_Valid_1_delay_7_16;
    io_A_Valid_1_delay_9_14 <= io_A_Valid_1_delay_8_15;
    io_A_Valid_1_delay_10_13 <= io_A_Valid_1_delay_9_14;
    io_A_Valid_1_delay_11_12 <= io_A_Valid_1_delay_10_13;
    io_A_Valid_1_delay_12_11 <= io_A_Valid_1_delay_11_12;
    io_A_Valid_1_delay_13_10 <= io_A_Valid_1_delay_12_11;
    io_A_Valid_1_delay_14_9 <= io_A_Valid_1_delay_13_10;
    io_A_Valid_1_delay_15_8 <= io_A_Valid_1_delay_14_9;
    io_A_Valid_1_delay_16_7 <= io_A_Valid_1_delay_15_8;
    io_A_Valid_1_delay_17_6 <= io_A_Valid_1_delay_16_7;
    io_A_Valid_1_delay_18_5 <= io_A_Valid_1_delay_17_6;
    io_A_Valid_1_delay_19_4 <= io_A_Valid_1_delay_18_5;
    io_A_Valid_1_delay_20_3 <= io_A_Valid_1_delay_19_4;
    io_A_Valid_1_delay_21_2 <= io_A_Valid_1_delay_20_3;
    io_A_Valid_1_delay_22_1 <= io_A_Valid_1_delay_21_2;
    io_A_Valid_1_delay_23 <= io_A_Valid_1_delay_22_1;
    io_B_Valid_23_delay_1 <= io_B_Valid_23;
    io_A_Valid_1_delay_1_23 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_22 <= io_A_Valid_1_delay_1_23;
    io_A_Valid_1_delay_3_21 <= io_A_Valid_1_delay_2_22;
    io_A_Valid_1_delay_4_20 <= io_A_Valid_1_delay_3_21;
    io_A_Valid_1_delay_5_19 <= io_A_Valid_1_delay_4_20;
    io_A_Valid_1_delay_6_18 <= io_A_Valid_1_delay_5_19;
    io_A_Valid_1_delay_7_17 <= io_A_Valid_1_delay_6_18;
    io_A_Valid_1_delay_8_16 <= io_A_Valid_1_delay_7_17;
    io_A_Valid_1_delay_9_15 <= io_A_Valid_1_delay_8_16;
    io_A_Valid_1_delay_10_14 <= io_A_Valid_1_delay_9_15;
    io_A_Valid_1_delay_11_13 <= io_A_Valid_1_delay_10_14;
    io_A_Valid_1_delay_12_12 <= io_A_Valid_1_delay_11_13;
    io_A_Valid_1_delay_13_11 <= io_A_Valid_1_delay_12_12;
    io_A_Valid_1_delay_14_10 <= io_A_Valid_1_delay_13_11;
    io_A_Valid_1_delay_15_9 <= io_A_Valid_1_delay_14_10;
    io_A_Valid_1_delay_16_8 <= io_A_Valid_1_delay_15_9;
    io_A_Valid_1_delay_17_7 <= io_A_Valid_1_delay_16_8;
    io_A_Valid_1_delay_18_6 <= io_A_Valid_1_delay_17_7;
    io_A_Valid_1_delay_19_5 <= io_A_Valid_1_delay_18_6;
    io_A_Valid_1_delay_20_4 <= io_A_Valid_1_delay_19_5;
    io_A_Valid_1_delay_21_3 <= io_A_Valid_1_delay_20_4;
    io_A_Valid_1_delay_22_2 <= io_A_Valid_1_delay_21_3;
    io_A_Valid_1_delay_23_1 <= io_A_Valid_1_delay_22_2;
    io_A_Valid_1_delay_24 <= io_A_Valid_1_delay_23_1;
    io_B_Valid_24_delay_1 <= io_B_Valid_24;
    io_A_Valid_1_delay_1_24 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_23 <= io_A_Valid_1_delay_1_24;
    io_A_Valid_1_delay_3_22 <= io_A_Valid_1_delay_2_23;
    io_A_Valid_1_delay_4_21 <= io_A_Valid_1_delay_3_22;
    io_A_Valid_1_delay_5_20 <= io_A_Valid_1_delay_4_21;
    io_A_Valid_1_delay_6_19 <= io_A_Valid_1_delay_5_20;
    io_A_Valid_1_delay_7_18 <= io_A_Valid_1_delay_6_19;
    io_A_Valid_1_delay_8_17 <= io_A_Valid_1_delay_7_18;
    io_A_Valid_1_delay_9_16 <= io_A_Valid_1_delay_8_17;
    io_A_Valid_1_delay_10_15 <= io_A_Valid_1_delay_9_16;
    io_A_Valid_1_delay_11_14 <= io_A_Valid_1_delay_10_15;
    io_A_Valid_1_delay_12_13 <= io_A_Valid_1_delay_11_14;
    io_A_Valid_1_delay_13_12 <= io_A_Valid_1_delay_12_13;
    io_A_Valid_1_delay_14_11 <= io_A_Valid_1_delay_13_12;
    io_A_Valid_1_delay_15_10 <= io_A_Valid_1_delay_14_11;
    io_A_Valid_1_delay_16_9 <= io_A_Valid_1_delay_15_10;
    io_A_Valid_1_delay_17_8 <= io_A_Valid_1_delay_16_9;
    io_A_Valid_1_delay_18_7 <= io_A_Valid_1_delay_17_8;
    io_A_Valid_1_delay_19_6 <= io_A_Valid_1_delay_18_7;
    io_A_Valid_1_delay_20_5 <= io_A_Valid_1_delay_19_6;
    io_A_Valid_1_delay_21_4 <= io_A_Valid_1_delay_20_5;
    io_A_Valid_1_delay_22_3 <= io_A_Valid_1_delay_21_4;
    io_A_Valid_1_delay_23_2 <= io_A_Valid_1_delay_22_3;
    io_A_Valid_1_delay_24_1 <= io_A_Valid_1_delay_23_2;
    io_A_Valid_1_delay_25 <= io_A_Valid_1_delay_24_1;
    io_B_Valid_25_delay_1 <= io_B_Valid_25;
    io_A_Valid_1_delay_1_25 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_24 <= io_A_Valid_1_delay_1_25;
    io_A_Valid_1_delay_3_23 <= io_A_Valid_1_delay_2_24;
    io_A_Valid_1_delay_4_22 <= io_A_Valid_1_delay_3_23;
    io_A_Valid_1_delay_5_21 <= io_A_Valid_1_delay_4_22;
    io_A_Valid_1_delay_6_20 <= io_A_Valid_1_delay_5_21;
    io_A_Valid_1_delay_7_19 <= io_A_Valid_1_delay_6_20;
    io_A_Valid_1_delay_8_18 <= io_A_Valid_1_delay_7_19;
    io_A_Valid_1_delay_9_17 <= io_A_Valid_1_delay_8_18;
    io_A_Valid_1_delay_10_16 <= io_A_Valid_1_delay_9_17;
    io_A_Valid_1_delay_11_15 <= io_A_Valid_1_delay_10_16;
    io_A_Valid_1_delay_12_14 <= io_A_Valid_1_delay_11_15;
    io_A_Valid_1_delay_13_13 <= io_A_Valid_1_delay_12_14;
    io_A_Valid_1_delay_14_12 <= io_A_Valid_1_delay_13_13;
    io_A_Valid_1_delay_15_11 <= io_A_Valid_1_delay_14_12;
    io_A_Valid_1_delay_16_10 <= io_A_Valid_1_delay_15_11;
    io_A_Valid_1_delay_17_9 <= io_A_Valid_1_delay_16_10;
    io_A_Valid_1_delay_18_8 <= io_A_Valid_1_delay_17_9;
    io_A_Valid_1_delay_19_7 <= io_A_Valid_1_delay_18_8;
    io_A_Valid_1_delay_20_6 <= io_A_Valid_1_delay_19_7;
    io_A_Valid_1_delay_21_5 <= io_A_Valid_1_delay_20_6;
    io_A_Valid_1_delay_22_4 <= io_A_Valid_1_delay_21_5;
    io_A_Valid_1_delay_23_3 <= io_A_Valid_1_delay_22_4;
    io_A_Valid_1_delay_24_2 <= io_A_Valid_1_delay_23_3;
    io_A_Valid_1_delay_25_1 <= io_A_Valid_1_delay_24_2;
    io_A_Valid_1_delay_26 <= io_A_Valid_1_delay_25_1;
    io_B_Valid_26_delay_1 <= io_B_Valid_26;
    io_A_Valid_1_delay_1_26 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_25 <= io_A_Valid_1_delay_1_26;
    io_A_Valid_1_delay_3_24 <= io_A_Valid_1_delay_2_25;
    io_A_Valid_1_delay_4_23 <= io_A_Valid_1_delay_3_24;
    io_A_Valid_1_delay_5_22 <= io_A_Valid_1_delay_4_23;
    io_A_Valid_1_delay_6_21 <= io_A_Valid_1_delay_5_22;
    io_A_Valid_1_delay_7_20 <= io_A_Valid_1_delay_6_21;
    io_A_Valid_1_delay_8_19 <= io_A_Valid_1_delay_7_20;
    io_A_Valid_1_delay_9_18 <= io_A_Valid_1_delay_8_19;
    io_A_Valid_1_delay_10_17 <= io_A_Valid_1_delay_9_18;
    io_A_Valid_1_delay_11_16 <= io_A_Valid_1_delay_10_17;
    io_A_Valid_1_delay_12_15 <= io_A_Valid_1_delay_11_16;
    io_A_Valid_1_delay_13_14 <= io_A_Valid_1_delay_12_15;
    io_A_Valid_1_delay_14_13 <= io_A_Valid_1_delay_13_14;
    io_A_Valid_1_delay_15_12 <= io_A_Valid_1_delay_14_13;
    io_A_Valid_1_delay_16_11 <= io_A_Valid_1_delay_15_12;
    io_A_Valid_1_delay_17_10 <= io_A_Valid_1_delay_16_11;
    io_A_Valid_1_delay_18_9 <= io_A_Valid_1_delay_17_10;
    io_A_Valid_1_delay_19_8 <= io_A_Valid_1_delay_18_9;
    io_A_Valid_1_delay_20_7 <= io_A_Valid_1_delay_19_8;
    io_A_Valid_1_delay_21_6 <= io_A_Valid_1_delay_20_7;
    io_A_Valid_1_delay_22_5 <= io_A_Valid_1_delay_21_6;
    io_A_Valid_1_delay_23_4 <= io_A_Valid_1_delay_22_5;
    io_A_Valid_1_delay_24_3 <= io_A_Valid_1_delay_23_4;
    io_A_Valid_1_delay_25_2 <= io_A_Valid_1_delay_24_3;
    io_A_Valid_1_delay_26_1 <= io_A_Valid_1_delay_25_2;
    io_A_Valid_1_delay_27 <= io_A_Valid_1_delay_26_1;
    io_B_Valid_27_delay_1 <= io_B_Valid_27;
    io_A_Valid_1_delay_1_27 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_26 <= io_A_Valid_1_delay_1_27;
    io_A_Valid_1_delay_3_25 <= io_A_Valid_1_delay_2_26;
    io_A_Valid_1_delay_4_24 <= io_A_Valid_1_delay_3_25;
    io_A_Valid_1_delay_5_23 <= io_A_Valid_1_delay_4_24;
    io_A_Valid_1_delay_6_22 <= io_A_Valid_1_delay_5_23;
    io_A_Valid_1_delay_7_21 <= io_A_Valid_1_delay_6_22;
    io_A_Valid_1_delay_8_20 <= io_A_Valid_1_delay_7_21;
    io_A_Valid_1_delay_9_19 <= io_A_Valid_1_delay_8_20;
    io_A_Valid_1_delay_10_18 <= io_A_Valid_1_delay_9_19;
    io_A_Valid_1_delay_11_17 <= io_A_Valid_1_delay_10_18;
    io_A_Valid_1_delay_12_16 <= io_A_Valid_1_delay_11_17;
    io_A_Valid_1_delay_13_15 <= io_A_Valid_1_delay_12_16;
    io_A_Valid_1_delay_14_14 <= io_A_Valid_1_delay_13_15;
    io_A_Valid_1_delay_15_13 <= io_A_Valid_1_delay_14_14;
    io_A_Valid_1_delay_16_12 <= io_A_Valid_1_delay_15_13;
    io_A_Valid_1_delay_17_11 <= io_A_Valid_1_delay_16_12;
    io_A_Valid_1_delay_18_10 <= io_A_Valid_1_delay_17_11;
    io_A_Valid_1_delay_19_9 <= io_A_Valid_1_delay_18_10;
    io_A_Valid_1_delay_20_8 <= io_A_Valid_1_delay_19_9;
    io_A_Valid_1_delay_21_7 <= io_A_Valid_1_delay_20_8;
    io_A_Valid_1_delay_22_6 <= io_A_Valid_1_delay_21_7;
    io_A_Valid_1_delay_23_5 <= io_A_Valid_1_delay_22_6;
    io_A_Valid_1_delay_24_4 <= io_A_Valid_1_delay_23_5;
    io_A_Valid_1_delay_25_3 <= io_A_Valid_1_delay_24_4;
    io_A_Valid_1_delay_26_2 <= io_A_Valid_1_delay_25_3;
    io_A_Valid_1_delay_27_1 <= io_A_Valid_1_delay_26_2;
    io_A_Valid_1_delay_28 <= io_A_Valid_1_delay_27_1;
    io_B_Valid_28_delay_1 <= io_B_Valid_28;
    io_A_Valid_1_delay_1_28 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_27 <= io_A_Valid_1_delay_1_28;
    io_A_Valid_1_delay_3_26 <= io_A_Valid_1_delay_2_27;
    io_A_Valid_1_delay_4_25 <= io_A_Valid_1_delay_3_26;
    io_A_Valid_1_delay_5_24 <= io_A_Valid_1_delay_4_25;
    io_A_Valid_1_delay_6_23 <= io_A_Valid_1_delay_5_24;
    io_A_Valid_1_delay_7_22 <= io_A_Valid_1_delay_6_23;
    io_A_Valid_1_delay_8_21 <= io_A_Valid_1_delay_7_22;
    io_A_Valid_1_delay_9_20 <= io_A_Valid_1_delay_8_21;
    io_A_Valid_1_delay_10_19 <= io_A_Valid_1_delay_9_20;
    io_A_Valid_1_delay_11_18 <= io_A_Valid_1_delay_10_19;
    io_A_Valid_1_delay_12_17 <= io_A_Valid_1_delay_11_18;
    io_A_Valid_1_delay_13_16 <= io_A_Valid_1_delay_12_17;
    io_A_Valid_1_delay_14_15 <= io_A_Valid_1_delay_13_16;
    io_A_Valid_1_delay_15_14 <= io_A_Valid_1_delay_14_15;
    io_A_Valid_1_delay_16_13 <= io_A_Valid_1_delay_15_14;
    io_A_Valid_1_delay_17_12 <= io_A_Valid_1_delay_16_13;
    io_A_Valid_1_delay_18_11 <= io_A_Valid_1_delay_17_12;
    io_A_Valid_1_delay_19_10 <= io_A_Valid_1_delay_18_11;
    io_A_Valid_1_delay_20_9 <= io_A_Valid_1_delay_19_10;
    io_A_Valid_1_delay_21_8 <= io_A_Valid_1_delay_20_9;
    io_A_Valid_1_delay_22_7 <= io_A_Valid_1_delay_21_8;
    io_A_Valid_1_delay_23_6 <= io_A_Valid_1_delay_22_7;
    io_A_Valid_1_delay_24_5 <= io_A_Valid_1_delay_23_6;
    io_A_Valid_1_delay_25_4 <= io_A_Valid_1_delay_24_5;
    io_A_Valid_1_delay_26_3 <= io_A_Valid_1_delay_25_4;
    io_A_Valid_1_delay_27_2 <= io_A_Valid_1_delay_26_3;
    io_A_Valid_1_delay_28_1 <= io_A_Valid_1_delay_27_2;
    io_A_Valid_1_delay_29 <= io_A_Valid_1_delay_28_1;
    io_B_Valid_29_delay_1 <= io_B_Valid_29;
    io_A_Valid_1_delay_1_29 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_28 <= io_A_Valid_1_delay_1_29;
    io_A_Valid_1_delay_3_27 <= io_A_Valid_1_delay_2_28;
    io_A_Valid_1_delay_4_26 <= io_A_Valid_1_delay_3_27;
    io_A_Valid_1_delay_5_25 <= io_A_Valid_1_delay_4_26;
    io_A_Valid_1_delay_6_24 <= io_A_Valid_1_delay_5_25;
    io_A_Valid_1_delay_7_23 <= io_A_Valid_1_delay_6_24;
    io_A_Valid_1_delay_8_22 <= io_A_Valid_1_delay_7_23;
    io_A_Valid_1_delay_9_21 <= io_A_Valid_1_delay_8_22;
    io_A_Valid_1_delay_10_20 <= io_A_Valid_1_delay_9_21;
    io_A_Valid_1_delay_11_19 <= io_A_Valid_1_delay_10_20;
    io_A_Valid_1_delay_12_18 <= io_A_Valid_1_delay_11_19;
    io_A_Valid_1_delay_13_17 <= io_A_Valid_1_delay_12_18;
    io_A_Valid_1_delay_14_16 <= io_A_Valid_1_delay_13_17;
    io_A_Valid_1_delay_15_15 <= io_A_Valid_1_delay_14_16;
    io_A_Valid_1_delay_16_14 <= io_A_Valid_1_delay_15_15;
    io_A_Valid_1_delay_17_13 <= io_A_Valid_1_delay_16_14;
    io_A_Valid_1_delay_18_12 <= io_A_Valid_1_delay_17_13;
    io_A_Valid_1_delay_19_11 <= io_A_Valid_1_delay_18_12;
    io_A_Valid_1_delay_20_10 <= io_A_Valid_1_delay_19_11;
    io_A_Valid_1_delay_21_9 <= io_A_Valid_1_delay_20_10;
    io_A_Valid_1_delay_22_8 <= io_A_Valid_1_delay_21_9;
    io_A_Valid_1_delay_23_7 <= io_A_Valid_1_delay_22_8;
    io_A_Valid_1_delay_24_6 <= io_A_Valid_1_delay_23_7;
    io_A_Valid_1_delay_25_5 <= io_A_Valid_1_delay_24_6;
    io_A_Valid_1_delay_26_4 <= io_A_Valid_1_delay_25_5;
    io_A_Valid_1_delay_27_3 <= io_A_Valid_1_delay_26_4;
    io_A_Valid_1_delay_28_2 <= io_A_Valid_1_delay_27_3;
    io_A_Valid_1_delay_29_1 <= io_A_Valid_1_delay_28_2;
    io_A_Valid_1_delay_30 <= io_A_Valid_1_delay_29_1;
    io_B_Valid_30_delay_1 <= io_B_Valid_30;
    io_A_Valid_1_delay_1_30 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_29 <= io_A_Valid_1_delay_1_30;
    io_A_Valid_1_delay_3_28 <= io_A_Valid_1_delay_2_29;
    io_A_Valid_1_delay_4_27 <= io_A_Valid_1_delay_3_28;
    io_A_Valid_1_delay_5_26 <= io_A_Valid_1_delay_4_27;
    io_A_Valid_1_delay_6_25 <= io_A_Valid_1_delay_5_26;
    io_A_Valid_1_delay_7_24 <= io_A_Valid_1_delay_6_25;
    io_A_Valid_1_delay_8_23 <= io_A_Valid_1_delay_7_24;
    io_A_Valid_1_delay_9_22 <= io_A_Valid_1_delay_8_23;
    io_A_Valid_1_delay_10_21 <= io_A_Valid_1_delay_9_22;
    io_A_Valid_1_delay_11_20 <= io_A_Valid_1_delay_10_21;
    io_A_Valid_1_delay_12_19 <= io_A_Valid_1_delay_11_20;
    io_A_Valid_1_delay_13_18 <= io_A_Valid_1_delay_12_19;
    io_A_Valid_1_delay_14_17 <= io_A_Valid_1_delay_13_18;
    io_A_Valid_1_delay_15_16 <= io_A_Valid_1_delay_14_17;
    io_A_Valid_1_delay_16_15 <= io_A_Valid_1_delay_15_16;
    io_A_Valid_1_delay_17_14 <= io_A_Valid_1_delay_16_15;
    io_A_Valid_1_delay_18_13 <= io_A_Valid_1_delay_17_14;
    io_A_Valid_1_delay_19_12 <= io_A_Valid_1_delay_18_13;
    io_A_Valid_1_delay_20_11 <= io_A_Valid_1_delay_19_12;
    io_A_Valid_1_delay_21_10 <= io_A_Valid_1_delay_20_11;
    io_A_Valid_1_delay_22_9 <= io_A_Valid_1_delay_21_10;
    io_A_Valid_1_delay_23_8 <= io_A_Valid_1_delay_22_9;
    io_A_Valid_1_delay_24_7 <= io_A_Valid_1_delay_23_8;
    io_A_Valid_1_delay_25_6 <= io_A_Valid_1_delay_24_7;
    io_A_Valid_1_delay_26_5 <= io_A_Valid_1_delay_25_6;
    io_A_Valid_1_delay_27_4 <= io_A_Valid_1_delay_26_5;
    io_A_Valid_1_delay_28_3 <= io_A_Valid_1_delay_27_4;
    io_A_Valid_1_delay_29_2 <= io_A_Valid_1_delay_28_3;
    io_A_Valid_1_delay_30_1 <= io_A_Valid_1_delay_29_2;
    io_A_Valid_1_delay_31 <= io_A_Valid_1_delay_30_1;
    io_B_Valid_31_delay_1 <= io_B_Valid_31;
    io_A_Valid_1_delay_1_31 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_30 <= io_A_Valid_1_delay_1_31;
    io_A_Valid_1_delay_3_29 <= io_A_Valid_1_delay_2_30;
    io_A_Valid_1_delay_4_28 <= io_A_Valid_1_delay_3_29;
    io_A_Valid_1_delay_5_27 <= io_A_Valid_1_delay_4_28;
    io_A_Valid_1_delay_6_26 <= io_A_Valid_1_delay_5_27;
    io_A_Valid_1_delay_7_25 <= io_A_Valid_1_delay_6_26;
    io_A_Valid_1_delay_8_24 <= io_A_Valid_1_delay_7_25;
    io_A_Valid_1_delay_9_23 <= io_A_Valid_1_delay_8_24;
    io_A_Valid_1_delay_10_22 <= io_A_Valid_1_delay_9_23;
    io_A_Valid_1_delay_11_21 <= io_A_Valid_1_delay_10_22;
    io_A_Valid_1_delay_12_20 <= io_A_Valid_1_delay_11_21;
    io_A_Valid_1_delay_13_19 <= io_A_Valid_1_delay_12_20;
    io_A_Valid_1_delay_14_18 <= io_A_Valid_1_delay_13_19;
    io_A_Valid_1_delay_15_17 <= io_A_Valid_1_delay_14_18;
    io_A_Valid_1_delay_16_16 <= io_A_Valid_1_delay_15_17;
    io_A_Valid_1_delay_17_15 <= io_A_Valid_1_delay_16_16;
    io_A_Valid_1_delay_18_14 <= io_A_Valid_1_delay_17_15;
    io_A_Valid_1_delay_19_13 <= io_A_Valid_1_delay_18_14;
    io_A_Valid_1_delay_20_12 <= io_A_Valid_1_delay_19_13;
    io_A_Valid_1_delay_21_11 <= io_A_Valid_1_delay_20_12;
    io_A_Valid_1_delay_22_10 <= io_A_Valid_1_delay_21_11;
    io_A_Valid_1_delay_23_9 <= io_A_Valid_1_delay_22_10;
    io_A_Valid_1_delay_24_8 <= io_A_Valid_1_delay_23_9;
    io_A_Valid_1_delay_25_7 <= io_A_Valid_1_delay_24_8;
    io_A_Valid_1_delay_26_6 <= io_A_Valid_1_delay_25_7;
    io_A_Valid_1_delay_27_5 <= io_A_Valid_1_delay_26_6;
    io_A_Valid_1_delay_28_4 <= io_A_Valid_1_delay_27_5;
    io_A_Valid_1_delay_29_3 <= io_A_Valid_1_delay_28_4;
    io_A_Valid_1_delay_30_2 <= io_A_Valid_1_delay_29_3;
    io_A_Valid_1_delay_31_1 <= io_A_Valid_1_delay_30_2;
    io_A_Valid_1_delay_32 <= io_A_Valid_1_delay_31_1;
    io_B_Valid_32_delay_1 <= io_B_Valid_32;
    io_A_Valid_1_delay_1_32 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_31 <= io_A_Valid_1_delay_1_32;
    io_A_Valid_1_delay_3_30 <= io_A_Valid_1_delay_2_31;
    io_A_Valid_1_delay_4_29 <= io_A_Valid_1_delay_3_30;
    io_A_Valid_1_delay_5_28 <= io_A_Valid_1_delay_4_29;
    io_A_Valid_1_delay_6_27 <= io_A_Valid_1_delay_5_28;
    io_A_Valid_1_delay_7_26 <= io_A_Valid_1_delay_6_27;
    io_A_Valid_1_delay_8_25 <= io_A_Valid_1_delay_7_26;
    io_A_Valid_1_delay_9_24 <= io_A_Valid_1_delay_8_25;
    io_A_Valid_1_delay_10_23 <= io_A_Valid_1_delay_9_24;
    io_A_Valid_1_delay_11_22 <= io_A_Valid_1_delay_10_23;
    io_A_Valid_1_delay_12_21 <= io_A_Valid_1_delay_11_22;
    io_A_Valid_1_delay_13_20 <= io_A_Valid_1_delay_12_21;
    io_A_Valid_1_delay_14_19 <= io_A_Valid_1_delay_13_20;
    io_A_Valid_1_delay_15_18 <= io_A_Valid_1_delay_14_19;
    io_A_Valid_1_delay_16_17 <= io_A_Valid_1_delay_15_18;
    io_A_Valid_1_delay_17_16 <= io_A_Valid_1_delay_16_17;
    io_A_Valid_1_delay_18_15 <= io_A_Valid_1_delay_17_16;
    io_A_Valid_1_delay_19_14 <= io_A_Valid_1_delay_18_15;
    io_A_Valid_1_delay_20_13 <= io_A_Valid_1_delay_19_14;
    io_A_Valid_1_delay_21_12 <= io_A_Valid_1_delay_20_13;
    io_A_Valid_1_delay_22_11 <= io_A_Valid_1_delay_21_12;
    io_A_Valid_1_delay_23_10 <= io_A_Valid_1_delay_22_11;
    io_A_Valid_1_delay_24_9 <= io_A_Valid_1_delay_23_10;
    io_A_Valid_1_delay_25_8 <= io_A_Valid_1_delay_24_9;
    io_A_Valid_1_delay_26_7 <= io_A_Valid_1_delay_25_8;
    io_A_Valid_1_delay_27_6 <= io_A_Valid_1_delay_26_7;
    io_A_Valid_1_delay_28_5 <= io_A_Valid_1_delay_27_6;
    io_A_Valid_1_delay_29_4 <= io_A_Valid_1_delay_28_5;
    io_A_Valid_1_delay_30_3 <= io_A_Valid_1_delay_29_4;
    io_A_Valid_1_delay_31_2 <= io_A_Valid_1_delay_30_3;
    io_A_Valid_1_delay_32_1 <= io_A_Valid_1_delay_31_2;
    io_A_Valid_1_delay_33 <= io_A_Valid_1_delay_32_1;
    io_B_Valid_33_delay_1 <= io_B_Valid_33;
    io_A_Valid_1_delay_1_33 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_32 <= io_A_Valid_1_delay_1_33;
    io_A_Valid_1_delay_3_31 <= io_A_Valid_1_delay_2_32;
    io_A_Valid_1_delay_4_30 <= io_A_Valid_1_delay_3_31;
    io_A_Valid_1_delay_5_29 <= io_A_Valid_1_delay_4_30;
    io_A_Valid_1_delay_6_28 <= io_A_Valid_1_delay_5_29;
    io_A_Valid_1_delay_7_27 <= io_A_Valid_1_delay_6_28;
    io_A_Valid_1_delay_8_26 <= io_A_Valid_1_delay_7_27;
    io_A_Valid_1_delay_9_25 <= io_A_Valid_1_delay_8_26;
    io_A_Valid_1_delay_10_24 <= io_A_Valid_1_delay_9_25;
    io_A_Valid_1_delay_11_23 <= io_A_Valid_1_delay_10_24;
    io_A_Valid_1_delay_12_22 <= io_A_Valid_1_delay_11_23;
    io_A_Valid_1_delay_13_21 <= io_A_Valid_1_delay_12_22;
    io_A_Valid_1_delay_14_20 <= io_A_Valid_1_delay_13_21;
    io_A_Valid_1_delay_15_19 <= io_A_Valid_1_delay_14_20;
    io_A_Valid_1_delay_16_18 <= io_A_Valid_1_delay_15_19;
    io_A_Valid_1_delay_17_17 <= io_A_Valid_1_delay_16_18;
    io_A_Valid_1_delay_18_16 <= io_A_Valid_1_delay_17_17;
    io_A_Valid_1_delay_19_15 <= io_A_Valid_1_delay_18_16;
    io_A_Valid_1_delay_20_14 <= io_A_Valid_1_delay_19_15;
    io_A_Valid_1_delay_21_13 <= io_A_Valid_1_delay_20_14;
    io_A_Valid_1_delay_22_12 <= io_A_Valid_1_delay_21_13;
    io_A_Valid_1_delay_23_11 <= io_A_Valid_1_delay_22_12;
    io_A_Valid_1_delay_24_10 <= io_A_Valid_1_delay_23_11;
    io_A_Valid_1_delay_25_9 <= io_A_Valid_1_delay_24_10;
    io_A_Valid_1_delay_26_8 <= io_A_Valid_1_delay_25_9;
    io_A_Valid_1_delay_27_7 <= io_A_Valid_1_delay_26_8;
    io_A_Valid_1_delay_28_6 <= io_A_Valid_1_delay_27_7;
    io_A_Valid_1_delay_29_5 <= io_A_Valid_1_delay_28_6;
    io_A_Valid_1_delay_30_4 <= io_A_Valid_1_delay_29_5;
    io_A_Valid_1_delay_31_3 <= io_A_Valid_1_delay_30_4;
    io_A_Valid_1_delay_32_2 <= io_A_Valid_1_delay_31_3;
    io_A_Valid_1_delay_33_1 <= io_A_Valid_1_delay_32_2;
    io_A_Valid_1_delay_34 <= io_A_Valid_1_delay_33_1;
    io_B_Valid_34_delay_1 <= io_B_Valid_34;
    io_A_Valid_1_delay_1_34 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_33 <= io_A_Valid_1_delay_1_34;
    io_A_Valid_1_delay_3_32 <= io_A_Valid_1_delay_2_33;
    io_A_Valid_1_delay_4_31 <= io_A_Valid_1_delay_3_32;
    io_A_Valid_1_delay_5_30 <= io_A_Valid_1_delay_4_31;
    io_A_Valid_1_delay_6_29 <= io_A_Valid_1_delay_5_30;
    io_A_Valid_1_delay_7_28 <= io_A_Valid_1_delay_6_29;
    io_A_Valid_1_delay_8_27 <= io_A_Valid_1_delay_7_28;
    io_A_Valid_1_delay_9_26 <= io_A_Valid_1_delay_8_27;
    io_A_Valid_1_delay_10_25 <= io_A_Valid_1_delay_9_26;
    io_A_Valid_1_delay_11_24 <= io_A_Valid_1_delay_10_25;
    io_A_Valid_1_delay_12_23 <= io_A_Valid_1_delay_11_24;
    io_A_Valid_1_delay_13_22 <= io_A_Valid_1_delay_12_23;
    io_A_Valid_1_delay_14_21 <= io_A_Valid_1_delay_13_22;
    io_A_Valid_1_delay_15_20 <= io_A_Valid_1_delay_14_21;
    io_A_Valid_1_delay_16_19 <= io_A_Valid_1_delay_15_20;
    io_A_Valid_1_delay_17_18 <= io_A_Valid_1_delay_16_19;
    io_A_Valid_1_delay_18_17 <= io_A_Valid_1_delay_17_18;
    io_A_Valid_1_delay_19_16 <= io_A_Valid_1_delay_18_17;
    io_A_Valid_1_delay_20_15 <= io_A_Valid_1_delay_19_16;
    io_A_Valid_1_delay_21_14 <= io_A_Valid_1_delay_20_15;
    io_A_Valid_1_delay_22_13 <= io_A_Valid_1_delay_21_14;
    io_A_Valid_1_delay_23_12 <= io_A_Valid_1_delay_22_13;
    io_A_Valid_1_delay_24_11 <= io_A_Valid_1_delay_23_12;
    io_A_Valid_1_delay_25_10 <= io_A_Valid_1_delay_24_11;
    io_A_Valid_1_delay_26_9 <= io_A_Valid_1_delay_25_10;
    io_A_Valid_1_delay_27_8 <= io_A_Valid_1_delay_26_9;
    io_A_Valid_1_delay_28_7 <= io_A_Valid_1_delay_27_8;
    io_A_Valid_1_delay_29_6 <= io_A_Valid_1_delay_28_7;
    io_A_Valid_1_delay_30_5 <= io_A_Valid_1_delay_29_6;
    io_A_Valid_1_delay_31_4 <= io_A_Valid_1_delay_30_5;
    io_A_Valid_1_delay_32_3 <= io_A_Valid_1_delay_31_4;
    io_A_Valid_1_delay_33_2 <= io_A_Valid_1_delay_32_3;
    io_A_Valid_1_delay_34_1 <= io_A_Valid_1_delay_33_2;
    io_A_Valid_1_delay_35 <= io_A_Valid_1_delay_34_1;
    io_B_Valid_35_delay_1 <= io_B_Valid_35;
    io_A_Valid_1_delay_1_35 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_34 <= io_A_Valid_1_delay_1_35;
    io_A_Valid_1_delay_3_33 <= io_A_Valid_1_delay_2_34;
    io_A_Valid_1_delay_4_32 <= io_A_Valid_1_delay_3_33;
    io_A_Valid_1_delay_5_31 <= io_A_Valid_1_delay_4_32;
    io_A_Valid_1_delay_6_30 <= io_A_Valid_1_delay_5_31;
    io_A_Valid_1_delay_7_29 <= io_A_Valid_1_delay_6_30;
    io_A_Valid_1_delay_8_28 <= io_A_Valid_1_delay_7_29;
    io_A_Valid_1_delay_9_27 <= io_A_Valid_1_delay_8_28;
    io_A_Valid_1_delay_10_26 <= io_A_Valid_1_delay_9_27;
    io_A_Valid_1_delay_11_25 <= io_A_Valid_1_delay_10_26;
    io_A_Valid_1_delay_12_24 <= io_A_Valid_1_delay_11_25;
    io_A_Valid_1_delay_13_23 <= io_A_Valid_1_delay_12_24;
    io_A_Valid_1_delay_14_22 <= io_A_Valid_1_delay_13_23;
    io_A_Valid_1_delay_15_21 <= io_A_Valid_1_delay_14_22;
    io_A_Valid_1_delay_16_20 <= io_A_Valid_1_delay_15_21;
    io_A_Valid_1_delay_17_19 <= io_A_Valid_1_delay_16_20;
    io_A_Valid_1_delay_18_18 <= io_A_Valid_1_delay_17_19;
    io_A_Valid_1_delay_19_17 <= io_A_Valid_1_delay_18_18;
    io_A_Valid_1_delay_20_16 <= io_A_Valid_1_delay_19_17;
    io_A_Valid_1_delay_21_15 <= io_A_Valid_1_delay_20_16;
    io_A_Valid_1_delay_22_14 <= io_A_Valid_1_delay_21_15;
    io_A_Valid_1_delay_23_13 <= io_A_Valid_1_delay_22_14;
    io_A_Valid_1_delay_24_12 <= io_A_Valid_1_delay_23_13;
    io_A_Valid_1_delay_25_11 <= io_A_Valid_1_delay_24_12;
    io_A_Valid_1_delay_26_10 <= io_A_Valid_1_delay_25_11;
    io_A_Valid_1_delay_27_9 <= io_A_Valid_1_delay_26_10;
    io_A_Valid_1_delay_28_8 <= io_A_Valid_1_delay_27_9;
    io_A_Valid_1_delay_29_7 <= io_A_Valid_1_delay_28_8;
    io_A_Valid_1_delay_30_6 <= io_A_Valid_1_delay_29_7;
    io_A_Valid_1_delay_31_5 <= io_A_Valid_1_delay_30_6;
    io_A_Valid_1_delay_32_4 <= io_A_Valid_1_delay_31_5;
    io_A_Valid_1_delay_33_3 <= io_A_Valid_1_delay_32_4;
    io_A_Valid_1_delay_34_2 <= io_A_Valid_1_delay_33_3;
    io_A_Valid_1_delay_35_1 <= io_A_Valid_1_delay_34_2;
    io_A_Valid_1_delay_36 <= io_A_Valid_1_delay_35_1;
    io_B_Valid_36_delay_1 <= io_B_Valid_36;
    io_A_Valid_1_delay_1_36 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_35 <= io_A_Valid_1_delay_1_36;
    io_A_Valid_1_delay_3_34 <= io_A_Valid_1_delay_2_35;
    io_A_Valid_1_delay_4_33 <= io_A_Valid_1_delay_3_34;
    io_A_Valid_1_delay_5_32 <= io_A_Valid_1_delay_4_33;
    io_A_Valid_1_delay_6_31 <= io_A_Valid_1_delay_5_32;
    io_A_Valid_1_delay_7_30 <= io_A_Valid_1_delay_6_31;
    io_A_Valid_1_delay_8_29 <= io_A_Valid_1_delay_7_30;
    io_A_Valid_1_delay_9_28 <= io_A_Valid_1_delay_8_29;
    io_A_Valid_1_delay_10_27 <= io_A_Valid_1_delay_9_28;
    io_A_Valid_1_delay_11_26 <= io_A_Valid_1_delay_10_27;
    io_A_Valid_1_delay_12_25 <= io_A_Valid_1_delay_11_26;
    io_A_Valid_1_delay_13_24 <= io_A_Valid_1_delay_12_25;
    io_A_Valid_1_delay_14_23 <= io_A_Valid_1_delay_13_24;
    io_A_Valid_1_delay_15_22 <= io_A_Valid_1_delay_14_23;
    io_A_Valid_1_delay_16_21 <= io_A_Valid_1_delay_15_22;
    io_A_Valid_1_delay_17_20 <= io_A_Valid_1_delay_16_21;
    io_A_Valid_1_delay_18_19 <= io_A_Valid_1_delay_17_20;
    io_A_Valid_1_delay_19_18 <= io_A_Valid_1_delay_18_19;
    io_A_Valid_1_delay_20_17 <= io_A_Valid_1_delay_19_18;
    io_A_Valid_1_delay_21_16 <= io_A_Valid_1_delay_20_17;
    io_A_Valid_1_delay_22_15 <= io_A_Valid_1_delay_21_16;
    io_A_Valid_1_delay_23_14 <= io_A_Valid_1_delay_22_15;
    io_A_Valid_1_delay_24_13 <= io_A_Valid_1_delay_23_14;
    io_A_Valid_1_delay_25_12 <= io_A_Valid_1_delay_24_13;
    io_A_Valid_1_delay_26_11 <= io_A_Valid_1_delay_25_12;
    io_A_Valid_1_delay_27_10 <= io_A_Valid_1_delay_26_11;
    io_A_Valid_1_delay_28_9 <= io_A_Valid_1_delay_27_10;
    io_A_Valid_1_delay_29_8 <= io_A_Valid_1_delay_28_9;
    io_A_Valid_1_delay_30_7 <= io_A_Valid_1_delay_29_8;
    io_A_Valid_1_delay_31_6 <= io_A_Valid_1_delay_30_7;
    io_A_Valid_1_delay_32_5 <= io_A_Valid_1_delay_31_6;
    io_A_Valid_1_delay_33_4 <= io_A_Valid_1_delay_32_5;
    io_A_Valid_1_delay_34_3 <= io_A_Valid_1_delay_33_4;
    io_A_Valid_1_delay_35_2 <= io_A_Valid_1_delay_34_3;
    io_A_Valid_1_delay_36_1 <= io_A_Valid_1_delay_35_2;
    io_A_Valid_1_delay_37 <= io_A_Valid_1_delay_36_1;
    io_B_Valid_37_delay_1 <= io_B_Valid_37;
    io_A_Valid_1_delay_1_37 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_36 <= io_A_Valid_1_delay_1_37;
    io_A_Valid_1_delay_3_35 <= io_A_Valid_1_delay_2_36;
    io_A_Valid_1_delay_4_34 <= io_A_Valid_1_delay_3_35;
    io_A_Valid_1_delay_5_33 <= io_A_Valid_1_delay_4_34;
    io_A_Valid_1_delay_6_32 <= io_A_Valid_1_delay_5_33;
    io_A_Valid_1_delay_7_31 <= io_A_Valid_1_delay_6_32;
    io_A_Valid_1_delay_8_30 <= io_A_Valid_1_delay_7_31;
    io_A_Valid_1_delay_9_29 <= io_A_Valid_1_delay_8_30;
    io_A_Valid_1_delay_10_28 <= io_A_Valid_1_delay_9_29;
    io_A_Valid_1_delay_11_27 <= io_A_Valid_1_delay_10_28;
    io_A_Valid_1_delay_12_26 <= io_A_Valid_1_delay_11_27;
    io_A_Valid_1_delay_13_25 <= io_A_Valid_1_delay_12_26;
    io_A_Valid_1_delay_14_24 <= io_A_Valid_1_delay_13_25;
    io_A_Valid_1_delay_15_23 <= io_A_Valid_1_delay_14_24;
    io_A_Valid_1_delay_16_22 <= io_A_Valid_1_delay_15_23;
    io_A_Valid_1_delay_17_21 <= io_A_Valid_1_delay_16_22;
    io_A_Valid_1_delay_18_20 <= io_A_Valid_1_delay_17_21;
    io_A_Valid_1_delay_19_19 <= io_A_Valid_1_delay_18_20;
    io_A_Valid_1_delay_20_18 <= io_A_Valid_1_delay_19_19;
    io_A_Valid_1_delay_21_17 <= io_A_Valid_1_delay_20_18;
    io_A_Valid_1_delay_22_16 <= io_A_Valid_1_delay_21_17;
    io_A_Valid_1_delay_23_15 <= io_A_Valid_1_delay_22_16;
    io_A_Valid_1_delay_24_14 <= io_A_Valid_1_delay_23_15;
    io_A_Valid_1_delay_25_13 <= io_A_Valid_1_delay_24_14;
    io_A_Valid_1_delay_26_12 <= io_A_Valid_1_delay_25_13;
    io_A_Valid_1_delay_27_11 <= io_A_Valid_1_delay_26_12;
    io_A_Valid_1_delay_28_10 <= io_A_Valid_1_delay_27_11;
    io_A_Valid_1_delay_29_9 <= io_A_Valid_1_delay_28_10;
    io_A_Valid_1_delay_30_8 <= io_A_Valid_1_delay_29_9;
    io_A_Valid_1_delay_31_7 <= io_A_Valid_1_delay_30_8;
    io_A_Valid_1_delay_32_6 <= io_A_Valid_1_delay_31_7;
    io_A_Valid_1_delay_33_5 <= io_A_Valid_1_delay_32_6;
    io_A_Valid_1_delay_34_4 <= io_A_Valid_1_delay_33_5;
    io_A_Valid_1_delay_35_3 <= io_A_Valid_1_delay_34_4;
    io_A_Valid_1_delay_36_2 <= io_A_Valid_1_delay_35_3;
    io_A_Valid_1_delay_37_1 <= io_A_Valid_1_delay_36_2;
    io_A_Valid_1_delay_38 <= io_A_Valid_1_delay_37_1;
    io_B_Valid_38_delay_1 <= io_B_Valid_38;
    io_A_Valid_1_delay_1_38 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_37 <= io_A_Valid_1_delay_1_38;
    io_A_Valid_1_delay_3_36 <= io_A_Valid_1_delay_2_37;
    io_A_Valid_1_delay_4_35 <= io_A_Valid_1_delay_3_36;
    io_A_Valid_1_delay_5_34 <= io_A_Valid_1_delay_4_35;
    io_A_Valid_1_delay_6_33 <= io_A_Valid_1_delay_5_34;
    io_A_Valid_1_delay_7_32 <= io_A_Valid_1_delay_6_33;
    io_A_Valid_1_delay_8_31 <= io_A_Valid_1_delay_7_32;
    io_A_Valid_1_delay_9_30 <= io_A_Valid_1_delay_8_31;
    io_A_Valid_1_delay_10_29 <= io_A_Valid_1_delay_9_30;
    io_A_Valid_1_delay_11_28 <= io_A_Valid_1_delay_10_29;
    io_A_Valid_1_delay_12_27 <= io_A_Valid_1_delay_11_28;
    io_A_Valid_1_delay_13_26 <= io_A_Valid_1_delay_12_27;
    io_A_Valid_1_delay_14_25 <= io_A_Valid_1_delay_13_26;
    io_A_Valid_1_delay_15_24 <= io_A_Valid_1_delay_14_25;
    io_A_Valid_1_delay_16_23 <= io_A_Valid_1_delay_15_24;
    io_A_Valid_1_delay_17_22 <= io_A_Valid_1_delay_16_23;
    io_A_Valid_1_delay_18_21 <= io_A_Valid_1_delay_17_22;
    io_A_Valid_1_delay_19_20 <= io_A_Valid_1_delay_18_21;
    io_A_Valid_1_delay_20_19 <= io_A_Valid_1_delay_19_20;
    io_A_Valid_1_delay_21_18 <= io_A_Valid_1_delay_20_19;
    io_A_Valid_1_delay_22_17 <= io_A_Valid_1_delay_21_18;
    io_A_Valid_1_delay_23_16 <= io_A_Valid_1_delay_22_17;
    io_A_Valid_1_delay_24_15 <= io_A_Valid_1_delay_23_16;
    io_A_Valid_1_delay_25_14 <= io_A_Valid_1_delay_24_15;
    io_A_Valid_1_delay_26_13 <= io_A_Valid_1_delay_25_14;
    io_A_Valid_1_delay_27_12 <= io_A_Valid_1_delay_26_13;
    io_A_Valid_1_delay_28_11 <= io_A_Valid_1_delay_27_12;
    io_A_Valid_1_delay_29_10 <= io_A_Valid_1_delay_28_11;
    io_A_Valid_1_delay_30_9 <= io_A_Valid_1_delay_29_10;
    io_A_Valid_1_delay_31_8 <= io_A_Valid_1_delay_30_9;
    io_A_Valid_1_delay_32_7 <= io_A_Valid_1_delay_31_8;
    io_A_Valid_1_delay_33_6 <= io_A_Valid_1_delay_32_7;
    io_A_Valid_1_delay_34_5 <= io_A_Valid_1_delay_33_6;
    io_A_Valid_1_delay_35_4 <= io_A_Valid_1_delay_34_5;
    io_A_Valid_1_delay_36_3 <= io_A_Valid_1_delay_35_4;
    io_A_Valid_1_delay_37_2 <= io_A_Valid_1_delay_36_3;
    io_A_Valid_1_delay_38_1 <= io_A_Valid_1_delay_37_2;
    io_A_Valid_1_delay_39 <= io_A_Valid_1_delay_38_1;
    io_B_Valid_39_delay_1 <= io_B_Valid_39;
    io_A_Valid_1_delay_1_39 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_38 <= io_A_Valid_1_delay_1_39;
    io_A_Valid_1_delay_3_37 <= io_A_Valid_1_delay_2_38;
    io_A_Valid_1_delay_4_36 <= io_A_Valid_1_delay_3_37;
    io_A_Valid_1_delay_5_35 <= io_A_Valid_1_delay_4_36;
    io_A_Valid_1_delay_6_34 <= io_A_Valid_1_delay_5_35;
    io_A_Valid_1_delay_7_33 <= io_A_Valid_1_delay_6_34;
    io_A_Valid_1_delay_8_32 <= io_A_Valid_1_delay_7_33;
    io_A_Valid_1_delay_9_31 <= io_A_Valid_1_delay_8_32;
    io_A_Valid_1_delay_10_30 <= io_A_Valid_1_delay_9_31;
    io_A_Valid_1_delay_11_29 <= io_A_Valid_1_delay_10_30;
    io_A_Valid_1_delay_12_28 <= io_A_Valid_1_delay_11_29;
    io_A_Valid_1_delay_13_27 <= io_A_Valid_1_delay_12_28;
    io_A_Valid_1_delay_14_26 <= io_A_Valid_1_delay_13_27;
    io_A_Valid_1_delay_15_25 <= io_A_Valid_1_delay_14_26;
    io_A_Valid_1_delay_16_24 <= io_A_Valid_1_delay_15_25;
    io_A_Valid_1_delay_17_23 <= io_A_Valid_1_delay_16_24;
    io_A_Valid_1_delay_18_22 <= io_A_Valid_1_delay_17_23;
    io_A_Valid_1_delay_19_21 <= io_A_Valid_1_delay_18_22;
    io_A_Valid_1_delay_20_20 <= io_A_Valid_1_delay_19_21;
    io_A_Valid_1_delay_21_19 <= io_A_Valid_1_delay_20_20;
    io_A_Valid_1_delay_22_18 <= io_A_Valid_1_delay_21_19;
    io_A_Valid_1_delay_23_17 <= io_A_Valid_1_delay_22_18;
    io_A_Valid_1_delay_24_16 <= io_A_Valid_1_delay_23_17;
    io_A_Valid_1_delay_25_15 <= io_A_Valid_1_delay_24_16;
    io_A_Valid_1_delay_26_14 <= io_A_Valid_1_delay_25_15;
    io_A_Valid_1_delay_27_13 <= io_A_Valid_1_delay_26_14;
    io_A_Valid_1_delay_28_12 <= io_A_Valid_1_delay_27_13;
    io_A_Valid_1_delay_29_11 <= io_A_Valid_1_delay_28_12;
    io_A_Valid_1_delay_30_10 <= io_A_Valid_1_delay_29_11;
    io_A_Valid_1_delay_31_9 <= io_A_Valid_1_delay_30_10;
    io_A_Valid_1_delay_32_8 <= io_A_Valid_1_delay_31_9;
    io_A_Valid_1_delay_33_7 <= io_A_Valid_1_delay_32_8;
    io_A_Valid_1_delay_34_6 <= io_A_Valid_1_delay_33_7;
    io_A_Valid_1_delay_35_5 <= io_A_Valid_1_delay_34_6;
    io_A_Valid_1_delay_36_4 <= io_A_Valid_1_delay_35_5;
    io_A_Valid_1_delay_37_3 <= io_A_Valid_1_delay_36_4;
    io_A_Valid_1_delay_38_2 <= io_A_Valid_1_delay_37_3;
    io_A_Valid_1_delay_39_1 <= io_A_Valid_1_delay_38_2;
    io_A_Valid_1_delay_40 <= io_A_Valid_1_delay_39_1;
    io_B_Valid_40_delay_1 <= io_B_Valid_40;
    io_A_Valid_1_delay_1_40 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_39 <= io_A_Valid_1_delay_1_40;
    io_A_Valid_1_delay_3_38 <= io_A_Valid_1_delay_2_39;
    io_A_Valid_1_delay_4_37 <= io_A_Valid_1_delay_3_38;
    io_A_Valid_1_delay_5_36 <= io_A_Valid_1_delay_4_37;
    io_A_Valid_1_delay_6_35 <= io_A_Valid_1_delay_5_36;
    io_A_Valid_1_delay_7_34 <= io_A_Valid_1_delay_6_35;
    io_A_Valid_1_delay_8_33 <= io_A_Valid_1_delay_7_34;
    io_A_Valid_1_delay_9_32 <= io_A_Valid_1_delay_8_33;
    io_A_Valid_1_delay_10_31 <= io_A_Valid_1_delay_9_32;
    io_A_Valid_1_delay_11_30 <= io_A_Valid_1_delay_10_31;
    io_A_Valid_1_delay_12_29 <= io_A_Valid_1_delay_11_30;
    io_A_Valid_1_delay_13_28 <= io_A_Valid_1_delay_12_29;
    io_A_Valid_1_delay_14_27 <= io_A_Valid_1_delay_13_28;
    io_A_Valid_1_delay_15_26 <= io_A_Valid_1_delay_14_27;
    io_A_Valid_1_delay_16_25 <= io_A_Valid_1_delay_15_26;
    io_A_Valid_1_delay_17_24 <= io_A_Valid_1_delay_16_25;
    io_A_Valid_1_delay_18_23 <= io_A_Valid_1_delay_17_24;
    io_A_Valid_1_delay_19_22 <= io_A_Valid_1_delay_18_23;
    io_A_Valid_1_delay_20_21 <= io_A_Valid_1_delay_19_22;
    io_A_Valid_1_delay_21_20 <= io_A_Valid_1_delay_20_21;
    io_A_Valid_1_delay_22_19 <= io_A_Valid_1_delay_21_20;
    io_A_Valid_1_delay_23_18 <= io_A_Valid_1_delay_22_19;
    io_A_Valid_1_delay_24_17 <= io_A_Valid_1_delay_23_18;
    io_A_Valid_1_delay_25_16 <= io_A_Valid_1_delay_24_17;
    io_A_Valid_1_delay_26_15 <= io_A_Valid_1_delay_25_16;
    io_A_Valid_1_delay_27_14 <= io_A_Valid_1_delay_26_15;
    io_A_Valid_1_delay_28_13 <= io_A_Valid_1_delay_27_14;
    io_A_Valid_1_delay_29_12 <= io_A_Valid_1_delay_28_13;
    io_A_Valid_1_delay_30_11 <= io_A_Valid_1_delay_29_12;
    io_A_Valid_1_delay_31_10 <= io_A_Valid_1_delay_30_11;
    io_A_Valid_1_delay_32_9 <= io_A_Valid_1_delay_31_10;
    io_A_Valid_1_delay_33_8 <= io_A_Valid_1_delay_32_9;
    io_A_Valid_1_delay_34_7 <= io_A_Valid_1_delay_33_8;
    io_A_Valid_1_delay_35_6 <= io_A_Valid_1_delay_34_7;
    io_A_Valid_1_delay_36_5 <= io_A_Valid_1_delay_35_6;
    io_A_Valid_1_delay_37_4 <= io_A_Valid_1_delay_36_5;
    io_A_Valid_1_delay_38_3 <= io_A_Valid_1_delay_37_4;
    io_A_Valid_1_delay_39_2 <= io_A_Valid_1_delay_38_3;
    io_A_Valid_1_delay_40_1 <= io_A_Valid_1_delay_39_2;
    io_A_Valid_1_delay_41 <= io_A_Valid_1_delay_40_1;
    io_B_Valid_41_delay_1 <= io_B_Valid_41;
    io_A_Valid_1_delay_1_41 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_40 <= io_A_Valid_1_delay_1_41;
    io_A_Valid_1_delay_3_39 <= io_A_Valid_1_delay_2_40;
    io_A_Valid_1_delay_4_38 <= io_A_Valid_1_delay_3_39;
    io_A_Valid_1_delay_5_37 <= io_A_Valid_1_delay_4_38;
    io_A_Valid_1_delay_6_36 <= io_A_Valid_1_delay_5_37;
    io_A_Valid_1_delay_7_35 <= io_A_Valid_1_delay_6_36;
    io_A_Valid_1_delay_8_34 <= io_A_Valid_1_delay_7_35;
    io_A_Valid_1_delay_9_33 <= io_A_Valid_1_delay_8_34;
    io_A_Valid_1_delay_10_32 <= io_A_Valid_1_delay_9_33;
    io_A_Valid_1_delay_11_31 <= io_A_Valid_1_delay_10_32;
    io_A_Valid_1_delay_12_30 <= io_A_Valid_1_delay_11_31;
    io_A_Valid_1_delay_13_29 <= io_A_Valid_1_delay_12_30;
    io_A_Valid_1_delay_14_28 <= io_A_Valid_1_delay_13_29;
    io_A_Valid_1_delay_15_27 <= io_A_Valid_1_delay_14_28;
    io_A_Valid_1_delay_16_26 <= io_A_Valid_1_delay_15_27;
    io_A_Valid_1_delay_17_25 <= io_A_Valid_1_delay_16_26;
    io_A_Valid_1_delay_18_24 <= io_A_Valid_1_delay_17_25;
    io_A_Valid_1_delay_19_23 <= io_A_Valid_1_delay_18_24;
    io_A_Valid_1_delay_20_22 <= io_A_Valid_1_delay_19_23;
    io_A_Valid_1_delay_21_21 <= io_A_Valid_1_delay_20_22;
    io_A_Valid_1_delay_22_20 <= io_A_Valid_1_delay_21_21;
    io_A_Valid_1_delay_23_19 <= io_A_Valid_1_delay_22_20;
    io_A_Valid_1_delay_24_18 <= io_A_Valid_1_delay_23_19;
    io_A_Valid_1_delay_25_17 <= io_A_Valid_1_delay_24_18;
    io_A_Valid_1_delay_26_16 <= io_A_Valid_1_delay_25_17;
    io_A_Valid_1_delay_27_15 <= io_A_Valid_1_delay_26_16;
    io_A_Valid_1_delay_28_14 <= io_A_Valid_1_delay_27_15;
    io_A_Valid_1_delay_29_13 <= io_A_Valid_1_delay_28_14;
    io_A_Valid_1_delay_30_12 <= io_A_Valid_1_delay_29_13;
    io_A_Valid_1_delay_31_11 <= io_A_Valid_1_delay_30_12;
    io_A_Valid_1_delay_32_10 <= io_A_Valid_1_delay_31_11;
    io_A_Valid_1_delay_33_9 <= io_A_Valid_1_delay_32_10;
    io_A_Valid_1_delay_34_8 <= io_A_Valid_1_delay_33_9;
    io_A_Valid_1_delay_35_7 <= io_A_Valid_1_delay_34_8;
    io_A_Valid_1_delay_36_6 <= io_A_Valid_1_delay_35_7;
    io_A_Valid_1_delay_37_5 <= io_A_Valid_1_delay_36_6;
    io_A_Valid_1_delay_38_4 <= io_A_Valid_1_delay_37_5;
    io_A_Valid_1_delay_39_3 <= io_A_Valid_1_delay_38_4;
    io_A_Valid_1_delay_40_2 <= io_A_Valid_1_delay_39_3;
    io_A_Valid_1_delay_41_1 <= io_A_Valid_1_delay_40_2;
    io_A_Valid_1_delay_42 <= io_A_Valid_1_delay_41_1;
    io_B_Valid_42_delay_1 <= io_B_Valid_42;
    io_A_Valid_1_delay_1_42 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_41 <= io_A_Valid_1_delay_1_42;
    io_A_Valid_1_delay_3_40 <= io_A_Valid_1_delay_2_41;
    io_A_Valid_1_delay_4_39 <= io_A_Valid_1_delay_3_40;
    io_A_Valid_1_delay_5_38 <= io_A_Valid_1_delay_4_39;
    io_A_Valid_1_delay_6_37 <= io_A_Valid_1_delay_5_38;
    io_A_Valid_1_delay_7_36 <= io_A_Valid_1_delay_6_37;
    io_A_Valid_1_delay_8_35 <= io_A_Valid_1_delay_7_36;
    io_A_Valid_1_delay_9_34 <= io_A_Valid_1_delay_8_35;
    io_A_Valid_1_delay_10_33 <= io_A_Valid_1_delay_9_34;
    io_A_Valid_1_delay_11_32 <= io_A_Valid_1_delay_10_33;
    io_A_Valid_1_delay_12_31 <= io_A_Valid_1_delay_11_32;
    io_A_Valid_1_delay_13_30 <= io_A_Valid_1_delay_12_31;
    io_A_Valid_1_delay_14_29 <= io_A_Valid_1_delay_13_30;
    io_A_Valid_1_delay_15_28 <= io_A_Valid_1_delay_14_29;
    io_A_Valid_1_delay_16_27 <= io_A_Valid_1_delay_15_28;
    io_A_Valid_1_delay_17_26 <= io_A_Valid_1_delay_16_27;
    io_A_Valid_1_delay_18_25 <= io_A_Valid_1_delay_17_26;
    io_A_Valid_1_delay_19_24 <= io_A_Valid_1_delay_18_25;
    io_A_Valid_1_delay_20_23 <= io_A_Valid_1_delay_19_24;
    io_A_Valid_1_delay_21_22 <= io_A_Valid_1_delay_20_23;
    io_A_Valid_1_delay_22_21 <= io_A_Valid_1_delay_21_22;
    io_A_Valid_1_delay_23_20 <= io_A_Valid_1_delay_22_21;
    io_A_Valid_1_delay_24_19 <= io_A_Valid_1_delay_23_20;
    io_A_Valid_1_delay_25_18 <= io_A_Valid_1_delay_24_19;
    io_A_Valid_1_delay_26_17 <= io_A_Valid_1_delay_25_18;
    io_A_Valid_1_delay_27_16 <= io_A_Valid_1_delay_26_17;
    io_A_Valid_1_delay_28_15 <= io_A_Valid_1_delay_27_16;
    io_A_Valid_1_delay_29_14 <= io_A_Valid_1_delay_28_15;
    io_A_Valid_1_delay_30_13 <= io_A_Valid_1_delay_29_14;
    io_A_Valid_1_delay_31_12 <= io_A_Valid_1_delay_30_13;
    io_A_Valid_1_delay_32_11 <= io_A_Valid_1_delay_31_12;
    io_A_Valid_1_delay_33_10 <= io_A_Valid_1_delay_32_11;
    io_A_Valid_1_delay_34_9 <= io_A_Valid_1_delay_33_10;
    io_A_Valid_1_delay_35_8 <= io_A_Valid_1_delay_34_9;
    io_A_Valid_1_delay_36_7 <= io_A_Valid_1_delay_35_8;
    io_A_Valid_1_delay_37_6 <= io_A_Valid_1_delay_36_7;
    io_A_Valid_1_delay_38_5 <= io_A_Valid_1_delay_37_6;
    io_A_Valid_1_delay_39_4 <= io_A_Valid_1_delay_38_5;
    io_A_Valid_1_delay_40_3 <= io_A_Valid_1_delay_39_4;
    io_A_Valid_1_delay_41_2 <= io_A_Valid_1_delay_40_3;
    io_A_Valid_1_delay_42_1 <= io_A_Valid_1_delay_41_2;
    io_A_Valid_1_delay_43 <= io_A_Valid_1_delay_42_1;
    io_B_Valid_43_delay_1 <= io_B_Valid_43;
    io_A_Valid_1_delay_1_43 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_42 <= io_A_Valid_1_delay_1_43;
    io_A_Valid_1_delay_3_41 <= io_A_Valid_1_delay_2_42;
    io_A_Valid_1_delay_4_40 <= io_A_Valid_1_delay_3_41;
    io_A_Valid_1_delay_5_39 <= io_A_Valid_1_delay_4_40;
    io_A_Valid_1_delay_6_38 <= io_A_Valid_1_delay_5_39;
    io_A_Valid_1_delay_7_37 <= io_A_Valid_1_delay_6_38;
    io_A_Valid_1_delay_8_36 <= io_A_Valid_1_delay_7_37;
    io_A_Valid_1_delay_9_35 <= io_A_Valid_1_delay_8_36;
    io_A_Valid_1_delay_10_34 <= io_A_Valid_1_delay_9_35;
    io_A_Valid_1_delay_11_33 <= io_A_Valid_1_delay_10_34;
    io_A_Valid_1_delay_12_32 <= io_A_Valid_1_delay_11_33;
    io_A_Valid_1_delay_13_31 <= io_A_Valid_1_delay_12_32;
    io_A_Valid_1_delay_14_30 <= io_A_Valid_1_delay_13_31;
    io_A_Valid_1_delay_15_29 <= io_A_Valid_1_delay_14_30;
    io_A_Valid_1_delay_16_28 <= io_A_Valid_1_delay_15_29;
    io_A_Valid_1_delay_17_27 <= io_A_Valid_1_delay_16_28;
    io_A_Valid_1_delay_18_26 <= io_A_Valid_1_delay_17_27;
    io_A_Valid_1_delay_19_25 <= io_A_Valid_1_delay_18_26;
    io_A_Valid_1_delay_20_24 <= io_A_Valid_1_delay_19_25;
    io_A_Valid_1_delay_21_23 <= io_A_Valid_1_delay_20_24;
    io_A_Valid_1_delay_22_22 <= io_A_Valid_1_delay_21_23;
    io_A_Valid_1_delay_23_21 <= io_A_Valid_1_delay_22_22;
    io_A_Valid_1_delay_24_20 <= io_A_Valid_1_delay_23_21;
    io_A_Valid_1_delay_25_19 <= io_A_Valid_1_delay_24_20;
    io_A_Valid_1_delay_26_18 <= io_A_Valid_1_delay_25_19;
    io_A_Valid_1_delay_27_17 <= io_A_Valid_1_delay_26_18;
    io_A_Valid_1_delay_28_16 <= io_A_Valid_1_delay_27_17;
    io_A_Valid_1_delay_29_15 <= io_A_Valid_1_delay_28_16;
    io_A_Valid_1_delay_30_14 <= io_A_Valid_1_delay_29_15;
    io_A_Valid_1_delay_31_13 <= io_A_Valid_1_delay_30_14;
    io_A_Valid_1_delay_32_12 <= io_A_Valid_1_delay_31_13;
    io_A_Valid_1_delay_33_11 <= io_A_Valid_1_delay_32_12;
    io_A_Valid_1_delay_34_10 <= io_A_Valid_1_delay_33_11;
    io_A_Valid_1_delay_35_9 <= io_A_Valid_1_delay_34_10;
    io_A_Valid_1_delay_36_8 <= io_A_Valid_1_delay_35_9;
    io_A_Valid_1_delay_37_7 <= io_A_Valid_1_delay_36_8;
    io_A_Valid_1_delay_38_6 <= io_A_Valid_1_delay_37_7;
    io_A_Valid_1_delay_39_5 <= io_A_Valid_1_delay_38_6;
    io_A_Valid_1_delay_40_4 <= io_A_Valid_1_delay_39_5;
    io_A_Valid_1_delay_41_3 <= io_A_Valid_1_delay_40_4;
    io_A_Valid_1_delay_42_2 <= io_A_Valid_1_delay_41_3;
    io_A_Valid_1_delay_43_1 <= io_A_Valid_1_delay_42_2;
    io_A_Valid_1_delay_44 <= io_A_Valid_1_delay_43_1;
    io_B_Valid_44_delay_1 <= io_B_Valid_44;
    io_A_Valid_1_delay_1_44 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_43 <= io_A_Valid_1_delay_1_44;
    io_A_Valid_1_delay_3_42 <= io_A_Valid_1_delay_2_43;
    io_A_Valid_1_delay_4_41 <= io_A_Valid_1_delay_3_42;
    io_A_Valid_1_delay_5_40 <= io_A_Valid_1_delay_4_41;
    io_A_Valid_1_delay_6_39 <= io_A_Valid_1_delay_5_40;
    io_A_Valid_1_delay_7_38 <= io_A_Valid_1_delay_6_39;
    io_A_Valid_1_delay_8_37 <= io_A_Valid_1_delay_7_38;
    io_A_Valid_1_delay_9_36 <= io_A_Valid_1_delay_8_37;
    io_A_Valid_1_delay_10_35 <= io_A_Valid_1_delay_9_36;
    io_A_Valid_1_delay_11_34 <= io_A_Valid_1_delay_10_35;
    io_A_Valid_1_delay_12_33 <= io_A_Valid_1_delay_11_34;
    io_A_Valid_1_delay_13_32 <= io_A_Valid_1_delay_12_33;
    io_A_Valid_1_delay_14_31 <= io_A_Valid_1_delay_13_32;
    io_A_Valid_1_delay_15_30 <= io_A_Valid_1_delay_14_31;
    io_A_Valid_1_delay_16_29 <= io_A_Valid_1_delay_15_30;
    io_A_Valid_1_delay_17_28 <= io_A_Valid_1_delay_16_29;
    io_A_Valid_1_delay_18_27 <= io_A_Valid_1_delay_17_28;
    io_A_Valid_1_delay_19_26 <= io_A_Valid_1_delay_18_27;
    io_A_Valid_1_delay_20_25 <= io_A_Valid_1_delay_19_26;
    io_A_Valid_1_delay_21_24 <= io_A_Valid_1_delay_20_25;
    io_A_Valid_1_delay_22_23 <= io_A_Valid_1_delay_21_24;
    io_A_Valid_1_delay_23_22 <= io_A_Valid_1_delay_22_23;
    io_A_Valid_1_delay_24_21 <= io_A_Valid_1_delay_23_22;
    io_A_Valid_1_delay_25_20 <= io_A_Valid_1_delay_24_21;
    io_A_Valid_1_delay_26_19 <= io_A_Valid_1_delay_25_20;
    io_A_Valid_1_delay_27_18 <= io_A_Valid_1_delay_26_19;
    io_A_Valid_1_delay_28_17 <= io_A_Valid_1_delay_27_18;
    io_A_Valid_1_delay_29_16 <= io_A_Valid_1_delay_28_17;
    io_A_Valid_1_delay_30_15 <= io_A_Valid_1_delay_29_16;
    io_A_Valid_1_delay_31_14 <= io_A_Valid_1_delay_30_15;
    io_A_Valid_1_delay_32_13 <= io_A_Valid_1_delay_31_14;
    io_A_Valid_1_delay_33_12 <= io_A_Valid_1_delay_32_13;
    io_A_Valid_1_delay_34_11 <= io_A_Valid_1_delay_33_12;
    io_A_Valid_1_delay_35_10 <= io_A_Valid_1_delay_34_11;
    io_A_Valid_1_delay_36_9 <= io_A_Valid_1_delay_35_10;
    io_A_Valid_1_delay_37_8 <= io_A_Valid_1_delay_36_9;
    io_A_Valid_1_delay_38_7 <= io_A_Valid_1_delay_37_8;
    io_A_Valid_1_delay_39_6 <= io_A_Valid_1_delay_38_7;
    io_A_Valid_1_delay_40_5 <= io_A_Valid_1_delay_39_6;
    io_A_Valid_1_delay_41_4 <= io_A_Valid_1_delay_40_5;
    io_A_Valid_1_delay_42_3 <= io_A_Valid_1_delay_41_4;
    io_A_Valid_1_delay_43_2 <= io_A_Valid_1_delay_42_3;
    io_A_Valid_1_delay_44_1 <= io_A_Valid_1_delay_43_2;
    io_A_Valid_1_delay_45 <= io_A_Valid_1_delay_44_1;
    io_B_Valid_45_delay_1 <= io_B_Valid_45;
    io_A_Valid_1_delay_1_45 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_44 <= io_A_Valid_1_delay_1_45;
    io_A_Valid_1_delay_3_43 <= io_A_Valid_1_delay_2_44;
    io_A_Valid_1_delay_4_42 <= io_A_Valid_1_delay_3_43;
    io_A_Valid_1_delay_5_41 <= io_A_Valid_1_delay_4_42;
    io_A_Valid_1_delay_6_40 <= io_A_Valid_1_delay_5_41;
    io_A_Valid_1_delay_7_39 <= io_A_Valid_1_delay_6_40;
    io_A_Valid_1_delay_8_38 <= io_A_Valid_1_delay_7_39;
    io_A_Valid_1_delay_9_37 <= io_A_Valid_1_delay_8_38;
    io_A_Valid_1_delay_10_36 <= io_A_Valid_1_delay_9_37;
    io_A_Valid_1_delay_11_35 <= io_A_Valid_1_delay_10_36;
    io_A_Valid_1_delay_12_34 <= io_A_Valid_1_delay_11_35;
    io_A_Valid_1_delay_13_33 <= io_A_Valid_1_delay_12_34;
    io_A_Valid_1_delay_14_32 <= io_A_Valid_1_delay_13_33;
    io_A_Valid_1_delay_15_31 <= io_A_Valid_1_delay_14_32;
    io_A_Valid_1_delay_16_30 <= io_A_Valid_1_delay_15_31;
    io_A_Valid_1_delay_17_29 <= io_A_Valid_1_delay_16_30;
    io_A_Valid_1_delay_18_28 <= io_A_Valid_1_delay_17_29;
    io_A_Valid_1_delay_19_27 <= io_A_Valid_1_delay_18_28;
    io_A_Valid_1_delay_20_26 <= io_A_Valid_1_delay_19_27;
    io_A_Valid_1_delay_21_25 <= io_A_Valid_1_delay_20_26;
    io_A_Valid_1_delay_22_24 <= io_A_Valid_1_delay_21_25;
    io_A_Valid_1_delay_23_23 <= io_A_Valid_1_delay_22_24;
    io_A_Valid_1_delay_24_22 <= io_A_Valid_1_delay_23_23;
    io_A_Valid_1_delay_25_21 <= io_A_Valid_1_delay_24_22;
    io_A_Valid_1_delay_26_20 <= io_A_Valid_1_delay_25_21;
    io_A_Valid_1_delay_27_19 <= io_A_Valid_1_delay_26_20;
    io_A_Valid_1_delay_28_18 <= io_A_Valid_1_delay_27_19;
    io_A_Valid_1_delay_29_17 <= io_A_Valid_1_delay_28_18;
    io_A_Valid_1_delay_30_16 <= io_A_Valid_1_delay_29_17;
    io_A_Valid_1_delay_31_15 <= io_A_Valid_1_delay_30_16;
    io_A_Valid_1_delay_32_14 <= io_A_Valid_1_delay_31_15;
    io_A_Valid_1_delay_33_13 <= io_A_Valid_1_delay_32_14;
    io_A_Valid_1_delay_34_12 <= io_A_Valid_1_delay_33_13;
    io_A_Valid_1_delay_35_11 <= io_A_Valid_1_delay_34_12;
    io_A_Valid_1_delay_36_10 <= io_A_Valid_1_delay_35_11;
    io_A_Valid_1_delay_37_9 <= io_A_Valid_1_delay_36_10;
    io_A_Valid_1_delay_38_8 <= io_A_Valid_1_delay_37_9;
    io_A_Valid_1_delay_39_7 <= io_A_Valid_1_delay_38_8;
    io_A_Valid_1_delay_40_6 <= io_A_Valid_1_delay_39_7;
    io_A_Valid_1_delay_41_5 <= io_A_Valid_1_delay_40_6;
    io_A_Valid_1_delay_42_4 <= io_A_Valid_1_delay_41_5;
    io_A_Valid_1_delay_43_3 <= io_A_Valid_1_delay_42_4;
    io_A_Valid_1_delay_44_2 <= io_A_Valid_1_delay_43_3;
    io_A_Valid_1_delay_45_1 <= io_A_Valid_1_delay_44_2;
    io_A_Valid_1_delay_46 <= io_A_Valid_1_delay_45_1;
    io_B_Valid_46_delay_1 <= io_B_Valid_46;
    io_A_Valid_1_delay_1_46 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_45 <= io_A_Valid_1_delay_1_46;
    io_A_Valid_1_delay_3_44 <= io_A_Valid_1_delay_2_45;
    io_A_Valid_1_delay_4_43 <= io_A_Valid_1_delay_3_44;
    io_A_Valid_1_delay_5_42 <= io_A_Valid_1_delay_4_43;
    io_A_Valid_1_delay_6_41 <= io_A_Valid_1_delay_5_42;
    io_A_Valid_1_delay_7_40 <= io_A_Valid_1_delay_6_41;
    io_A_Valid_1_delay_8_39 <= io_A_Valid_1_delay_7_40;
    io_A_Valid_1_delay_9_38 <= io_A_Valid_1_delay_8_39;
    io_A_Valid_1_delay_10_37 <= io_A_Valid_1_delay_9_38;
    io_A_Valid_1_delay_11_36 <= io_A_Valid_1_delay_10_37;
    io_A_Valid_1_delay_12_35 <= io_A_Valid_1_delay_11_36;
    io_A_Valid_1_delay_13_34 <= io_A_Valid_1_delay_12_35;
    io_A_Valid_1_delay_14_33 <= io_A_Valid_1_delay_13_34;
    io_A_Valid_1_delay_15_32 <= io_A_Valid_1_delay_14_33;
    io_A_Valid_1_delay_16_31 <= io_A_Valid_1_delay_15_32;
    io_A_Valid_1_delay_17_30 <= io_A_Valid_1_delay_16_31;
    io_A_Valid_1_delay_18_29 <= io_A_Valid_1_delay_17_30;
    io_A_Valid_1_delay_19_28 <= io_A_Valid_1_delay_18_29;
    io_A_Valid_1_delay_20_27 <= io_A_Valid_1_delay_19_28;
    io_A_Valid_1_delay_21_26 <= io_A_Valid_1_delay_20_27;
    io_A_Valid_1_delay_22_25 <= io_A_Valid_1_delay_21_26;
    io_A_Valid_1_delay_23_24 <= io_A_Valid_1_delay_22_25;
    io_A_Valid_1_delay_24_23 <= io_A_Valid_1_delay_23_24;
    io_A_Valid_1_delay_25_22 <= io_A_Valid_1_delay_24_23;
    io_A_Valid_1_delay_26_21 <= io_A_Valid_1_delay_25_22;
    io_A_Valid_1_delay_27_20 <= io_A_Valid_1_delay_26_21;
    io_A_Valid_1_delay_28_19 <= io_A_Valid_1_delay_27_20;
    io_A_Valid_1_delay_29_18 <= io_A_Valid_1_delay_28_19;
    io_A_Valid_1_delay_30_17 <= io_A_Valid_1_delay_29_18;
    io_A_Valid_1_delay_31_16 <= io_A_Valid_1_delay_30_17;
    io_A_Valid_1_delay_32_15 <= io_A_Valid_1_delay_31_16;
    io_A_Valid_1_delay_33_14 <= io_A_Valid_1_delay_32_15;
    io_A_Valid_1_delay_34_13 <= io_A_Valid_1_delay_33_14;
    io_A_Valid_1_delay_35_12 <= io_A_Valid_1_delay_34_13;
    io_A_Valid_1_delay_36_11 <= io_A_Valid_1_delay_35_12;
    io_A_Valid_1_delay_37_10 <= io_A_Valid_1_delay_36_11;
    io_A_Valid_1_delay_38_9 <= io_A_Valid_1_delay_37_10;
    io_A_Valid_1_delay_39_8 <= io_A_Valid_1_delay_38_9;
    io_A_Valid_1_delay_40_7 <= io_A_Valid_1_delay_39_8;
    io_A_Valid_1_delay_41_6 <= io_A_Valid_1_delay_40_7;
    io_A_Valid_1_delay_42_5 <= io_A_Valid_1_delay_41_6;
    io_A_Valid_1_delay_43_4 <= io_A_Valid_1_delay_42_5;
    io_A_Valid_1_delay_44_3 <= io_A_Valid_1_delay_43_4;
    io_A_Valid_1_delay_45_2 <= io_A_Valid_1_delay_44_3;
    io_A_Valid_1_delay_46_1 <= io_A_Valid_1_delay_45_2;
    io_A_Valid_1_delay_47 <= io_A_Valid_1_delay_46_1;
    io_B_Valid_47_delay_1 <= io_B_Valid_47;
    io_A_Valid_1_delay_1_47 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_46 <= io_A_Valid_1_delay_1_47;
    io_A_Valid_1_delay_3_45 <= io_A_Valid_1_delay_2_46;
    io_A_Valid_1_delay_4_44 <= io_A_Valid_1_delay_3_45;
    io_A_Valid_1_delay_5_43 <= io_A_Valid_1_delay_4_44;
    io_A_Valid_1_delay_6_42 <= io_A_Valid_1_delay_5_43;
    io_A_Valid_1_delay_7_41 <= io_A_Valid_1_delay_6_42;
    io_A_Valid_1_delay_8_40 <= io_A_Valid_1_delay_7_41;
    io_A_Valid_1_delay_9_39 <= io_A_Valid_1_delay_8_40;
    io_A_Valid_1_delay_10_38 <= io_A_Valid_1_delay_9_39;
    io_A_Valid_1_delay_11_37 <= io_A_Valid_1_delay_10_38;
    io_A_Valid_1_delay_12_36 <= io_A_Valid_1_delay_11_37;
    io_A_Valid_1_delay_13_35 <= io_A_Valid_1_delay_12_36;
    io_A_Valid_1_delay_14_34 <= io_A_Valid_1_delay_13_35;
    io_A_Valid_1_delay_15_33 <= io_A_Valid_1_delay_14_34;
    io_A_Valid_1_delay_16_32 <= io_A_Valid_1_delay_15_33;
    io_A_Valid_1_delay_17_31 <= io_A_Valid_1_delay_16_32;
    io_A_Valid_1_delay_18_30 <= io_A_Valid_1_delay_17_31;
    io_A_Valid_1_delay_19_29 <= io_A_Valid_1_delay_18_30;
    io_A_Valid_1_delay_20_28 <= io_A_Valid_1_delay_19_29;
    io_A_Valid_1_delay_21_27 <= io_A_Valid_1_delay_20_28;
    io_A_Valid_1_delay_22_26 <= io_A_Valid_1_delay_21_27;
    io_A_Valid_1_delay_23_25 <= io_A_Valid_1_delay_22_26;
    io_A_Valid_1_delay_24_24 <= io_A_Valid_1_delay_23_25;
    io_A_Valid_1_delay_25_23 <= io_A_Valid_1_delay_24_24;
    io_A_Valid_1_delay_26_22 <= io_A_Valid_1_delay_25_23;
    io_A_Valid_1_delay_27_21 <= io_A_Valid_1_delay_26_22;
    io_A_Valid_1_delay_28_20 <= io_A_Valid_1_delay_27_21;
    io_A_Valid_1_delay_29_19 <= io_A_Valid_1_delay_28_20;
    io_A_Valid_1_delay_30_18 <= io_A_Valid_1_delay_29_19;
    io_A_Valid_1_delay_31_17 <= io_A_Valid_1_delay_30_18;
    io_A_Valid_1_delay_32_16 <= io_A_Valid_1_delay_31_17;
    io_A_Valid_1_delay_33_15 <= io_A_Valid_1_delay_32_16;
    io_A_Valid_1_delay_34_14 <= io_A_Valid_1_delay_33_15;
    io_A_Valid_1_delay_35_13 <= io_A_Valid_1_delay_34_14;
    io_A_Valid_1_delay_36_12 <= io_A_Valid_1_delay_35_13;
    io_A_Valid_1_delay_37_11 <= io_A_Valid_1_delay_36_12;
    io_A_Valid_1_delay_38_10 <= io_A_Valid_1_delay_37_11;
    io_A_Valid_1_delay_39_9 <= io_A_Valid_1_delay_38_10;
    io_A_Valid_1_delay_40_8 <= io_A_Valid_1_delay_39_9;
    io_A_Valid_1_delay_41_7 <= io_A_Valid_1_delay_40_8;
    io_A_Valid_1_delay_42_6 <= io_A_Valid_1_delay_41_7;
    io_A_Valid_1_delay_43_5 <= io_A_Valid_1_delay_42_6;
    io_A_Valid_1_delay_44_4 <= io_A_Valid_1_delay_43_5;
    io_A_Valid_1_delay_45_3 <= io_A_Valid_1_delay_44_4;
    io_A_Valid_1_delay_46_2 <= io_A_Valid_1_delay_45_3;
    io_A_Valid_1_delay_47_1 <= io_A_Valid_1_delay_46_2;
    io_A_Valid_1_delay_48 <= io_A_Valid_1_delay_47_1;
    io_B_Valid_48_delay_1 <= io_B_Valid_48;
    io_A_Valid_1_delay_1_48 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_47 <= io_A_Valid_1_delay_1_48;
    io_A_Valid_1_delay_3_46 <= io_A_Valid_1_delay_2_47;
    io_A_Valid_1_delay_4_45 <= io_A_Valid_1_delay_3_46;
    io_A_Valid_1_delay_5_44 <= io_A_Valid_1_delay_4_45;
    io_A_Valid_1_delay_6_43 <= io_A_Valid_1_delay_5_44;
    io_A_Valid_1_delay_7_42 <= io_A_Valid_1_delay_6_43;
    io_A_Valid_1_delay_8_41 <= io_A_Valid_1_delay_7_42;
    io_A_Valid_1_delay_9_40 <= io_A_Valid_1_delay_8_41;
    io_A_Valid_1_delay_10_39 <= io_A_Valid_1_delay_9_40;
    io_A_Valid_1_delay_11_38 <= io_A_Valid_1_delay_10_39;
    io_A_Valid_1_delay_12_37 <= io_A_Valid_1_delay_11_38;
    io_A_Valid_1_delay_13_36 <= io_A_Valid_1_delay_12_37;
    io_A_Valid_1_delay_14_35 <= io_A_Valid_1_delay_13_36;
    io_A_Valid_1_delay_15_34 <= io_A_Valid_1_delay_14_35;
    io_A_Valid_1_delay_16_33 <= io_A_Valid_1_delay_15_34;
    io_A_Valid_1_delay_17_32 <= io_A_Valid_1_delay_16_33;
    io_A_Valid_1_delay_18_31 <= io_A_Valid_1_delay_17_32;
    io_A_Valid_1_delay_19_30 <= io_A_Valid_1_delay_18_31;
    io_A_Valid_1_delay_20_29 <= io_A_Valid_1_delay_19_30;
    io_A_Valid_1_delay_21_28 <= io_A_Valid_1_delay_20_29;
    io_A_Valid_1_delay_22_27 <= io_A_Valid_1_delay_21_28;
    io_A_Valid_1_delay_23_26 <= io_A_Valid_1_delay_22_27;
    io_A_Valid_1_delay_24_25 <= io_A_Valid_1_delay_23_26;
    io_A_Valid_1_delay_25_24 <= io_A_Valid_1_delay_24_25;
    io_A_Valid_1_delay_26_23 <= io_A_Valid_1_delay_25_24;
    io_A_Valid_1_delay_27_22 <= io_A_Valid_1_delay_26_23;
    io_A_Valid_1_delay_28_21 <= io_A_Valid_1_delay_27_22;
    io_A_Valid_1_delay_29_20 <= io_A_Valid_1_delay_28_21;
    io_A_Valid_1_delay_30_19 <= io_A_Valid_1_delay_29_20;
    io_A_Valid_1_delay_31_18 <= io_A_Valid_1_delay_30_19;
    io_A_Valid_1_delay_32_17 <= io_A_Valid_1_delay_31_18;
    io_A_Valid_1_delay_33_16 <= io_A_Valid_1_delay_32_17;
    io_A_Valid_1_delay_34_15 <= io_A_Valid_1_delay_33_16;
    io_A_Valid_1_delay_35_14 <= io_A_Valid_1_delay_34_15;
    io_A_Valid_1_delay_36_13 <= io_A_Valid_1_delay_35_14;
    io_A_Valid_1_delay_37_12 <= io_A_Valid_1_delay_36_13;
    io_A_Valid_1_delay_38_11 <= io_A_Valid_1_delay_37_12;
    io_A_Valid_1_delay_39_10 <= io_A_Valid_1_delay_38_11;
    io_A_Valid_1_delay_40_9 <= io_A_Valid_1_delay_39_10;
    io_A_Valid_1_delay_41_8 <= io_A_Valid_1_delay_40_9;
    io_A_Valid_1_delay_42_7 <= io_A_Valid_1_delay_41_8;
    io_A_Valid_1_delay_43_6 <= io_A_Valid_1_delay_42_7;
    io_A_Valid_1_delay_44_5 <= io_A_Valid_1_delay_43_6;
    io_A_Valid_1_delay_45_4 <= io_A_Valid_1_delay_44_5;
    io_A_Valid_1_delay_46_3 <= io_A_Valid_1_delay_45_4;
    io_A_Valid_1_delay_47_2 <= io_A_Valid_1_delay_46_3;
    io_A_Valid_1_delay_48_1 <= io_A_Valid_1_delay_47_2;
    io_A_Valid_1_delay_49 <= io_A_Valid_1_delay_48_1;
    io_B_Valid_49_delay_1 <= io_B_Valid_49;
    io_A_Valid_1_delay_1_49 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_48 <= io_A_Valid_1_delay_1_49;
    io_A_Valid_1_delay_3_47 <= io_A_Valid_1_delay_2_48;
    io_A_Valid_1_delay_4_46 <= io_A_Valid_1_delay_3_47;
    io_A_Valid_1_delay_5_45 <= io_A_Valid_1_delay_4_46;
    io_A_Valid_1_delay_6_44 <= io_A_Valid_1_delay_5_45;
    io_A_Valid_1_delay_7_43 <= io_A_Valid_1_delay_6_44;
    io_A_Valid_1_delay_8_42 <= io_A_Valid_1_delay_7_43;
    io_A_Valid_1_delay_9_41 <= io_A_Valid_1_delay_8_42;
    io_A_Valid_1_delay_10_40 <= io_A_Valid_1_delay_9_41;
    io_A_Valid_1_delay_11_39 <= io_A_Valid_1_delay_10_40;
    io_A_Valid_1_delay_12_38 <= io_A_Valid_1_delay_11_39;
    io_A_Valid_1_delay_13_37 <= io_A_Valid_1_delay_12_38;
    io_A_Valid_1_delay_14_36 <= io_A_Valid_1_delay_13_37;
    io_A_Valid_1_delay_15_35 <= io_A_Valid_1_delay_14_36;
    io_A_Valid_1_delay_16_34 <= io_A_Valid_1_delay_15_35;
    io_A_Valid_1_delay_17_33 <= io_A_Valid_1_delay_16_34;
    io_A_Valid_1_delay_18_32 <= io_A_Valid_1_delay_17_33;
    io_A_Valid_1_delay_19_31 <= io_A_Valid_1_delay_18_32;
    io_A_Valid_1_delay_20_30 <= io_A_Valid_1_delay_19_31;
    io_A_Valid_1_delay_21_29 <= io_A_Valid_1_delay_20_30;
    io_A_Valid_1_delay_22_28 <= io_A_Valid_1_delay_21_29;
    io_A_Valid_1_delay_23_27 <= io_A_Valid_1_delay_22_28;
    io_A_Valid_1_delay_24_26 <= io_A_Valid_1_delay_23_27;
    io_A_Valid_1_delay_25_25 <= io_A_Valid_1_delay_24_26;
    io_A_Valid_1_delay_26_24 <= io_A_Valid_1_delay_25_25;
    io_A_Valid_1_delay_27_23 <= io_A_Valid_1_delay_26_24;
    io_A_Valid_1_delay_28_22 <= io_A_Valid_1_delay_27_23;
    io_A_Valid_1_delay_29_21 <= io_A_Valid_1_delay_28_22;
    io_A_Valid_1_delay_30_20 <= io_A_Valid_1_delay_29_21;
    io_A_Valid_1_delay_31_19 <= io_A_Valid_1_delay_30_20;
    io_A_Valid_1_delay_32_18 <= io_A_Valid_1_delay_31_19;
    io_A_Valid_1_delay_33_17 <= io_A_Valid_1_delay_32_18;
    io_A_Valid_1_delay_34_16 <= io_A_Valid_1_delay_33_17;
    io_A_Valid_1_delay_35_15 <= io_A_Valid_1_delay_34_16;
    io_A_Valid_1_delay_36_14 <= io_A_Valid_1_delay_35_15;
    io_A_Valid_1_delay_37_13 <= io_A_Valid_1_delay_36_14;
    io_A_Valid_1_delay_38_12 <= io_A_Valid_1_delay_37_13;
    io_A_Valid_1_delay_39_11 <= io_A_Valid_1_delay_38_12;
    io_A_Valid_1_delay_40_10 <= io_A_Valid_1_delay_39_11;
    io_A_Valid_1_delay_41_9 <= io_A_Valid_1_delay_40_10;
    io_A_Valid_1_delay_42_8 <= io_A_Valid_1_delay_41_9;
    io_A_Valid_1_delay_43_7 <= io_A_Valid_1_delay_42_8;
    io_A_Valid_1_delay_44_6 <= io_A_Valid_1_delay_43_7;
    io_A_Valid_1_delay_45_5 <= io_A_Valid_1_delay_44_6;
    io_A_Valid_1_delay_46_4 <= io_A_Valid_1_delay_45_5;
    io_A_Valid_1_delay_47_3 <= io_A_Valid_1_delay_46_4;
    io_A_Valid_1_delay_48_2 <= io_A_Valid_1_delay_47_3;
    io_A_Valid_1_delay_49_1 <= io_A_Valid_1_delay_48_2;
    io_A_Valid_1_delay_50 <= io_A_Valid_1_delay_49_1;
    io_B_Valid_50_delay_1 <= io_B_Valid_50;
    io_A_Valid_1_delay_1_50 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_49 <= io_A_Valid_1_delay_1_50;
    io_A_Valid_1_delay_3_48 <= io_A_Valid_1_delay_2_49;
    io_A_Valid_1_delay_4_47 <= io_A_Valid_1_delay_3_48;
    io_A_Valid_1_delay_5_46 <= io_A_Valid_1_delay_4_47;
    io_A_Valid_1_delay_6_45 <= io_A_Valid_1_delay_5_46;
    io_A_Valid_1_delay_7_44 <= io_A_Valid_1_delay_6_45;
    io_A_Valid_1_delay_8_43 <= io_A_Valid_1_delay_7_44;
    io_A_Valid_1_delay_9_42 <= io_A_Valid_1_delay_8_43;
    io_A_Valid_1_delay_10_41 <= io_A_Valid_1_delay_9_42;
    io_A_Valid_1_delay_11_40 <= io_A_Valid_1_delay_10_41;
    io_A_Valid_1_delay_12_39 <= io_A_Valid_1_delay_11_40;
    io_A_Valid_1_delay_13_38 <= io_A_Valid_1_delay_12_39;
    io_A_Valid_1_delay_14_37 <= io_A_Valid_1_delay_13_38;
    io_A_Valid_1_delay_15_36 <= io_A_Valid_1_delay_14_37;
    io_A_Valid_1_delay_16_35 <= io_A_Valid_1_delay_15_36;
    io_A_Valid_1_delay_17_34 <= io_A_Valid_1_delay_16_35;
    io_A_Valid_1_delay_18_33 <= io_A_Valid_1_delay_17_34;
    io_A_Valid_1_delay_19_32 <= io_A_Valid_1_delay_18_33;
    io_A_Valid_1_delay_20_31 <= io_A_Valid_1_delay_19_32;
    io_A_Valid_1_delay_21_30 <= io_A_Valid_1_delay_20_31;
    io_A_Valid_1_delay_22_29 <= io_A_Valid_1_delay_21_30;
    io_A_Valid_1_delay_23_28 <= io_A_Valid_1_delay_22_29;
    io_A_Valid_1_delay_24_27 <= io_A_Valid_1_delay_23_28;
    io_A_Valid_1_delay_25_26 <= io_A_Valid_1_delay_24_27;
    io_A_Valid_1_delay_26_25 <= io_A_Valid_1_delay_25_26;
    io_A_Valid_1_delay_27_24 <= io_A_Valid_1_delay_26_25;
    io_A_Valid_1_delay_28_23 <= io_A_Valid_1_delay_27_24;
    io_A_Valid_1_delay_29_22 <= io_A_Valid_1_delay_28_23;
    io_A_Valid_1_delay_30_21 <= io_A_Valid_1_delay_29_22;
    io_A_Valid_1_delay_31_20 <= io_A_Valid_1_delay_30_21;
    io_A_Valid_1_delay_32_19 <= io_A_Valid_1_delay_31_20;
    io_A_Valid_1_delay_33_18 <= io_A_Valid_1_delay_32_19;
    io_A_Valid_1_delay_34_17 <= io_A_Valid_1_delay_33_18;
    io_A_Valid_1_delay_35_16 <= io_A_Valid_1_delay_34_17;
    io_A_Valid_1_delay_36_15 <= io_A_Valid_1_delay_35_16;
    io_A_Valid_1_delay_37_14 <= io_A_Valid_1_delay_36_15;
    io_A_Valid_1_delay_38_13 <= io_A_Valid_1_delay_37_14;
    io_A_Valid_1_delay_39_12 <= io_A_Valid_1_delay_38_13;
    io_A_Valid_1_delay_40_11 <= io_A_Valid_1_delay_39_12;
    io_A_Valid_1_delay_41_10 <= io_A_Valid_1_delay_40_11;
    io_A_Valid_1_delay_42_9 <= io_A_Valid_1_delay_41_10;
    io_A_Valid_1_delay_43_8 <= io_A_Valid_1_delay_42_9;
    io_A_Valid_1_delay_44_7 <= io_A_Valid_1_delay_43_8;
    io_A_Valid_1_delay_45_6 <= io_A_Valid_1_delay_44_7;
    io_A_Valid_1_delay_46_5 <= io_A_Valid_1_delay_45_6;
    io_A_Valid_1_delay_47_4 <= io_A_Valid_1_delay_46_5;
    io_A_Valid_1_delay_48_3 <= io_A_Valid_1_delay_47_4;
    io_A_Valid_1_delay_49_2 <= io_A_Valid_1_delay_48_3;
    io_A_Valid_1_delay_50_1 <= io_A_Valid_1_delay_49_2;
    io_A_Valid_1_delay_51 <= io_A_Valid_1_delay_50_1;
    io_B_Valid_51_delay_1 <= io_B_Valid_51;
    io_A_Valid_1_delay_1_51 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_50 <= io_A_Valid_1_delay_1_51;
    io_A_Valid_1_delay_3_49 <= io_A_Valid_1_delay_2_50;
    io_A_Valid_1_delay_4_48 <= io_A_Valid_1_delay_3_49;
    io_A_Valid_1_delay_5_47 <= io_A_Valid_1_delay_4_48;
    io_A_Valid_1_delay_6_46 <= io_A_Valid_1_delay_5_47;
    io_A_Valid_1_delay_7_45 <= io_A_Valid_1_delay_6_46;
    io_A_Valid_1_delay_8_44 <= io_A_Valid_1_delay_7_45;
    io_A_Valid_1_delay_9_43 <= io_A_Valid_1_delay_8_44;
    io_A_Valid_1_delay_10_42 <= io_A_Valid_1_delay_9_43;
    io_A_Valid_1_delay_11_41 <= io_A_Valid_1_delay_10_42;
    io_A_Valid_1_delay_12_40 <= io_A_Valid_1_delay_11_41;
    io_A_Valid_1_delay_13_39 <= io_A_Valid_1_delay_12_40;
    io_A_Valid_1_delay_14_38 <= io_A_Valid_1_delay_13_39;
    io_A_Valid_1_delay_15_37 <= io_A_Valid_1_delay_14_38;
    io_A_Valid_1_delay_16_36 <= io_A_Valid_1_delay_15_37;
    io_A_Valid_1_delay_17_35 <= io_A_Valid_1_delay_16_36;
    io_A_Valid_1_delay_18_34 <= io_A_Valid_1_delay_17_35;
    io_A_Valid_1_delay_19_33 <= io_A_Valid_1_delay_18_34;
    io_A_Valid_1_delay_20_32 <= io_A_Valid_1_delay_19_33;
    io_A_Valid_1_delay_21_31 <= io_A_Valid_1_delay_20_32;
    io_A_Valid_1_delay_22_30 <= io_A_Valid_1_delay_21_31;
    io_A_Valid_1_delay_23_29 <= io_A_Valid_1_delay_22_30;
    io_A_Valid_1_delay_24_28 <= io_A_Valid_1_delay_23_29;
    io_A_Valid_1_delay_25_27 <= io_A_Valid_1_delay_24_28;
    io_A_Valid_1_delay_26_26 <= io_A_Valid_1_delay_25_27;
    io_A_Valid_1_delay_27_25 <= io_A_Valid_1_delay_26_26;
    io_A_Valid_1_delay_28_24 <= io_A_Valid_1_delay_27_25;
    io_A_Valid_1_delay_29_23 <= io_A_Valid_1_delay_28_24;
    io_A_Valid_1_delay_30_22 <= io_A_Valid_1_delay_29_23;
    io_A_Valid_1_delay_31_21 <= io_A_Valid_1_delay_30_22;
    io_A_Valid_1_delay_32_20 <= io_A_Valid_1_delay_31_21;
    io_A_Valid_1_delay_33_19 <= io_A_Valid_1_delay_32_20;
    io_A_Valid_1_delay_34_18 <= io_A_Valid_1_delay_33_19;
    io_A_Valid_1_delay_35_17 <= io_A_Valid_1_delay_34_18;
    io_A_Valid_1_delay_36_16 <= io_A_Valid_1_delay_35_17;
    io_A_Valid_1_delay_37_15 <= io_A_Valid_1_delay_36_16;
    io_A_Valid_1_delay_38_14 <= io_A_Valid_1_delay_37_15;
    io_A_Valid_1_delay_39_13 <= io_A_Valid_1_delay_38_14;
    io_A_Valid_1_delay_40_12 <= io_A_Valid_1_delay_39_13;
    io_A_Valid_1_delay_41_11 <= io_A_Valid_1_delay_40_12;
    io_A_Valid_1_delay_42_10 <= io_A_Valid_1_delay_41_11;
    io_A_Valid_1_delay_43_9 <= io_A_Valid_1_delay_42_10;
    io_A_Valid_1_delay_44_8 <= io_A_Valid_1_delay_43_9;
    io_A_Valid_1_delay_45_7 <= io_A_Valid_1_delay_44_8;
    io_A_Valid_1_delay_46_6 <= io_A_Valid_1_delay_45_7;
    io_A_Valid_1_delay_47_5 <= io_A_Valid_1_delay_46_6;
    io_A_Valid_1_delay_48_4 <= io_A_Valid_1_delay_47_5;
    io_A_Valid_1_delay_49_3 <= io_A_Valid_1_delay_48_4;
    io_A_Valid_1_delay_50_2 <= io_A_Valid_1_delay_49_3;
    io_A_Valid_1_delay_51_1 <= io_A_Valid_1_delay_50_2;
    io_A_Valid_1_delay_52 <= io_A_Valid_1_delay_51_1;
    io_B_Valid_52_delay_1 <= io_B_Valid_52;
    io_A_Valid_1_delay_1_52 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_51 <= io_A_Valid_1_delay_1_52;
    io_A_Valid_1_delay_3_50 <= io_A_Valid_1_delay_2_51;
    io_A_Valid_1_delay_4_49 <= io_A_Valid_1_delay_3_50;
    io_A_Valid_1_delay_5_48 <= io_A_Valid_1_delay_4_49;
    io_A_Valid_1_delay_6_47 <= io_A_Valid_1_delay_5_48;
    io_A_Valid_1_delay_7_46 <= io_A_Valid_1_delay_6_47;
    io_A_Valid_1_delay_8_45 <= io_A_Valid_1_delay_7_46;
    io_A_Valid_1_delay_9_44 <= io_A_Valid_1_delay_8_45;
    io_A_Valid_1_delay_10_43 <= io_A_Valid_1_delay_9_44;
    io_A_Valid_1_delay_11_42 <= io_A_Valid_1_delay_10_43;
    io_A_Valid_1_delay_12_41 <= io_A_Valid_1_delay_11_42;
    io_A_Valid_1_delay_13_40 <= io_A_Valid_1_delay_12_41;
    io_A_Valid_1_delay_14_39 <= io_A_Valid_1_delay_13_40;
    io_A_Valid_1_delay_15_38 <= io_A_Valid_1_delay_14_39;
    io_A_Valid_1_delay_16_37 <= io_A_Valid_1_delay_15_38;
    io_A_Valid_1_delay_17_36 <= io_A_Valid_1_delay_16_37;
    io_A_Valid_1_delay_18_35 <= io_A_Valid_1_delay_17_36;
    io_A_Valid_1_delay_19_34 <= io_A_Valid_1_delay_18_35;
    io_A_Valid_1_delay_20_33 <= io_A_Valid_1_delay_19_34;
    io_A_Valid_1_delay_21_32 <= io_A_Valid_1_delay_20_33;
    io_A_Valid_1_delay_22_31 <= io_A_Valid_1_delay_21_32;
    io_A_Valid_1_delay_23_30 <= io_A_Valid_1_delay_22_31;
    io_A_Valid_1_delay_24_29 <= io_A_Valid_1_delay_23_30;
    io_A_Valid_1_delay_25_28 <= io_A_Valid_1_delay_24_29;
    io_A_Valid_1_delay_26_27 <= io_A_Valid_1_delay_25_28;
    io_A_Valid_1_delay_27_26 <= io_A_Valid_1_delay_26_27;
    io_A_Valid_1_delay_28_25 <= io_A_Valid_1_delay_27_26;
    io_A_Valid_1_delay_29_24 <= io_A_Valid_1_delay_28_25;
    io_A_Valid_1_delay_30_23 <= io_A_Valid_1_delay_29_24;
    io_A_Valid_1_delay_31_22 <= io_A_Valid_1_delay_30_23;
    io_A_Valid_1_delay_32_21 <= io_A_Valid_1_delay_31_22;
    io_A_Valid_1_delay_33_20 <= io_A_Valid_1_delay_32_21;
    io_A_Valid_1_delay_34_19 <= io_A_Valid_1_delay_33_20;
    io_A_Valid_1_delay_35_18 <= io_A_Valid_1_delay_34_19;
    io_A_Valid_1_delay_36_17 <= io_A_Valid_1_delay_35_18;
    io_A_Valid_1_delay_37_16 <= io_A_Valid_1_delay_36_17;
    io_A_Valid_1_delay_38_15 <= io_A_Valid_1_delay_37_16;
    io_A_Valid_1_delay_39_14 <= io_A_Valid_1_delay_38_15;
    io_A_Valid_1_delay_40_13 <= io_A_Valid_1_delay_39_14;
    io_A_Valid_1_delay_41_12 <= io_A_Valid_1_delay_40_13;
    io_A_Valid_1_delay_42_11 <= io_A_Valid_1_delay_41_12;
    io_A_Valid_1_delay_43_10 <= io_A_Valid_1_delay_42_11;
    io_A_Valid_1_delay_44_9 <= io_A_Valid_1_delay_43_10;
    io_A_Valid_1_delay_45_8 <= io_A_Valid_1_delay_44_9;
    io_A_Valid_1_delay_46_7 <= io_A_Valid_1_delay_45_8;
    io_A_Valid_1_delay_47_6 <= io_A_Valid_1_delay_46_7;
    io_A_Valid_1_delay_48_5 <= io_A_Valid_1_delay_47_6;
    io_A_Valid_1_delay_49_4 <= io_A_Valid_1_delay_48_5;
    io_A_Valid_1_delay_50_3 <= io_A_Valid_1_delay_49_4;
    io_A_Valid_1_delay_51_2 <= io_A_Valid_1_delay_50_3;
    io_A_Valid_1_delay_52_1 <= io_A_Valid_1_delay_51_2;
    io_A_Valid_1_delay_53 <= io_A_Valid_1_delay_52_1;
    io_B_Valid_53_delay_1 <= io_B_Valid_53;
    io_A_Valid_1_delay_1_53 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_52 <= io_A_Valid_1_delay_1_53;
    io_A_Valid_1_delay_3_51 <= io_A_Valid_1_delay_2_52;
    io_A_Valid_1_delay_4_50 <= io_A_Valid_1_delay_3_51;
    io_A_Valid_1_delay_5_49 <= io_A_Valid_1_delay_4_50;
    io_A_Valid_1_delay_6_48 <= io_A_Valid_1_delay_5_49;
    io_A_Valid_1_delay_7_47 <= io_A_Valid_1_delay_6_48;
    io_A_Valid_1_delay_8_46 <= io_A_Valid_1_delay_7_47;
    io_A_Valid_1_delay_9_45 <= io_A_Valid_1_delay_8_46;
    io_A_Valid_1_delay_10_44 <= io_A_Valid_1_delay_9_45;
    io_A_Valid_1_delay_11_43 <= io_A_Valid_1_delay_10_44;
    io_A_Valid_1_delay_12_42 <= io_A_Valid_1_delay_11_43;
    io_A_Valid_1_delay_13_41 <= io_A_Valid_1_delay_12_42;
    io_A_Valid_1_delay_14_40 <= io_A_Valid_1_delay_13_41;
    io_A_Valid_1_delay_15_39 <= io_A_Valid_1_delay_14_40;
    io_A_Valid_1_delay_16_38 <= io_A_Valid_1_delay_15_39;
    io_A_Valid_1_delay_17_37 <= io_A_Valid_1_delay_16_38;
    io_A_Valid_1_delay_18_36 <= io_A_Valid_1_delay_17_37;
    io_A_Valid_1_delay_19_35 <= io_A_Valid_1_delay_18_36;
    io_A_Valid_1_delay_20_34 <= io_A_Valid_1_delay_19_35;
    io_A_Valid_1_delay_21_33 <= io_A_Valid_1_delay_20_34;
    io_A_Valid_1_delay_22_32 <= io_A_Valid_1_delay_21_33;
    io_A_Valid_1_delay_23_31 <= io_A_Valid_1_delay_22_32;
    io_A_Valid_1_delay_24_30 <= io_A_Valid_1_delay_23_31;
    io_A_Valid_1_delay_25_29 <= io_A_Valid_1_delay_24_30;
    io_A_Valid_1_delay_26_28 <= io_A_Valid_1_delay_25_29;
    io_A_Valid_1_delay_27_27 <= io_A_Valid_1_delay_26_28;
    io_A_Valid_1_delay_28_26 <= io_A_Valid_1_delay_27_27;
    io_A_Valid_1_delay_29_25 <= io_A_Valid_1_delay_28_26;
    io_A_Valid_1_delay_30_24 <= io_A_Valid_1_delay_29_25;
    io_A_Valid_1_delay_31_23 <= io_A_Valid_1_delay_30_24;
    io_A_Valid_1_delay_32_22 <= io_A_Valid_1_delay_31_23;
    io_A_Valid_1_delay_33_21 <= io_A_Valid_1_delay_32_22;
    io_A_Valid_1_delay_34_20 <= io_A_Valid_1_delay_33_21;
    io_A_Valid_1_delay_35_19 <= io_A_Valid_1_delay_34_20;
    io_A_Valid_1_delay_36_18 <= io_A_Valid_1_delay_35_19;
    io_A_Valid_1_delay_37_17 <= io_A_Valid_1_delay_36_18;
    io_A_Valid_1_delay_38_16 <= io_A_Valid_1_delay_37_17;
    io_A_Valid_1_delay_39_15 <= io_A_Valid_1_delay_38_16;
    io_A_Valid_1_delay_40_14 <= io_A_Valid_1_delay_39_15;
    io_A_Valid_1_delay_41_13 <= io_A_Valid_1_delay_40_14;
    io_A_Valid_1_delay_42_12 <= io_A_Valid_1_delay_41_13;
    io_A_Valid_1_delay_43_11 <= io_A_Valid_1_delay_42_12;
    io_A_Valid_1_delay_44_10 <= io_A_Valid_1_delay_43_11;
    io_A_Valid_1_delay_45_9 <= io_A_Valid_1_delay_44_10;
    io_A_Valid_1_delay_46_8 <= io_A_Valid_1_delay_45_9;
    io_A_Valid_1_delay_47_7 <= io_A_Valid_1_delay_46_8;
    io_A_Valid_1_delay_48_6 <= io_A_Valid_1_delay_47_7;
    io_A_Valid_1_delay_49_5 <= io_A_Valid_1_delay_48_6;
    io_A_Valid_1_delay_50_4 <= io_A_Valid_1_delay_49_5;
    io_A_Valid_1_delay_51_3 <= io_A_Valid_1_delay_50_4;
    io_A_Valid_1_delay_52_2 <= io_A_Valid_1_delay_51_3;
    io_A_Valid_1_delay_53_1 <= io_A_Valid_1_delay_52_2;
    io_A_Valid_1_delay_54 <= io_A_Valid_1_delay_53_1;
    io_B_Valid_54_delay_1 <= io_B_Valid_54;
    io_A_Valid_1_delay_1_54 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_53 <= io_A_Valid_1_delay_1_54;
    io_A_Valid_1_delay_3_52 <= io_A_Valid_1_delay_2_53;
    io_A_Valid_1_delay_4_51 <= io_A_Valid_1_delay_3_52;
    io_A_Valid_1_delay_5_50 <= io_A_Valid_1_delay_4_51;
    io_A_Valid_1_delay_6_49 <= io_A_Valid_1_delay_5_50;
    io_A_Valid_1_delay_7_48 <= io_A_Valid_1_delay_6_49;
    io_A_Valid_1_delay_8_47 <= io_A_Valid_1_delay_7_48;
    io_A_Valid_1_delay_9_46 <= io_A_Valid_1_delay_8_47;
    io_A_Valid_1_delay_10_45 <= io_A_Valid_1_delay_9_46;
    io_A_Valid_1_delay_11_44 <= io_A_Valid_1_delay_10_45;
    io_A_Valid_1_delay_12_43 <= io_A_Valid_1_delay_11_44;
    io_A_Valid_1_delay_13_42 <= io_A_Valid_1_delay_12_43;
    io_A_Valid_1_delay_14_41 <= io_A_Valid_1_delay_13_42;
    io_A_Valid_1_delay_15_40 <= io_A_Valid_1_delay_14_41;
    io_A_Valid_1_delay_16_39 <= io_A_Valid_1_delay_15_40;
    io_A_Valid_1_delay_17_38 <= io_A_Valid_1_delay_16_39;
    io_A_Valid_1_delay_18_37 <= io_A_Valid_1_delay_17_38;
    io_A_Valid_1_delay_19_36 <= io_A_Valid_1_delay_18_37;
    io_A_Valid_1_delay_20_35 <= io_A_Valid_1_delay_19_36;
    io_A_Valid_1_delay_21_34 <= io_A_Valid_1_delay_20_35;
    io_A_Valid_1_delay_22_33 <= io_A_Valid_1_delay_21_34;
    io_A_Valid_1_delay_23_32 <= io_A_Valid_1_delay_22_33;
    io_A_Valid_1_delay_24_31 <= io_A_Valid_1_delay_23_32;
    io_A_Valid_1_delay_25_30 <= io_A_Valid_1_delay_24_31;
    io_A_Valid_1_delay_26_29 <= io_A_Valid_1_delay_25_30;
    io_A_Valid_1_delay_27_28 <= io_A_Valid_1_delay_26_29;
    io_A_Valid_1_delay_28_27 <= io_A_Valid_1_delay_27_28;
    io_A_Valid_1_delay_29_26 <= io_A_Valid_1_delay_28_27;
    io_A_Valid_1_delay_30_25 <= io_A_Valid_1_delay_29_26;
    io_A_Valid_1_delay_31_24 <= io_A_Valid_1_delay_30_25;
    io_A_Valid_1_delay_32_23 <= io_A_Valid_1_delay_31_24;
    io_A_Valid_1_delay_33_22 <= io_A_Valid_1_delay_32_23;
    io_A_Valid_1_delay_34_21 <= io_A_Valid_1_delay_33_22;
    io_A_Valid_1_delay_35_20 <= io_A_Valid_1_delay_34_21;
    io_A_Valid_1_delay_36_19 <= io_A_Valid_1_delay_35_20;
    io_A_Valid_1_delay_37_18 <= io_A_Valid_1_delay_36_19;
    io_A_Valid_1_delay_38_17 <= io_A_Valid_1_delay_37_18;
    io_A_Valid_1_delay_39_16 <= io_A_Valid_1_delay_38_17;
    io_A_Valid_1_delay_40_15 <= io_A_Valid_1_delay_39_16;
    io_A_Valid_1_delay_41_14 <= io_A_Valid_1_delay_40_15;
    io_A_Valid_1_delay_42_13 <= io_A_Valid_1_delay_41_14;
    io_A_Valid_1_delay_43_12 <= io_A_Valid_1_delay_42_13;
    io_A_Valid_1_delay_44_11 <= io_A_Valid_1_delay_43_12;
    io_A_Valid_1_delay_45_10 <= io_A_Valid_1_delay_44_11;
    io_A_Valid_1_delay_46_9 <= io_A_Valid_1_delay_45_10;
    io_A_Valid_1_delay_47_8 <= io_A_Valid_1_delay_46_9;
    io_A_Valid_1_delay_48_7 <= io_A_Valid_1_delay_47_8;
    io_A_Valid_1_delay_49_6 <= io_A_Valid_1_delay_48_7;
    io_A_Valid_1_delay_50_5 <= io_A_Valid_1_delay_49_6;
    io_A_Valid_1_delay_51_4 <= io_A_Valid_1_delay_50_5;
    io_A_Valid_1_delay_52_3 <= io_A_Valid_1_delay_51_4;
    io_A_Valid_1_delay_53_2 <= io_A_Valid_1_delay_52_3;
    io_A_Valid_1_delay_54_1 <= io_A_Valid_1_delay_53_2;
    io_A_Valid_1_delay_55 <= io_A_Valid_1_delay_54_1;
    io_B_Valid_55_delay_1 <= io_B_Valid_55;
    io_A_Valid_1_delay_1_55 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_54 <= io_A_Valid_1_delay_1_55;
    io_A_Valid_1_delay_3_53 <= io_A_Valid_1_delay_2_54;
    io_A_Valid_1_delay_4_52 <= io_A_Valid_1_delay_3_53;
    io_A_Valid_1_delay_5_51 <= io_A_Valid_1_delay_4_52;
    io_A_Valid_1_delay_6_50 <= io_A_Valid_1_delay_5_51;
    io_A_Valid_1_delay_7_49 <= io_A_Valid_1_delay_6_50;
    io_A_Valid_1_delay_8_48 <= io_A_Valid_1_delay_7_49;
    io_A_Valid_1_delay_9_47 <= io_A_Valid_1_delay_8_48;
    io_A_Valid_1_delay_10_46 <= io_A_Valid_1_delay_9_47;
    io_A_Valid_1_delay_11_45 <= io_A_Valid_1_delay_10_46;
    io_A_Valid_1_delay_12_44 <= io_A_Valid_1_delay_11_45;
    io_A_Valid_1_delay_13_43 <= io_A_Valid_1_delay_12_44;
    io_A_Valid_1_delay_14_42 <= io_A_Valid_1_delay_13_43;
    io_A_Valid_1_delay_15_41 <= io_A_Valid_1_delay_14_42;
    io_A_Valid_1_delay_16_40 <= io_A_Valid_1_delay_15_41;
    io_A_Valid_1_delay_17_39 <= io_A_Valid_1_delay_16_40;
    io_A_Valid_1_delay_18_38 <= io_A_Valid_1_delay_17_39;
    io_A_Valid_1_delay_19_37 <= io_A_Valid_1_delay_18_38;
    io_A_Valid_1_delay_20_36 <= io_A_Valid_1_delay_19_37;
    io_A_Valid_1_delay_21_35 <= io_A_Valid_1_delay_20_36;
    io_A_Valid_1_delay_22_34 <= io_A_Valid_1_delay_21_35;
    io_A_Valid_1_delay_23_33 <= io_A_Valid_1_delay_22_34;
    io_A_Valid_1_delay_24_32 <= io_A_Valid_1_delay_23_33;
    io_A_Valid_1_delay_25_31 <= io_A_Valid_1_delay_24_32;
    io_A_Valid_1_delay_26_30 <= io_A_Valid_1_delay_25_31;
    io_A_Valid_1_delay_27_29 <= io_A_Valid_1_delay_26_30;
    io_A_Valid_1_delay_28_28 <= io_A_Valid_1_delay_27_29;
    io_A_Valid_1_delay_29_27 <= io_A_Valid_1_delay_28_28;
    io_A_Valid_1_delay_30_26 <= io_A_Valid_1_delay_29_27;
    io_A_Valid_1_delay_31_25 <= io_A_Valid_1_delay_30_26;
    io_A_Valid_1_delay_32_24 <= io_A_Valid_1_delay_31_25;
    io_A_Valid_1_delay_33_23 <= io_A_Valid_1_delay_32_24;
    io_A_Valid_1_delay_34_22 <= io_A_Valid_1_delay_33_23;
    io_A_Valid_1_delay_35_21 <= io_A_Valid_1_delay_34_22;
    io_A_Valid_1_delay_36_20 <= io_A_Valid_1_delay_35_21;
    io_A_Valid_1_delay_37_19 <= io_A_Valid_1_delay_36_20;
    io_A_Valid_1_delay_38_18 <= io_A_Valid_1_delay_37_19;
    io_A_Valid_1_delay_39_17 <= io_A_Valid_1_delay_38_18;
    io_A_Valid_1_delay_40_16 <= io_A_Valid_1_delay_39_17;
    io_A_Valid_1_delay_41_15 <= io_A_Valid_1_delay_40_16;
    io_A_Valid_1_delay_42_14 <= io_A_Valid_1_delay_41_15;
    io_A_Valid_1_delay_43_13 <= io_A_Valid_1_delay_42_14;
    io_A_Valid_1_delay_44_12 <= io_A_Valid_1_delay_43_13;
    io_A_Valid_1_delay_45_11 <= io_A_Valid_1_delay_44_12;
    io_A_Valid_1_delay_46_10 <= io_A_Valid_1_delay_45_11;
    io_A_Valid_1_delay_47_9 <= io_A_Valid_1_delay_46_10;
    io_A_Valid_1_delay_48_8 <= io_A_Valid_1_delay_47_9;
    io_A_Valid_1_delay_49_7 <= io_A_Valid_1_delay_48_8;
    io_A_Valid_1_delay_50_6 <= io_A_Valid_1_delay_49_7;
    io_A_Valid_1_delay_51_5 <= io_A_Valid_1_delay_50_6;
    io_A_Valid_1_delay_52_4 <= io_A_Valid_1_delay_51_5;
    io_A_Valid_1_delay_53_3 <= io_A_Valid_1_delay_52_4;
    io_A_Valid_1_delay_54_2 <= io_A_Valid_1_delay_53_3;
    io_A_Valid_1_delay_55_1 <= io_A_Valid_1_delay_54_2;
    io_A_Valid_1_delay_56 <= io_A_Valid_1_delay_55_1;
    io_B_Valid_56_delay_1 <= io_B_Valid_56;
    io_A_Valid_1_delay_1_56 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_55 <= io_A_Valid_1_delay_1_56;
    io_A_Valid_1_delay_3_54 <= io_A_Valid_1_delay_2_55;
    io_A_Valid_1_delay_4_53 <= io_A_Valid_1_delay_3_54;
    io_A_Valid_1_delay_5_52 <= io_A_Valid_1_delay_4_53;
    io_A_Valid_1_delay_6_51 <= io_A_Valid_1_delay_5_52;
    io_A_Valid_1_delay_7_50 <= io_A_Valid_1_delay_6_51;
    io_A_Valid_1_delay_8_49 <= io_A_Valid_1_delay_7_50;
    io_A_Valid_1_delay_9_48 <= io_A_Valid_1_delay_8_49;
    io_A_Valid_1_delay_10_47 <= io_A_Valid_1_delay_9_48;
    io_A_Valid_1_delay_11_46 <= io_A_Valid_1_delay_10_47;
    io_A_Valid_1_delay_12_45 <= io_A_Valid_1_delay_11_46;
    io_A_Valid_1_delay_13_44 <= io_A_Valid_1_delay_12_45;
    io_A_Valid_1_delay_14_43 <= io_A_Valid_1_delay_13_44;
    io_A_Valid_1_delay_15_42 <= io_A_Valid_1_delay_14_43;
    io_A_Valid_1_delay_16_41 <= io_A_Valid_1_delay_15_42;
    io_A_Valid_1_delay_17_40 <= io_A_Valid_1_delay_16_41;
    io_A_Valid_1_delay_18_39 <= io_A_Valid_1_delay_17_40;
    io_A_Valid_1_delay_19_38 <= io_A_Valid_1_delay_18_39;
    io_A_Valid_1_delay_20_37 <= io_A_Valid_1_delay_19_38;
    io_A_Valid_1_delay_21_36 <= io_A_Valid_1_delay_20_37;
    io_A_Valid_1_delay_22_35 <= io_A_Valid_1_delay_21_36;
    io_A_Valid_1_delay_23_34 <= io_A_Valid_1_delay_22_35;
    io_A_Valid_1_delay_24_33 <= io_A_Valid_1_delay_23_34;
    io_A_Valid_1_delay_25_32 <= io_A_Valid_1_delay_24_33;
    io_A_Valid_1_delay_26_31 <= io_A_Valid_1_delay_25_32;
    io_A_Valid_1_delay_27_30 <= io_A_Valid_1_delay_26_31;
    io_A_Valid_1_delay_28_29 <= io_A_Valid_1_delay_27_30;
    io_A_Valid_1_delay_29_28 <= io_A_Valid_1_delay_28_29;
    io_A_Valid_1_delay_30_27 <= io_A_Valid_1_delay_29_28;
    io_A_Valid_1_delay_31_26 <= io_A_Valid_1_delay_30_27;
    io_A_Valid_1_delay_32_25 <= io_A_Valid_1_delay_31_26;
    io_A_Valid_1_delay_33_24 <= io_A_Valid_1_delay_32_25;
    io_A_Valid_1_delay_34_23 <= io_A_Valid_1_delay_33_24;
    io_A_Valid_1_delay_35_22 <= io_A_Valid_1_delay_34_23;
    io_A_Valid_1_delay_36_21 <= io_A_Valid_1_delay_35_22;
    io_A_Valid_1_delay_37_20 <= io_A_Valid_1_delay_36_21;
    io_A_Valid_1_delay_38_19 <= io_A_Valid_1_delay_37_20;
    io_A_Valid_1_delay_39_18 <= io_A_Valid_1_delay_38_19;
    io_A_Valid_1_delay_40_17 <= io_A_Valid_1_delay_39_18;
    io_A_Valid_1_delay_41_16 <= io_A_Valid_1_delay_40_17;
    io_A_Valid_1_delay_42_15 <= io_A_Valid_1_delay_41_16;
    io_A_Valid_1_delay_43_14 <= io_A_Valid_1_delay_42_15;
    io_A_Valid_1_delay_44_13 <= io_A_Valid_1_delay_43_14;
    io_A_Valid_1_delay_45_12 <= io_A_Valid_1_delay_44_13;
    io_A_Valid_1_delay_46_11 <= io_A_Valid_1_delay_45_12;
    io_A_Valid_1_delay_47_10 <= io_A_Valid_1_delay_46_11;
    io_A_Valid_1_delay_48_9 <= io_A_Valid_1_delay_47_10;
    io_A_Valid_1_delay_49_8 <= io_A_Valid_1_delay_48_9;
    io_A_Valid_1_delay_50_7 <= io_A_Valid_1_delay_49_8;
    io_A_Valid_1_delay_51_6 <= io_A_Valid_1_delay_50_7;
    io_A_Valid_1_delay_52_5 <= io_A_Valid_1_delay_51_6;
    io_A_Valid_1_delay_53_4 <= io_A_Valid_1_delay_52_5;
    io_A_Valid_1_delay_54_3 <= io_A_Valid_1_delay_53_4;
    io_A_Valid_1_delay_55_2 <= io_A_Valid_1_delay_54_3;
    io_A_Valid_1_delay_56_1 <= io_A_Valid_1_delay_55_2;
    io_A_Valid_1_delay_57 <= io_A_Valid_1_delay_56_1;
    io_B_Valid_57_delay_1 <= io_B_Valid_57;
    io_A_Valid_1_delay_1_57 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_56 <= io_A_Valid_1_delay_1_57;
    io_A_Valid_1_delay_3_55 <= io_A_Valid_1_delay_2_56;
    io_A_Valid_1_delay_4_54 <= io_A_Valid_1_delay_3_55;
    io_A_Valid_1_delay_5_53 <= io_A_Valid_1_delay_4_54;
    io_A_Valid_1_delay_6_52 <= io_A_Valid_1_delay_5_53;
    io_A_Valid_1_delay_7_51 <= io_A_Valid_1_delay_6_52;
    io_A_Valid_1_delay_8_50 <= io_A_Valid_1_delay_7_51;
    io_A_Valid_1_delay_9_49 <= io_A_Valid_1_delay_8_50;
    io_A_Valid_1_delay_10_48 <= io_A_Valid_1_delay_9_49;
    io_A_Valid_1_delay_11_47 <= io_A_Valid_1_delay_10_48;
    io_A_Valid_1_delay_12_46 <= io_A_Valid_1_delay_11_47;
    io_A_Valid_1_delay_13_45 <= io_A_Valid_1_delay_12_46;
    io_A_Valid_1_delay_14_44 <= io_A_Valid_1_delay_13_45;
    io_A_Valid_1_delay_15_43 <= io_A_Valid_1_delay_14_44;
    io_A_Valid_1_delay_16_42 <= io_A_Valid_1_delay_15_43;
    io_A_Valid_1_delay_17_41 <= io_A_Valid_1_delay_16_42;
    io_A_Valid_1_delay_18_40 <= io_A_Valid_1_delay_17_41;
    io_A_Valid_1_delay_19_39 <= io_A_Valid_1_delay_18_40;
    io_A_Valid_1_delay_20_38 <= io_A_Valid_1_delay_19_39;
    io_A_Valid_1_delay_21_37 <= io_A_Valid_1_delay_20_38;
    io_A_Valid_1_delay_22_36 <= io_A_Valid_1_delay_21_37;
    io_A_Valid_1_delay_23_35 <= io_A_Valid_1_delay_22_36;
    io_A_Valid_1_delay_24_34 <= io_A_Valid_1_delay_23_35;
    io_A_Valid_1_delay_25_33 <= io_A_Valid_1_delay_24_34;
    io_A_Valid_1_delay_26_32 <= io_A_Valid_1_delay_25_33;
    io_A_Valid_1_delay_27_31 <= io_A_Valid_1_delay_26_32;
    io_A_Valid_1_delay_28_30 <= io_A_Valid_1_delay_27_31;
    io_A_Valid_1_delay_29_29 <= io_A_Valid_1_delay_28_30;
    io_A_Valid_1_delay_30_28 <= io_A_Valid_1_delay_29_29;
    io_A_Valid_1_delay_31_27 <= io_A_Valid_1_delay_30_28;
    io_A_Valid_1_delay_32_26 <= io_A_Valid_1_delay_31_27;
    io_A_Valid_1_delay_33_25 <= io_A_Valid_1_delay_32_26;
    io_A_Valid_1_delay_34_24 <= io_A_Valid_1_delay_33_25;
    io_A_Valid_1_delay_35_23 <= io_A_Valid_1_delay_34_24;
    io_A_Valid_1_delay_36_22 <= io_A_Valid_1_delay_35_23;
    io_A_Valid_1_delay_37_21 <= io_A_Valid_1_delay_36_22;
    io_A_Valid_1_delay_38_20 <= io_A_Valid_1_delay_37_21;
    io_A_Valid_1_delay_39_19 <= io_A_Valid_1_delay_38_20;
    io_A_Valid_1_delay_40_18 <= io_A_Valid_1_delay_39_19;
    io_A_Valid_1_delay_41_17 <= io_A_Valid_1_delay_40_18;
    io_A_Valid_1_delay_42_16 <= io_A_Valid_1_delay_41_17;
    io_A_Valid_1_delay_43_15 <= io_A_Valid_1_delay_42_16;
    io_A_Valid_1_delay_44_14 <= io_A_Valid_1_delay_43_15;
    io_A_Valid_1_delay_45_13 <= io_A_Valid_1_delay_44_14;
    io_A_Valid_1_delay_46_12 <= io_A_Valid_1_delay_45_13;
    io_A_Valid_1_delay_47_11 <= io_A_Valid_1_delay_46_12;
    io_A_Valid_1_delay_48_10 <= io_A_Valid_1_delay_47_11;
    io_A_Valid_1_delay_49_9 <= io_A_Valid_1_delay_48_10;
    io_A_Valid_1_delay_50_8 <= io_A_Valid_1_delay_49_9;
    io_A_Valid_1_delay_51_7 <= io_A_Valid_1_delay_50_8;
    io_A_Valid_1_delay_52_6 <= io_A_Valid_1_delay_51_7;
    io_A_Valid_1_delay_53_5 <= io_A_Valid_1_delay_52_6;
    io_A_Valid_1_delay_54_4 <= io_A_Valid_1_delay_53_5;
    io_A_Valid_1_delay_55_3 <= io_A_Valid_1_delay_54_4;
    io_A_Valid_1_delay_56_2 <= io_A_Valid_1_delay_55_3;
    io_A_Valid_1_delay_57_1 <= io_A_Valid_1_delay_56_2;
    io_A_Valid_1_delay_58 <= io_A_Valid_1_delay_57_1;
    io_B_Valid_58_delay_1 <= io_B_Valid_58;
    io_A_Valid_1_delay_1_58 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_57 <= io_A_Valid_1_delay_1_58;
    io_A_Valid_1_delay_3_56 <= io_A_Valid_1_delay_2_57;
    io_A_Valid_1_delay_4_55 <= io_A_Valid_1_delay_3_56;
    io_A_Valid_1_delay_5_54 <= io_A_Valid_1_delay_4_55;
    io_A_Valid_1_delay_6_53 <= io_A_Valid_1_delay_5_54;
    io_A_Valid_1_delay_7_52 <= io_A_Valid_1_delay_6_53;
    io_A_Valid_1_delay_8_51 <= io_A_Valid_1_delay_7_52;
    io_A_Valid_1_delay_9_50 <= io_A_Valid_1_delay_8_51;
    io_A_Valid_1_delay_10_49 <= io_A_Valid_1_delay_9_50;
    io_A_Valid_1_delay_11_48 <= io_A_Valid_1_delay_10_49;
    io_A_Valid_1_delay_12_47 <= io_A_Valid_1_delay_11_48;
    io_A_Valid_1_delay_13_46 <= io_A_Valid_1_delay_12_47;
    io_A_Valid_1_delay_14_45 <= io_A_Valid_1_delay_13_46;
    io_A_Valid_1_delay_15_44 <= io_A_Valid_1_delay_14_45;
    io_A_Valid_1_delay_16_43 <= io_A_Valid_1_delay_15_44;
    io_A_Valid_1_delay_17_42 <= io_A_Valid_1_delay_16_43;
    io_A_Valid_1_delay_18_41 <= io_A_Valid_1_delay_17_42;
    io_A_Valid_1_delay_19_40 <= io_A_Valid_1_delay_18_41;
    io_A_Valid_1_delay_20_39 <= io_A_Valid_1_delay_19_40;
    io_A_Valid_1_delay_21_38 <= io_A_Valid_1_delay_20_39;
    io_A_Valid_1_delay_22_37 <= io_A_Valid_1_delay_21_38;
    io_A_Valid_1_delay_23_36 <= io_A_Valid_1_delay_22_37;
    io_A_Valid_1_delay_24_35 <= io_A_Valid_1_delay_23_36;
    io_A_Valid_1_delay_25_34 <= io_A_Valid_1_delay_24_35;
    io_A_Valid_1_delay_26_33 <= io_A_Valid_1_delay_25_34;
    io_A_Valid_1_delay_27_32 <= io_A_Valid_1_delay_26_33;
    io_A_Valid_1_delay_28_31 <= io_A_Valid_1_delay_27_32;
    io_A_Valid_1_delay_29_30 <= io_A_Valid_1_delay_28_31;
    io_A_Valid_1_delay_30_29 <= io_A_Valid_1_delay_29_30;
    io_A_Valid_1_delay_31_28 <= io_A_Valid_1_delay_30_29;
    io_A_Valid_1_delay_32_27 <= io_A_Valid_1_delay_31_28;
    io_A_Valid_1_delay_33_26 <= io_A_Valid_1_delay_32_27;
    io_A_Valid_1_delay_34_25 <= io_A_Valid_1_delay_33_26;
    io_A_Valid_1_delay_35_24 <= io_A_Valid_1_delay_34_25;
    io_A_Valid_1_delay_36_23 <= io_A_Valid_1_delay_35_24;
    io_A_Valid_1_delay_37_22 <= io_A_Valid_1_delay_36_23;
    io_A_Valid_1_delay_38_21 <= io_A_Valid_1_delay_37_22;
    io_A_Valid_1_delay_39_20 <= io_A_Valid_1_delay_38_21;
    io_A_Valid_1_delay_40_19 <= io_A_Valid_1_delay_39_20;
    io_A_Valid_1_delay_41_18 <= io_A_Valid_1_delay_40_19;
    io_A_Valid_1_delay_42_17 <= io_A_Valid_1_delay_41_18;
    io_A_Valid_1_delay_43_16 <= io_A_Valid_1_delay_42_17;
    io_A_Valid_1_delay_44_15 <= io_A_Valid_1_delay_43_16;
    io_A_Valid_1_delay_45_14 <= io_A_Valid_1_delay_44_15;
    io_A_Valid_1_delay_46_13 <= io_A_Valid_1_delay_45_14;
    io_A_Valid_1_delay_47_12 <= io_A_Valid_1_delay_46_13;
    io_A_Valid_1_delay_48_11 <= io_A_Valid_1_delay_47_12;
    io_A_Valid_1_delay_49_10 <= io_A_Valid_1_delay_48_11;
    io_A_Valid_1_delay_50_9 <= io_A_Valid_1_delay_49_10;
    io_A_Valid_1_delay_51_8 <= io_A_Valid_1_delay_50_9;
    io_A_Valid_1_delay_52_7 <= io_A_Valid_1_delay_51_8;
    io_A_Valid_1_delay_53_6 <= io_A_Valid_1_delay_52_7;
    io_A_Valid_1_delay_54_5 <= io_A_Valid_1_delay_53_6;
    io_A_Valid_1_delay_55_4 <= io_A_Valid_1_delay_54_5;
    io_A_Valid_1_delay_56_3 <= io_A_Valid_1_delay_55_4;
    io_A_Valid_1_delay_57_2 <= io_A_Valid_1_delay_56_3;
    io_A_Valid_1_delay_58_1 <= io_A_Valid_1_delay_57_2;
    io_A_Valid_1_delay_59 <= io_A_Valid_1_delay_58_1;
    io_B_Valid_59_delay_1 <= io_B_Valid_59;
    io_A_Valid_1_delay_1_59 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_58 <= io_A_Valid_1_delay_1_59;
    io_A_Valid_1_delay_3_57 <= io_A_Valid_1_delay_2_58;
    io_A_Valid_1_delay_4_56 <= io_A_Valid_1_delay_3_57;
    io_A_Valid_1_delay_5_55 <= io_A_Valid_1_delay_4_56;
    io_A_Valid_1_delay_6_54 <= io_A_Valid_1_delay_5_55;
    io_A_Valid_1_delay_7_53 <= io_A_Valid_1_delay_6_54;
    io_A_Valid_1_delay_8_52 <= io_A_Valid_1_delay_7_53;
    io_A_Valid_1_delay_9_51 <= io_A_Valid_1_delay_8_52;
    io_A_Valid_1_delay_10_50 <= io_A_Valid_1_delay_9_51;
    io_A_Valid_1_delay_11_49 <= io_A_Valid_1_delay_10_50;
    io_A_Valid_1_delay_12_48 <= io_A_Valid_1_delay_11_49;
    io_A_Valid_1_delay_13_47 <= io_A_Valid_1_delay_12_48;
    io_A_Valid_1_delay_14_46 <= io_A_Valid_1_delay_13_47;
    io_A_Valid_1_delay_15_45 <= io_A_Valid_1_delay_14_46;
    io_A_Valid_1_delay_16_44 <= io_A_Valid_1_delay_15_45;
    io_A_Valid_1_delay_17_43 <= io_A_Valid_1_delay_16_44;
    io_A_Valid_1_delay_18_42 <= io_A_Valid_1_delay_17_43;
    io_A_Valid_1_delay_19_41 <= io_A_Valid_1_delay_18_42;
    io_A_Valid_1_delay_20_40 <= io_A_Valid_1_delay_19_41;
    io_A_Valid_1_delay_21_39 <= io_A_Valid_1_delay_20_40;
    io_A_Valid_1_delay_22_38 <= io_A_Valid_1_delay_21_39;
    io_A_Valid_1_delay_23_37 <= io_A_Valid_1_delay_22_38;
    io_A_Valid_1_delay_24_36 <= io_A_Valid_1_delay_23_37;
    io_A_Valid_1_delay_25_35 <= io_A_Valid_1_delay_24_36;
    io_A_Valid_1_delay_26_34 <= io_A_Valid_1_delay_25_35;
    io_A_Valid_1_delay_27_33 <= io_A_Valid_1_delay_26_34;
    io_A_Valid_1_delay_28_32 <= io_A_Valid_1_delay_27_33;
    io_A_Valid_1_delay_29_31 <= io_A_Valid_1_delay_28_32;
    io_A_Valid_1_delay_30_30 <= io_A_Valid_1_delay_29_31;
    io_A_Valid_1_delay_31_29 <= io_A_Valid_1_delay_30_30;
    io_A_Valid_1_delay_32_28 <= io_A_Valid_1_delay_31_29;
    io_A_Valid_1_delay_33_27 <= io_A_Valid_1_delay_32_28;
    io_A_Valid_1_delay_34_26 <= io_A_Valid_1_delay_33_27;
    io_A_Valid_1_delay_35_25 <= io_A_Valid_1_delay_34_26;
    io_A_Valid_1_delay_36_24 <= io_A_Valid_1_delay_35_25;
    io_A_Valid_1_delay_37_23 <= io_A_Valid_1_delay_36_24;
    io_A_Valid_1_delay_38_22 <= io_A_Valid_1_delay_37_23;
    io_A_Valid_1_delay_39_21 <= io_A_Valid_1_delay_38_22;
    io_A_Valid_1_delay_40_20 <= io_A_Valid_1_delay_39_21;
    io_A_Valid_1_delay_41_19 <= io_A_Valid_1_delay_40_20;
    io_A_Valid_1_delay_42_18 <= io_A_Valid_1_delay_41_19;
    io_A_Valid_1_delay_43_17 <= io_A_Valid_1_delay_42_18;
    io_A_Valid_1_delay_44_16 <= io_A_Valid_1_delay_43_17;
    io_A_Valid_1_delay_45_15 <= io_A_Valid_1_delay_44_16;
    io_A_Valid_1_delay_46_14 <= io_A_Valid_1_delay_45_15;
    io_A_Valid_1_delay_47_13 <= io_A_Valid_1_delay_46_14;
    io_A_Valid_1_delay_48_12 <= io_A_Valid_1_delay_47_13;
    io_A_Valid_1_delay_49_11 <= io_A_Valid_1_delay_48_12;
    io_A_Valid_1_delay_50_10 <= io_A_Valid_1_delay_49_11;
    io_A_Valid_1_delay_51_9 <= io_A_Valid_1_delay_50_10;
    io_A_Valid_1_delay_52_8 <= io_A_Valid_1_delay_51_9;
    io_A_Valid_1_delay_53_7 <= io_A_Valid_1_delay_52_8;
    io_A_Valid_1_delay_54_6 <= io_A_Valid_1_delay_53_7;
    io_A_Valid_1_delay_55_5 <= io_A_Valid_1_delay_54_6;
    io_A_Valid_1_delay_56_4 <= io_A_Valid_1_delay_55_5;
    io_A_Valid_1_delay_57_3 <= io_A_Valid_1_delay_56_4;
    io_A_Valid_1_delay_58_2 <= io_A_Valid_1_delay_57_3;
    io_A_Valid_1_delay_59_1 <= io_A_Valid_1_delay_58_2;
    io_A_Valid_1_delay_60 <= io_A_Valid_1_delay_59_1;
    io_B_Valid_60_delay_1 <= io_B_Valid_60;
    io_A_Valid_1_delay_1_60 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_59 <= io_A_Valid_1_delay_1_60;
    io_A_Valid_1_delay_3_58 <= io_A_Valid_1_delay_2_59;
    io_A_Valid_1_delay_4_57 <= io_A_Valid_1_delay_3_58;
    io_A_Valid_1_delay_5_56 <= io_A_Valid_1_delay_4_57;
    io_A_Valid_1_delay_6_55 <= io_A_Valid_1_delay_5_56;
    io_A_Valid_1_delay_7_54 <= io_A_Valid_1_delay_6_55;
    io_A_Valid_1_delay_8_53 <= io_A_Valid_1_delay_7_54;
    io_A_Valid_1_delay_9_52 <= io_A_Valid_1_delay_8_53;
    io_A_Valid_1_delay_10_51 <= io_A_Valid_1_delay_9_52;
    io_A_Valid_1_delay_11_50 <= io_A_Valid_1_delay_10_51;
    io_A_Valid_1_delay_12_49 <= io_A_Valid_1_delay_11_50;
    io_A_Valid_1_delay_13_48 <= io_A_Valid_1_delay_12_49;
    io_A_Valid_1_delay_14_47 <= io_A_Valid_1_delay_13_48;
    io_A_Valid_1_delay_15_46 <= io_A_Valid_1_delay_14_47;
    io_A_Valid_1_delay_16_45 <= io_A_Valid_1_delay_15_46;
    io_A_Valid_1_delay_17_44 <= io_A_Valid_1_delay_16_45;
    io_A_Valid_1_delay_18_43 <= io_A_Valid_1_delay_17_44;
    io_A_Valid_1_delay_19_42 <= io_A_Valid_1_delay_18_43;
    io_A_Valid_1_delay_20_41 <= io_A_Valid_1_delay_19_42;
    io_A_Valid_1_delay_21_40 <= io_A_Valid_1_delay_20_41;
    io_A_Valid_1_delay_22_39 <= io_A_Valid_1_delay_21_40;
    io_A_Valid_1_delay_23_38 <= io_A_Valid_1_delay_22_39;
    io_A_Valid_1_delay_24_37 <= io_A_Valid_1_delay_23_38;
    io_A_Valid_1_delay_25_36 <= io_A_Valid_1_delay_24_37;
    io_A_Valid_1_delay_26_35 <= io_A_Valid_1_delay_25_36;
    io_A_Valid_1_delay_27_34 <= io_A_Valid_1_delay_26_35;
    io_A_Valid_1_delay_28_33 <= io_A_Valid_1_delay_27_34;
    io_A_Valid_1_delay_29_32 <= io_A_Valid_1_delay_28_33;
    io_A_Valid_1_delay_30_31 <= io_A_Valid_1_delay_29_32;
    io_A_Valid_1_delay_31_30 <= io_A_Valid_1_delay_30_31;
    io_A_Valid_1_delay_32_29 <= io_A_Valid_1_delay_31_30;
    io_A_Valid_1_delay_33_28 <= io_A_Valid_1_delay_32_29;
    io_A_Valid_1_delay_34_27 <= io_A_Valid_1_delay_33_28;
    io_A_Valid_1_delay_35_26 <= io_A_Valid_1_delay_34_27;
    io_A_Valid_1_delay_36_25 <= io_A_Valid_1_delay_35_26;
    io_A_Valid_1_delay_37_24 <= io_A_Valid_1_delay_36_25;
    io_A_Valid_1_delay_38_23 <= io_A_Valid_1_delay_37_24;
    io_A_Valid_1_delay_39_22 <= io_A_Valid_1_delay_38_23;
    io_A_Valid_1_delay_40_21 <= io_A_Valid_1_delay_39_22;
    io_A_Valid_1_delay_41_20 <= io_A_Valid_1_delay_40_21;
    io_A_Valid_1_delay_42_19 <= io_A_Valid_1_delay_41_20;
    io_A_Valid_1_delay_43_18 <= io_A_Valid_1_delay_42_19;
    io_A_Valid_1_delay_44_17 <= io_A_Valid_1_delay_43_18;
    io_A_Valid_1_delay_45_16 <= io_A_Valid_1_delay_44_17;
    io_A_Valid_1_delay_46_15 <= io_A_Valid_1_delay_45_16;
    io_A_Valid_1_delay_47_14 <= io_A_Valid_1_delay_46_15;
    io_A_Valid_1_delay_48_13 <= io_A_Valid_1_delay_47_14;
    io_A_Valid_1_delay_49_12 <= io_A_Valid_1_delay_48_13;
    io_A_Valid_1_delay_50_11 <= io_A_Valid_1_delay_49_12;
    io_A_Valid_1_delay_51_10 <= io_A_Valid_1_delay_50_11;
    io_A_Valid_1_delay_52_9 <= io_A_Valid_1_delay_51_10;
    io_A_Valid_1_delay_53_8 <= io_A_Valid_1_delay_52_9;
    io_A_Valid_1_delay_54_7 <= io_A_Valid_1_delay_53_8;
    io_A_Valid_1_delay_55_6 <= io_A_Valid_1_delay_54_7;
    io_A_Valid_1_delay_56_5 <= io_A_Valid_1_delay_55_6;
    io_A_Valid_1_delay_57_4 <= io_A_Valid_1_delay_56_5;
    io_A_Valid_1_delay_58_3 <= io_A_Valid_1_delay_57_4;
    io_A_Valid_1_delay_59_2 <= io_A_Valid_1_delay_58_3;
    io_A_Valid_1_delay_60_1 <= io_A_Valid_1_delay_59_2;
    io_A_Valid_1_delay_61 <= io_A_Valid_1_delay_60_1;
    io_B_Valid_61_delay_1 <= io_B_Valid_61;
    io_A_Valid_1_delay_1_61 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_60 <= io_A_Valid_1_delay_1_61;
    io_A_Valid_1_delay_3_59 <= io_A_Valid_1_delay_2_60;
    io_A_Valid_1_delay_4_58 <= io_A_Valid_1_delay_3_59;
    io_A_Valid_1_delay_5_57 <= io_A_Valid_1_delay_4_58;
    io_A_Valid_1_delay_6_56 <= io_A_Valid_1_delay_5_57;
    io_A_Valid_1_delay_7_55 <= io_A_Valid_1_delay_6_56;
    io_A_Valid_1_delay_8_54 <= io_A_Valid_1_delay_7_55;
    io_A_Valid_1_delay_9_53 <= io_A_Valid_1_delay_8_54;
    io_A_Valid_1_delay_10_52 <= io_A_Valid_1_delay_9_53;
    io_A_Valid_1_delay_11_51 <= io_A_Valid_1_delay_10_52;
    io_A_Valid_1_delay_12_50 <= io_A_Valid_1_delay_11_51;
    io_A_Valid_1_delay_13_49 <= io_A_Valid_1_delay_12_50;
    io_A_Valid_1_delay_14_48 <= io_A_Valid_1_delay_13_49;
    io_A_Valid_1_delay_15_47 <= io_A_Valid_1_delay_14_48;
    io_A_Valid_1_delay_16_46 <= io_A_Valid_1_delay_15_47;
    io_A_Valid_1_delay_17_45 <= io_A_Valid_1_delay_16_46;
    io_A_Valid_1_delay_18_44 <= io_A_Valid_1_delay_17_45;
    io_A_Valid_1_delay_19_43 <= io_A_Valid_1_delay_18_44;
    io_A_Valid_1_delay_20_42 <= io_A_Valid_1_delay_19_43;
    io_A_Valid_1_delay_21_41 <= io_A_Valid_1_delay_20_42;
    io_A_Valid_1_delay_22_40 <= io_A_Valid_1_delay_21_41;
    io_A_Valid_1_delay_23_39 <= io_A_Valid_1_delay_22_40;
    io_A_Valid_1_delay_24_38 <= io_A_Valid_1_delay_23_39;
    io_A_Valid_1_delay_25_37 <= io_A_Valid_1_delay_24_38;
    io_A_Valid_1_delay_26_36 <= io_A_Valid_1_delay_25_37;
    io_A_Valid_1_delay_27_35 <= io_A_Valid_1_delay_26_36;
    io_A_Valid_1_delay_28_34 <= io_A_Valid_1_delay_27_35;
    io_A_Valid_1_delay_29_33 <= io_A_Valid_1_delay_28_34;
    io_A_Valid_1_delay_30_32 <= io_A_Valid_1_delay_29_33;
    io_A_Valid_1_delay_31_31 <= io_A_Valid_1_delay_30_32;
    io_A_Valid_1_delay_32_30 <= io_A_Valid_1_delay_31_31;
    io_A_Valid_1_delay_33_29 <= io_A_Valid_1_delay_32_30;
    io_A_Valid_1_delay_34_28 <= io_A_Valid_1_delay_33_29;
    io_A_Valid_1_delay_35_27 <= io_A_Valid_1_delay_34_28;
    io_A_Valid_1_delay_36_26 <= io_A_Valid_1_delay_35_27;
    io_A_Valid_1_delay_37_25 <= io_A_Valid_1_delay_36_26;
    io_A_Valid_1_delay_38_24 <= io_A_Valid_1_delay_37_25;
    io_A_Valid_1_delay_39_23 <= io_A_Valid_1_delay_38_24;
    io_A_Valid_1_delay_40_22 <= io_A_Valid_1_delay_39_23;
    io_A_Valid_1_delay_41_21 <= io_A_Valid_1_delay_40_22;
    io_A_Valid_1_delay_42_20 <= io_A_Valid_1_delay_41_21;
    io_A_Valid_1_delay_43_19 <= io_A_Valid_1_delay_42_20;
    io_A_Valid_1_delay_44_18 <= io_A_Valid_1_delay_43_19;
    io_A_Valid_1_delay_45_17 <= io_A_Valid_1_delay_44_18;
    io_A_Valid_1_delay_46_16 <= io_A_Valid_1_delay_45_17;
    io_A_Valid_1_delay_47_15 <= io_A_Valid_1_delay_46_16;
    io_A_Valid_1_delay_48_14 <= io_A_Valid_1_delay_47_15;
    io_A_Valid_1_delay_49_13 <= io_A_Valid_1_delay_48_14;
    io_A_Valid_1_delay_50_12 <= io_A_Valid_1_delay_49_13;
    io_A_Valid_1_delay_51_11 <= io_A_Valid_1_delay_50_12;
    io_A_Valid_1_delay_52_10 <= io_A_Valid_1_delay_51_11;
    io_A_Valid_1_delay_53_9 <= io_A_Valid_1_delay_52_10;
    io_A_Valid_1_delay_54_8 <= io_A_Valid_1_delay_53_9;
    io_A_Valid_1_delay_55_7 <= io_A_Valid_1_delay_54_8;
    io_A_Valid_1_delay_56_6 <= io_A_Valid_1_delay_55_7;
    io_A_Valid_1_delay_57_5 <= io_A_Valid_1_delay_56_6;
    io_A_Valid_1_delay_58_4 <= io_A_Valid_1_delay_57_5;
    io_A_Valid_1_delay_59_3 <= io_A_Valid_1_delay_58_4;
    io_A_Valid_1_delay_60_2 <= io_A_Valid_1_delay_59_3;
    io_A_Valid_1_delay_61_1 <= io_A_Valid_1_delay_60_2;
    io_A_Valid_1_delay_62 <= io_A_Valid_1_delay_61_1;
    io_B_Valid_62_delay_1 <= io_B_Valid_62;
    io_A_Valid_1_delay_1_62 <= io_A_Valid_1;
    io_A_Valid_1_delay_2_61 <= io_A_Valid_1_delay_1_62;
    io_A_Valid_1_delay_3_60 <= io_A_Valid_1_delay_2_61;
    io_A_Valid_1_delay_4_59 <= io_A_Valid_1_delay_3_60;
    io_A_Valid_1_delay_5_58 <= io_A_Valid_1_delay_4_59;
    io_A_Valid_1_delay_6_57 <= io_A_Valid_1_delay_5_58;
    io_A_Valid_1_delay_7_56 <= io_A_Valid_1_delay_6_57;
    io_A_Valid_1_delay_8_55 <= io_A_Valid_1_delay_7_56;
    io_A_Valid_1_delay_9_54 <= io_A_Valid_1_delay_8_55;
    io_A_Valid_1_delay_10_53 <= io_A_Valid_1_delay_9_54;
    io_A_Valid_1_delay_11_52 <= io_A_Valid_1_delay_10_53;
    io_A_Valid_1_delay_12_51 <= io_A_Valid_1_delay_11_52;
    io_A_Valid_1_delay_13_50 <= io_A_Valid_1_delay_12_51;
    io_A_Valid_1_delay_14_49 <= io_A_Valid_1_delay_13_50;
    io_A_Valid_1_delay_15_48 <= io_A_Valid_1_delay_14_49;
    io_A_Valid_1_delay_16_47 <= io_A_Valid_1_delay_15_48;
    io_A_Valid_1_delay_17_46 <= io_A_Valid_1_delay_16_47;
    io_A_Valid_1_delay_18_45 <= io_A_Valid_1_delay_17_46;
    io_A_Valid_1_delay_19_44 <= io_A_Valid_1_delay_18_45;
    io_A_Valid_1_delay_20_43 <= io_A_Valid_1_delay_19_44;
    io_A_Valid_1_delay_21_42 <= io_A_Valid_1_delay_20_43;
    io_A_Valid_1_delay_22_41 <= io_A_Valid_1_delay_21_42;
    io_A_Valid_1_delay_23_40 <= io_A_Valid_1_delay_22_41;
    io_A_Valid_1_delay_24_39 <= io_A_Valid_1_delay_23_40;
    io_A_Valid_1_delay_25_38 <= io_A_Valid_1_delay_24_39;
    io_A_Valid_1_delay_26_37 <= io_A_Valid_1_delay_25_38;
    io_A_Valid_1_delay_27_36 <= io_A_Valid_1_delay_26_37;
    io_A_Valid_1_delay_28_35 <= io_A_Valid_1_delay_27_36;
    io_A_Valid_1_delay_29_34 <= io_A_Valid_1_delay_28_35;
    io_A_Valid_1_delay_30_33 <= io_A_Valid_1_delay_29_34;
    io_A_Valid_1_delay_31_32 <= io_A_Valid_1_delay_30_33;
    io_A_Valid_1_delay_32_31 <= io_A_Valid_1_delay_31_32;
    io_A_Valid_1_delay_33_30 <= io_A_Valid_1_delay_32_31;
    io_A_Valid_1_delay_34_29 <= io_A_Valid_1_delay_33_30;
    io_A_Valid_1_delay_35_28 <= io_A_Valid_1_delay_34_29;
    io_A_Valid_1_delay_36_27 <= io_A_Valid_1_delay_35_28;
    io_A_Valid_1_delay_37_26 <= io_A_Valid_1_delay_36_27;
    io_A_Valid_1_delay_38_25 <= io_A_Valid_1_delay_37_26;
    io_A_Valid_1_delay_39_24 <= io_A_Valid_1_delay_38_25;
    io_A_Valid_1_delay_40_23 <= io_A_Valid_1_delay_39_24;
    io_A_Valid_1_delay_41_22 <= io_A_Valid_1_delay_40_23;
    io_A_Valid_1_delay_42_21 <= io_A_Valid_1_delay_41_22;
    io_A_Valid_1_delay_43_20 <= io_A_Valid_1_delay_42_21;
    io_A_Valid_1_delay_44_19 <= io_A_Valid_1_delay_43_20;
    io_A_Valid_1_delay_45_18 <= io_A_Valid_1_delay_44_19;
    io_A_Valid_1_delay_46_17 <= io_A_Valid_1_delay_45_18;
    io_A_Valid_1_delay_47_16 <= io_A_Valid_1_delay_46_17;
    io_A_Valid_1_delay_48_15 <= io_A_Valid_1_delay_47_16;
    io_A_Valid_1_delay_49_14 <= io_A_Valid_1_delay_48_15;
    io_A_Valid_1_delay_50_13 <= io_A_Valid_1_delay_49_14;
    io_A_Valid_1_delay_51_12 <= io_A_Valid_1_delay_50_13;
    io_A_Valid_1_delay_52_11 <= io_A_Valid_1_delay_51_12;
    io_A_Valid_1_delay_53_10 <= io_A_Valid_1_delay_52_11;
    io_A_Valid_1_delay_54_9 <= io_A_Valid_1_delay_53_10;
    io_A_Valid_1_delay_55_8 <= io_A_Valid_1_delay_54_9;
    io_A_Valid_1_delay_56_7 <= io_A_Valid_1_delay_55_8;
    io_A_Valid_1_delay_57_6 <= io_A_Valid_1_delay_56_7;
    io_A_Valid_1_delay_58_5 <= io_A_Valid_1_delay_57_6;
    io_A_Valid_1_delay_59_4 <= io_A_Valid_1_delay_58_5;
    io_A_Valid_1_delay_60_3 <= io_A_Valid_1_delay_59_4;
    io_A_Valid_1_delay_61_2 <= io_A_Valid_1_delay_60_3;
    io_A_Valid_1_delay_62_1 <= io_A_Valid_1_delay_61_2;
    io_A_Valid_1_delay_63 <= io_A_Valid_1_delay_62_1;
    io_B_Valid_63_delay_1 <= io_B_Valid_63;
    io_B_Valid_0_delay_1_1 <= io_B_Valid_0;
    io_B_Valid_0_delay_2 <= io_B_Valid_0_delay_1_1;
    io_A_Valid_2_delay_1 <= io_A_Valid_2;
    io_B_Valid_1_delay_1_1 <= io_B_Valid_1;
    io_B_Valid_1_delay_2 <= io_B_Valid_1_delay_1_1;
    io_A_Valid_2_delay_1_1 <= io_A_Valid_2;
    io_A_Valid_2_delay_2 <= io_A_Valid_2_delay_1_1;
    io_B_Valid_2_delay_1_1 <= io_B_Valid_2;
    io_B_Valid_2_delay_2 <= io_B_Valid_2_delay_1_1;
    io_A_Valid_2_delay_1_2 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_1 <= io_A_Valid_2_delay_1_2;
    io_A_Valid_2_delay_3 <= io_A_Valid_2_delay_2_1;
    io_B_Valid_3_delay_1_1 <= io_B_Valid_3;
    io_B_Valid_3_delay_2 <= io_B_Valid_3_delay_1_1;
    io_A_Valid_2_delay_1_3 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_2 <= io_A_Valid_2_delay_1_3;
    io_A_Valid_2_delay_3_1 <= io_A_Valid_2_delay_2_2;
    io_A_Valid_2_delay_4 <= io_A_Valid_2_delay_3_1;
    io_B_Valid_4_delay_1_1 <= io_B_Valid_4;
    io_B_Valid_4_delay_2 <= io_B_Valid_4_delay_1_1;
    io_A_Valid_2_delay_1_4 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_3 <= io_A_Valid_2_delay_1_4;
    io_A_Valid_2_delay_3_2 <= io_A_Valid_2_delay_2_3;
    io_A_Valid_2_delay_4_1 <= io_A_Valid_2_delay_3_2;
    io_A_Valid_2_delay_5 <= io_A_Valid_2_delay_4_1;
    io_B_Valid_5_delay_1_1 <= io_B_Valid_5;
    io_B_Valid_5_delay_2 <= io_B_Valid_5_delay_1_1;
    io_A_Valid_2_delay_1_5 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_4 <= io_A_Valid_2_delay_1_5;
    io_A_Valid_2_delay_3_3 <= io_A_Valid_2_delay_2_4;
    io_A_Valid_2_delay_4_2 <= io_A_Valid_2_delay_3_3;
    io_A_Valid_2_delay_5_1 <= io_A_Valid_2_delay_4_2;
    io_A_Valid_2_delay_6 <= io_A_Valid_2_delay_5_1;
    io_B_Valid_6_delay_1_1 <= io_B_Valid_6;
    io_B_Valid_6_delay_2 <= io_B_Valid_6_delay_1_1;
    io_A_Valid_2_delay_1_6 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_5 <= io_A_Valid_2_delay_1_6;
    io_A_Valid_2_delay_3_4 <= io_A_Valid_2_delay_2_5;
    io_A_Valid_2_delay_4_3 <= io_A_Valid_2_delay_3_4;
    io_A_Valid_2_delay_5_2 <= io_A_Valid_2_delay_4_3;
    io_A_Valid_2_delay_6_1 <= io_A_Valid_2_delay_5_2;
    io_A_Valid_2_delay_7 <= io_A_Valid_2_delay_6_1;
    io_B_Valid_7_delay_1_1 <= io_B_Valid_7;
    io_B_Valid_7_delay_2 <= io_B_Valid_7_delay_1_1;
    io_A_Valid_2_delay_1_7 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_6 <= io_A_Valid_2_delay_1_7;
    io_A_Valid_2_delay_3_5 <= io_A_Valid_2_delay_2_6;
    io_A_Valid_2_delay_4_4 <= io_A_Valid_2_delay_3_5;
    io_A_Valid_2_delay_5_3 <= io_A_Valid_2_delay_4_4;
    io_A_Valid_2_delay_6_2 <= io_A_Valid_2_delay_5_3;
    io_A_Valid_2_delay_7_1 <= io_A_Valid_2_delay_6_2;
    io_A_Valid_2_delay_8 <= io_A_Valid_2_delay_7_1;
    io_B_Valid_8_delay_1_1 <= io_B_Valid_8;
    io_B_Valid_8_delay_2 <= io_B_Valid_8_delay_1_1;
    io_A_Valid_2_delay_1_8 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_7 <= io_A_Valid_2_delay_1_8;
    io_A_Valid_2_delay_3_6 <= io_A_Valid_2_delay_2_7;
    io_A_Valid_2_delay_4_5 <= io_A_Valid_2_delay_3_6;
    io_A_Valid_2_delay_5_4 <= io_A_Valid_2_delay_4_5;
    io_A_Valid_2_delay_6_3 <= io_A_Valid_2_delay_5_4;
    io_A_Valid_2_delay_7_2 <= io_A_Valid_2_delay_6_3;
    io_A_Valid_2_delay_8_1 <= io_A_Valid_2_delay_7_2;
    io_A_Valid_2_delay_9 <= io_A_Valid_2_delay_8_1;
    io_B_Valid_9_delay_1_1 <= io_B_Valid_9;
    io_B_Valid_9_delay_2 <= io_B_Valid_9_delay_1_1;
    io_A_Valid_2_delay_1_9 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_8 <= io_A_Valid_2_delay_1_9;
    io_A_Valid_2_delay_3_7 <= io_A_Valid_2_delay_2_8;
    io_A_Valid_2_delay_4_6 <= io_A_Valid_2_delay_3_7;
    io_A_Valid_2_delay_5_5 <= io_A_Valid_2_delay_4_6;
    io_A_Valid_2_delay_6_4 <= io_A_Valid_2_delay_5_5;
    io_A_Valid_2_delay_7_3 <= io_A_Valid_2_delay_6_4;
    io_A_Valid_2_delay_8_2 <= io_A_Valid_2_delay_7_3;
    io_A_Valid_2_delay_9_1 <= io_A_Valid_2_delay_8_2;
    io_A_Valid_2_delay_10 <= io_A_Valid_2_delay_9_1;
    io_B_Valid_10_delay_1_1 <= io_B_Valid_10;
    io_B_Valid_10_delay_2 <= io_B_Valid_10_delay_1_1;
    io_A_Valid_2_delay_1_10 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_9 <= io_A_Valid_2_delay_1_10;
    io_A_Valid_2_delay_3_8 <= io_A_Valid_2_delay_2_9;
    io_A_Valid_2_delay_4_7 <= io_A_Valid_2_delay_3_8;
    io_A_Valid_2_delay_5_6 <= io_A_Valid_2_delay_4_7;
    io_A_Valid_2_delay_6_5 <= io_A_Valid_2_delay_5_6;
    io_A_Valid_2_delay_7_4 <= io_A_Valid_2_delay_6_5;
    io_A_Valid_2_delay_8_3 <= io_A_Valid_2_delay_7_4;
    io_A_Valid_2_delay_9_2 <= io_A_Valid_2_delay_8_3;
    io_A_Valid_2_delay_10_1 <= io_A_Valid_2_delay_9_2;
    io_A_Valid_2_delay_11 <= io_A_Valid_2_delay_10_1;
    io_B_Valid_11_delay_1_1 <= io_B_Valid_11;
    io_B_Valid_11_delay_2 <= io_B_Valid_11_delay_1_1;
    io_A_Valid_2_delay_1_11 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_10 <= io_A_Valid_2_delay_1_11;
    io_A_Valid_2_delay_3_9 <= io_A_Valid_2_delay_2_10;
    io_A_Valid_2_delay_4_8 <= io_A_Valid_2_delay_3_9;
    io_A_Valid_2_delay_5_7 <= io_A_Valid_2_delay_4_8;
    io_A_Valid_2_delay_6_6 <= io_A_Valid_2_delay_5_7;
    io_A_Valid_2_delay_7_5 <= io_A_Valid_2_delay_6_6;
    io_A_Valid_2_delay_8_4 <= io_A_Valid_2_delay_7_5;
    io_A_Valid_2_delay_9_3 <= io_A_Valid_2_delay_8_4;
    io_A_Valid_2_delay_10_2 <= io_A_Valid_2_delay_9_3;
    io_A_Valid_2_delay_11_1 <= io_A_Valid_2_delay_10_2;
    io_A_Valid_2_delay_12 <= io_A_Valid_2_delay_11_1;
    io_B_Valid_12_delay_1_1 <= io_B_Valid_12;
    io_B_Valid_12_delay_2 <= io_B_Valid_12_delay_1_1;
    io_A_Valid_2_delay_1_12 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_11 <= io_A_Valid_2_delay_1_12;
    io_A_Valid_2_delay_3_10 <= io_A_Valid_2_delay_2_11;
    io_A_Valid_2_delay_4_9 <= io_A_Valid_2_delay_3_10;
    io_A_Valid_2_delay_5_8 <= io_A_Valid_2_delay_4_9;
    io_A_Valid_2_delay_6_7 <= io_A_Valid_2_delay_5_8;
    io_A_Valid_2_delay_7_6 <= io_A_Valid_2_delay_6_7;
    io_A_Valid_2_delay_8_5 <= io_A_Valid_2_delay_7_6;
    io_A_Valid_2_delay_9_4 <= io_A_Valid_2_delay_8_5;
    io_A_Valid_2_delay_10_3 <= io_A_Valid_2_delay_9_4;
    io_A_Valid_2_delay_11_2 <= io_A_Valid_2_delay_10_3;
    io_A_Valid_2_delay_12_1 <= io_A_Valid_2_delay_11_2;
    io_A_Valid_2_delay_13 <= io_A_Valid_2_delay_12_1;
    io_B_Valid_13_delay_1_1 <= io_B_Valid_13;
    io_B_Valid_13_delay_2 <= io_B_Valid_13_delay_1_1;
    io_A_Valid_2_delay_1_13 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_12 <= io_A_Valid_2_delay_1_13;
    io_A_Valid_2_delay_3_11 <= io_A_Valid_2_delay_2_12;
    io_A_Valid_2_delay_4_10 <= io_A_Valid_2_delay_3_11;
    io_A_Valid_2_delay_5_9 <= io_A_Valid_2_delay_4_10;
    io_A_Valid_2_delay_6_8 <= io_A_Valid_2_delay_5_9;
    io_A_Valid_2_delay_7_7 <= io_A_Valid_2_delay_6_8;
    io_A_Valid_2_delay_8_6 <= io_A_Valid_2_delay_7_7;
    io_A_Valid_2_delay_9_5 <= io_A_Valid_2_delay_8_6;
    io_A_Valid_2_delay_10_4 <= io_A_Valid_2_delay_9_5;
    io_A_Valid_2_delay_11_3 <= io_A_Valid_2_delay_10_4;
    io_A_Valid_2_delay_12_2 <= io_A_Valid_2_delay_11_3;
    io_A_Valid_2_delay_13_1 <= io_A_Valid_2_delay_12_2;
    io_A_Valid_2_delay_14 <= io_A_Valid_2_delay_13_1;
    io_B_Valid_14_delay_1_1 <= io_B_Valid_14;
    io_B_Valid_14_delay_2 <= io_B_Valid_14_delay_1_1;
    io_A_Valid_2_delay_1_14 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_13 <= io_A_Valid_2_delay_1_14;
    io_A_Valid_2_delay_3_12 <= io_A_Valid_2_delay_2_13;
    io_A_Valid_2_delay_4_11 <= io_A_Valid_2_delay_3_12;
    io_A_Valid_2_delay_5_10 <= io_A_Valid_2_delay_4_11;
    io_A_Valid_2_delay_6_9 <= io_A_Valid_2_delay_5_10;
    io_A_Valid_2_delay_7_8 <= io_A_Valid_2_delay_6_9;
    io_A_Valid_2_delay_8_7 <= io_A_Valid_2_delay_7_8;
    io_A_Valid_2_delay_9_6 <= io_A_Valid_2_delay_8_7;
    io_A_Valid_2_delay_10_5 <= io_A_Valid_2_delay_9_6;
    io_A_Valid_2_delay_11_4 <= io_A_Valid_2_delay_10_5;
    io_A_Valid_2_delay_12_3 <= io_A_Valid_2_delay_11_4;
    io_A_Valid_2_delay_13_2 <= io_A_Valid_2_delay_12_3;
    io_A_Valid_2_delay_14_1 <= io_A_Valid_2_delay_13_2;
    io_A_Valid_2_delay_15 <= io_A_Valid_2_delay_14_1;
    io_B_Valid_15_delay_1_1 <= io_B_Valid_15;
    io_B_Valid_15_delay_2 <= io_B_Valid_15_delay_1_1;
    io_A_Valid_2_delay_1_15 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_14 <= io_A_Valid_2_delay_1_15;
    io_A_Valid_2_delay_3_13 <= io_A_Valid_2_delay_2_14;
    io_A_Valid_2_delay_4_12 <= io_A_Valid_2_delay_3_13;
    io_A_Valid_2_delay_5_11 <= io_A_Valid_2_delay_4_12;
    io_A_Valid_2_delay_6_10 <= io_A_Valid_2_delay_5_11;
    io_A_Valid_2_delay_7_9 <= io_A_Valid_2_delay_6_10;
    io_A_Valid_2_delay_8_8 <= io_A_Valid_2_delay_7_9;
    io_A_Valid_2_delay_9_7 <= io_A_Valid_2_delay_8_8;
    io_A_Valid_2_delay_10_6 <= io_A_Valid_2_delay_9_7;
    io_A_Valid_2_delay_11_5 <= io_A_Valid_2_delay_10_6;
    io_A_Valid_2_delay_12_4 <= io_A_Valid_2_delay_11_5;
    io_A_Valid_2_delay_13_3 <= io_A_Valid_2_delay_12_4;
    io_A_Valid_2_delay_14_2 <= io_A_Valid_2_delay_13_3;
    io_A_Valid_2_delay_15_1 <= io_A_Valid_2_delay_14_2;
    io_A_Valid_2_delay_16 <= io_A_Valid_2_delay_15_1;
    io_B_Valid_16_delay_1_1 <= io_B_Valid_16;
    io_B_Valid_16_delay_2 <= io_B_Valid_16_delay_1_1;
    io_A_Valid_2_delay_1_16 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_15 <= io_A_Valid_2_delay_1_16;
    io_A_Valid_2_delay_3_14 <= io_A_Valid_2_delay_2_15;
    io_A_Valid_2_delay_4_13 <= io_A_Valid_2_delay_3_14;
    io_A_Valid_2_delay_5_12 <= io_A_Valid_2_delay_4_13;
    io_A_Valid_2_delay_6_11 <= io_A_Valid_2_delay_5_12;
    io_A_Valid_2_delay_7_10 <= io_A_Valid_2_delay_6_11;
    io_A_Valid_2_delay_8_9 <= io_A_Valid_2_delay_7_10;
    io_A_Valid_2_delay_9_8 <= io_A_Valid_2_delay_8_9;
    io_A_Valid_2_delay_10_7 <= io_A_Valid_2_delay_9_8;
    io_A_Valid_2_delay_11_6 <= io_A_Valid_2_delay_10_7;
    io_A_Valid_2_delay_12_5 <= io_A_Valid_2_delay_11_6;
    io_A_Valid_2_delay_13_4 <= io_A_Valid_2_delay_12_5;
    io_A_Valid_2_delay_14_3 <= io_A_Valid_2_delay_13_4;
    io_A_Valid_2_delay_15_2 <= io_A_Valid_2_delay_14_3;
    io_A_Valid_2_delay_16_1 <= io_A_Valid_2_delay_15_2;
    io_A_Valid_2_delay_17 <= io_A_Valid_2_delay_16_1;
    io_B_Valid_17_delay_1_1 <= io_B_Valid_17;
    io_B_Valid_17_delay_2 <= io_B_Valid_17_delay_1_1;
    io_A_Valid_2_delay_1_17 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_16 <= io_A_Valid_2_delay_1_17;
    io_A_Valid_2_delay_3_15 <= io_A_Valid_2_delay_2_16;
    io_A_Valid_2_delay_4_14 <= io_A_Valid_2_delay_3_15;
    io_A_Valid_2_delay_5_13 <= io_A_Valid_2_delay_4_14;
    io_A_Valid_2_delay_6_12 <= io_A_Valid_2_delay_5_13;
    io_A_Valid_2_delay_7_11 <= io_A_Valid_2_delay_6_12;
    io_A_Valid_2_delay_8_10 <= io_A_Valid_2_delay_7_11;
    io_A_Valid_2_delay_9_9 <= io_A_Valid_2_delay_8_10;
    io_A_Valid_2_delay_10_8 <= io_A_Valid_2_delay_9_9;
    io_A_Valid_2_delay_11_7 <= io_A_Valid_2_delay_10_8;
    io_A_Valid_2_delay_12_6 <= io_A_Valid_2_delay_11_7;
    io_A_Valid_2_delay_13_5 <= io_A_Valid_2_delay_12_6;
    io_A_Valid_2_delay_14_4 <= io_A_Valid_2_delay_13_5;
    io_A_Valid_2_delay_15_3 <= io_A_Valid_2_delay_14_4;
    io_A_Valid_2_delay_16_2 <= io_A_Valid_2_delay_15_3;
    io_A_Valid_2_delay_17_1 <= io_A_Valid_2_delay_16_2;
    io_A_Valid_2_delay_18 <= io_A_Valid_2_delay_17_1;
    io_B_Valid_18_delay_1_1 <= io_B_Valid_18;
    io_B_Valid_18_delay_2 <= io_B_Valid_18_delay_1_1;
    io_A_Valid_2_delay_1_18 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_17 <= io_A_Valid_2_delay_1_18;
    io_A_Valid_2_delay_3_16 <= io_A_Valid_2_delay_2_17;
    io_A_Valid_2_delay_4_15 <= io_A_Valid_2_delay_3_16;
    io_A_Valid_2_delay_5_14 <= io_A_Valid_2_delay_4_15;
    io_A_Valid_2_delay_6_13 <= io_A_Valid_2_delay_5_14;
    io_A_Valid_2_delay_7_12 <= io_A_Valid_2_delay_6_13;
    io_A_Valid_2_delay_8_11 <= io_A_Valid_2_delay_7_12;
    io_A_Valid_2_delay_9_10 <= io_A_Valid_2_delay_8_11;
    io_A_Valid_2_delay_10_9 <= io_A_Valid_2_delay_9_10;
    io_A_Valid_2_delay_11_8 <= io_A_Valid_2_delay_10_9;
    io_A_Valid_2_delay_12_7 <= io_A_Valid_2_delay_11_8;
    io_A_Valid_2_delay_13_6 <= io_A_Valid_2_delay_12_7;
    io_A_Valid_2_delay_14_5 <= io_A_Valid_2_delay_13_6;
    io_A_Valid_2_delay_15_4 <= io_A_Valid_2_delay_14_5;
    io_A_Valid_2_delay_16_3 <= io_A_Valid_2_delay_15_4;
    io_A_Valid_2_delay_17_2 <= io_A_Valid_2_delay_16_3;
    io_A_Valid_2_delay_18_1 <= io_A_Valid_2_delay_17_2;
    io_A_Valid_2_delay_19 <= io_A_Valid_2_delay_18_1;
    io_B_Valid_19_delay_1_1 <= io_B_Valid_19;
    io_B_Valid_19_delay_2 <= io_B_Valid_19_delay_1_1;
    io_A_Valid_2_delay_1_19 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_18 <= io_A_Valid_2_delay_1_19;
    io_A_Valid_2_delay_3_17 <= io_A_Valid_2_delay_2_18;
    io_A_Valid_2_delay_4_16 <= io_A_Valid_2_delay_3_17;
    io_A_Valid_2_delay_5_15 <= io_A_Valid_2_delay_4_16;
    io_A_Valid_2_delay_6_14 <= io_A_Valid_2_delay_5_15;
    io_A_Valid_2_delay_7_13 <= io_A_Valid_2_delay_6_14;
    io_A_Valid_2_delay_8_12 <= io_A_Valid_2_delay_7_13;
    io_A_Valid_2_delay_9_11 <= io_A_Valid_2_delay_8_12;
    io_A_Valid_2_delay_10_10 <= io_A_Valid_2_delay_9_11;
    io_A_Valid_2_delay_11_9 <= io_A_Valid_2_delay_10_10;
    io_A_Valid_2_delay_12_8 <= io_A_Valid_2_delay_11_9;
    io_A_Valid_2_delay_13_7 <= io_A_Valid_2_delay_12_8;
    io_A_Valid_2_delay_14_6 <= io_A_Valid_2_delay_13_7;
    io_A_Valid_2_delay_15_5 <= io_A_Valid_2_delay_14_6;
    io_A_Valid_2_delay_16_4 <= io_A_Valid_2_delay_15_5;
    io_A_Valid_2_delay_17_3 <= io_A_Valid_2_delay_16_4;
    io_A_Valid_2_delay_18_2 <= io_A_Valid_2_delay_17_3;
    io_A_Valid_2_delay_19_1 <= io_A_Valid_2_delay_18_2;
    io_A_Valid_2_delay_20 <= io_A_Valid_2_delay_19_1;
    io_B_Valid_20_delay_1_1 <= io_B_Valid_20;
    io_B_Valid_20_delay_2 <= io_B_Valid_20_delay_1_1;
    io_A_Valid_2_delay_1_20 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_19 <= io_A_Valid_2_delay_1_20;
    io_A_Valid_2_delay_3_18 <= io_A_Valid_2_delay_2_19;
    io_A_Valid_2_delay_4_17 <= io_A_Valid_2_delay_3_18;
    io_A_Valid_2_delay_5_16 <= io_A_Valid_2_delay_4_17;
    io_A_Valid_2_delay_6_15 <= io_A_Valid_2_delay_5_16;
    io_A_Valid_2_delay_7_14 <= io_A_Valid_2_delay_6_15;
    io_A_Valid_2_delay_8_13 <= io_A_Valid_2_delay_7_14;
    io_A_Valid_2_delay_9_12 <= io_A_Valid_2_delay_8_13;
    io_A_Valid_2_delay_10_11 <= io_A_Valid_2_delay_9_12;
    io_A_Valid_2_delay_11_10 <= io_A_Valid_2_delay_10_11;
    io_A_Valid_2_delay_12_9 <= io_A_Valid_2_delay_11_10;
    io_A_Valid_2_delay_13_8 <= io_A_Valid_2_delay_12_9;
    io_A_Valid_2_delay_14_7 <= io_A_Valid_2_delay_13_8;
    io_A_Valid_2_delay_15_6 <= io_A_Valid_2_delay_14_7;
    io_A_Valid_2_delay_16_5 <= io_A_Valid_2_delay_15_6;
    io_A_Valid_2_delay_17_4 <= io_A_Valid_2_delay_16_5;
    io_A_Valid_2_delay_18_3 <= io_A_Valid_2_delay_17_4;
    io_A_Valid_2_delay_19_2 <= io_A_Valid_2_delay_18_3;
    io_A_Valid_2_delay_20_1 <= io_A_Valid_2_delay_19_2;
    io_A_Valid_2_delay_21 <= io_A_Valid_2_delay_20_1;
    io_B_Valid_21_delay_1_1 <= io_B_Valid_21;
    io_B_Valid_21_delay_2 <= io_B_Valid_21_delay_1_1;
    io_A_Valid_2_delay_1_21 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_20 <= io_A_Valid_2_delay_1_21;
    io_A_Valid_2_delay_3_19 <= io_A_Valid_2_delay_2_20;
    io_A_Valid_2_delay_4_18 <= io_A_Valid_2_delay_3_19;
    io_A_Valid_2_delay_5_17 <= io_A_Valid_2_delay_4_18;
    io_A_Valid_2_delay_6_16 <= io_A_Valid_2_delay_5_17;
    io_A_Valid_2_delay_7_15 <= io_A_Valid_2_delay_6_16;
    io_A_Valid_2_delay_8_14 <= io_A_Valid_2_delay_7_15;
    io_A_Valid_2_delay_9_13 <= io_A_Valid_2_delay_8_14;
    io_A_Valid_2_delay_10_12 <= io_A_Valid_2_delay_9_13;
    io_A_Valid_2_delay_11_11 <= io_A_Valid_2_delay_10_12;
    io_A_Valid_2_delay_12_10 <= io_A_Valid_2_delay_11_11;
    io_A_Valid_2_delay_13_9 <= io_A_Valid_2_delay_12_10;
    io_A_Valid_2_delay_14_8 <= io_A_Valid_2_delay_13_9;
    io_A_Valid_2_delay_15_7 <= io_A_Valid_2_delay_14_8;
    io_A_Valid_2_delay_16_6 <= io_A_Valid_2_delay_15_7;
    io_A_Valid_2_delay_17_5 <= io_A_Valid_2_delay_16_6;
    io_A_Valid_2_delay_18_4 <= io_A_Valid_2_delay_17_5;
    io_A_Valid_2_delay_19_3 <= io_A_Valid_2_delay_18_4;
    io_A_Valid_2_delay_20_2 <= io_A_Valid_2_delay_19_3;
    io_A_Valid_2_delay_21_1 <= io_A_Valid_2_delay_20_2;
    io_A_Valid_2_delay_22 <= io_A_Valid_2_delay_21_1;
    io_B_Valid_22_delay_1_1 <= io_B_Valid_22;
    io_B_Valid_22_delay_2 <= io_B_Valid_22_delay_1_1;
    io_A_Valid_2_delay_1_22 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_21 <= io_A_Valid_2_delay_1_22;
    io_A_Valid_2_delay_3_20 <= io_A_Valid_2_delay_2_21;
    io_A_Valid_2_delay_4_19 <= io_A_Valid_2_delay_3_20;
    io_A_Valid_2_delay_5_18 <= io_A_Valid_2_delay_4_19;
    io_A_Valid_2_delay_6_17 <= io_A_Valid_2_delay_5_18;
    io_A_Valid_2_delay_7_16 <= io_A_Valid_2_delay_6_17;
    io_A_Valid_2_delay_8_15 <= io_A_Valid_2_delay_7_16;
    io_A_Valid_2_delay_9_14 <= io_A_Valid_2_delay_8_15;
    io_A_Valid_2_delay_10_13 <= io_A_Valid_2_delay_9_14;
    io_A_Valid_2_delay_11_12 <= io_A_Valid_2_delay_10_13;
    io_A_Valid_2_delay_12_11 <= io_A_Valid_2_delay_11_12;
    io_A_Valid_2_delay_13_10 <= io_A_Valid_2_delay_12_11;
    io_A_Valid_2_delay_14_9 <= io_A_Valid_2_delay_13_10;
    io_A_Valid_2_delay_15_8 <= io_A_Valid_2_delay_14_9;
    io_A_Valid_2_delay_16_7 <= io_A_Valid_2_delay_15_8;
    io_A_Valid_2_delay_17_6 <= io_A_Valid_2_delay_16_7;
    io_A_Valid_2_delay_18_5 <= io_A_Valid_2_delay_17_6;
    io_A_Valid_2_delay_19_4 <= io_A_Valid_2_delay_18_5;
    io_A_Valid_2_delay_20_3 <= io_A_Valid_2_delay_19_4;
    io_A_Valid_2_delay_21_2 <= io_A_Valid_2_delay_20_3;
    io_A_Valid_2_delay_22_1 <= io_A_Valid_2_delay_21_2;
    io_A_Valid_2_delay_23 <= io_A_Valid_2_delay_22_1;
    io_B_Valid_23_delay_1_1 <= io_B_Valid_23;
    io_B_Valid_23_delay_2 <= io_B_Valid_23_delay_1_1;
    io_A_Valid_2_delay_1_23 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_22 <= io_A_Valid_2_delay_1_23;
    io_A_Valid_2_delay_3_21 <= io_A_Valid_2_delay_2_22;
    io_A_Valid_2_delay_4_20 <= io_A_Valid_2_delay_3_21;
    io_A_Valid_2_delay_5_19 <= io_A_Valid_2_delay_4_20;
    io_A_Valid_2_delay_6_18 <= io_A_Valid_2_delay_5_19;
    io_A_Valid_2_delay_7_17 <= io_A_Valid_2_delay_6_18;
    io_A_Valid_2_delay_8_16 <= io_A_Valid_2_delay_7_17;
    io_A_Valid_2_delay_9_15 <= io_A_Valid_2_delay_8_16;
    io_A_Valid_2_delay_10_14 <= io_A_Valid_2_delay_9_15;
    io_A_Valid_2_delay_11_13 <= io_A_Valid_2_delay_10_14;
    io_A_Valid_2_delay_12_12 <= io_A_Valid_2_delay_11_13;
    io_A_Valid_2_delay_13_11 <= io_A_Valid_2_delay_12_12;
    io_A_Valid_2_delay_14_10 <= io_A_Valid_2_delay_13_11;
    io_A_Valid_2_delay_15_9 <= io_A_Valid_2_delay_14_10;
    io_A_Valid_2_delay_16_8 <= io_A_Valid_2_delay_15_9;
    io_A_Valid_2_delay_17_7 <= io_A_Valid_2_delay_16_8;
    io_A_Valid_2_delay_18_6 <= io_A_Valid_2_delay_17_7;
    io_A_Valid_2_delay_19_5 <= io_A_Valid_2_delay_18_6;
    io_A_Valid_2_delay_20_4 <= io_A_Valid_2_delay_19_5;
    io_A_Valid_2_delay_21_3 <= io_A_Valid_2_delay_20_4;
    io_A_Valid_2_delay_22_2 <= io_A_Valid_2_delay_21_3;
    io_A_Valid_2_delay_23_1 <= io_A_Valid_2_delay_22_2;
    io_A_Valid_2_delay_24 <= io_A_Valid_2_delay_23_1;
    io_B_Valid_24_delay_1_1 <= io_B_Valid_24;
    io_B_Valid_24_delay_2 <= io_B_Valid_24_delay_1_1;
    io_A_Valid_2_delay_1_24 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_23 <= io_A_Valid_2_delay_1_24;
    io_A_Valid_2_delay_3_22 <= io_A_Valid_2_delay_2_23;
    io_A_Valid_2_delay_4_21 <= io_A_Valid_2_delay_3_22;
    io_A_Valid_2_delay_5_20 <= io_A_Valid_2_delay_4_21;
    io_A_Valid_2_delay_6_19 <= io_A_Valid_2_delay_5_20;
    io_A_Valid_2_delay_7_18 <= io_A_Valid_2_delay_6_19;
    io_A_Valid_2_delay_8_17 <= io_A_Valid_2_delay_7_18;
    io_A_Valid_2_delay_9_16 <= io_A_Valid_2_delay_8_17;
    io_A_Valid_2_delay_10_15 <= io_A_Valid_2_delay_9_16;
    io_A_Valid_2_delay_11_14 <= io_A_Valid_2_delay_10_15;
    io_A_Valid_2_delay_12_13 <= io_A_Valid_2_delay_11_14;
    io_A_Valid_2_delay_13_12 <= io_A_Valid_2_delay_12_13;
    io_A_Valid_2_delay_14_11 <= io_A_Valid_2_delay_13_12;
    io_A_Valid_2_delay_15_10 <= io_A_Valid_2_delay_14_11;
    io_A_Valid_2_delay_16_9 <= io_A_Valid_2_delay_15_10;
    io_A_Valid_2_delay_17_8 <= io_A_Valid_2_delay_16_9;
    io_A_Valid_2_delay_18_7 <= io_A_Valid_2_delay_17_8;
    io_A_Valid_2_delay_19_6 <= io_A_Valid_2_delay_18_7;
    io_A_Valid_2_delay_20_5 <= io_A_Valid_2_delay_19_6;
    io_A_Valid_2_delay_21_4 <= io_A_Valid_2_delay_20_5;
    io_A_Valid_2_delay_22_3 <= io_A_Valid_2_delay_21_4;
    io_A_Valid_2_delay_23_2 <= io_A_Valid_2_delay_22_3;
    io_A_Valid_2_delay_24_1 <= io_A_Valid_2_delay_23_2;
    io_A_Valid_2_delay_25 <= io_A_Valid_2_delay_24_1;
    io_B_Valid_25_delay_1_1 <= io_B_Valid_25;
    io_B_Valid_25_delay_2 <= io_B_Valid_25_delay_1_1;
    io_A_Valid_2_delay_1_25 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_24 <= io_A_Valid_2_delay_1_25;
    io_A_Valid_2_delay_3_23 <= io_A_Valid_2_delay_2_24;
    io_A_Valid_2_delay_4_22 <= io_A_Valid_2_delay_3_23;
    io_A_Valid_2_delay_5_21 <= io_A_Valid_2_delay_4_22;
    io_A_Valid_2_delay_6_20 <= io_A_Valid_2_delay_5_21;
    io_A_Valid_2_delay_7_19 <= io_A_Valid_2_delay_6_20;
    io_A_Valid_2_delay_8_18 <= io_A_Valid_2_delay_7_19;
    io_A_Valid_2_delay_9_17 <= io_A_Valid_2_delay_8_18;
    io_A_Valid_2_delay_10_16 <= io_A_Valid_2_delay_9_17;
    io_A_Valid_2_delay_11_15 <= io_A_Valid_2_delay_10_16;
    io_A_Valid_2_delay_12_14 <= io_A_Valid_2_delay_11_15;
    io_A_Valid_2_delay_13_13 <= io_A_Valid_2_delay_12_14;
    io_A_Valid_2_delay_14_12 <= io_A_Valid_2_delay_13_13;
    io_A_Valid_2_delay_15_11 <= io_A_Valid_2_delay_14_12;
    io_A_Valid_2_delay_16_10 <= io_A_Valid_2_delay_15_11;
    io_A_Valid_2_delay_17_9 <= io_A_Valid_2_delay_16_10;
    io_A_Valid_2_delay_18_8 <= io_A_Valid_2_delay_17_9;
    io_A_Valid_2_delay_19_7 <= io_A_Valid_2_delay_18_8;
    io_A_Valid_2_delay_20_6 <= io_A_Valid_2_delay_19_7;
    io_A_Valid_2_delay_21_5 <= io_A_Valid_2_delay_20_6;
    io_A_Valid_2_delay_22_4 <= io_A_Valid_2_delay_21_5;
    io_A_Valid_2_delay_23_3 <= io_A_Valid_2_delay_22_4;
    io_A_Valid_2_delay_24_2 <= io_A_Valid_2_delay_23_3;
    io_A_Valid_2_delay_25_1 <= io_A_Valid_2_delay_24_2;
    io_A_Valid_2_delay_26 <= io_A_Valid_2_delay_25_1;
    io_B_Valid_26_delay_1_1 <= io_B_Valid_26;
    io_B_Valid_26_delay_2 <= io_B_Valid_26_delay_1_1;
    io_A_Valid_2_delay_1_26 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_25 <= io_A_Valid_2_delay_1_26;
    io_A_Valid_2_delay_3_24 <= io_A_Valid_2_delay_2_25;
    io_A_Valid_2_delay_4_23 <= io_A_Valid_2_delay_3_24;
    io_A_Valid_2_delay_5_22 <= io_A_Valid_2_delay_4_23;
    io_A_Valid_2_delay_6_21 <= io_A_Valid_2_delay_5_22;
    io_A_Valid_2_delay_7_20 <= io_A_Valid_2_delay_6_21;
    io_A_Valid_2_delay_8_19 <= io_A_Valid_2_delay_7_20;
    io_A_Valid_2_delay_9_18 <= io_A_Valid_2_delay_8_19;
    io_A_Valid_2_delay_10_17 <= io_A_Valid_2_delay_9_18;
    io_A_Valid_2_delay_11_16 <= io_A_Valid_2_delay_10_17;
    io_A_Valid_2_delay_12_15 <= io_A_Valid_2_delay_11_16;
    io_A_Valid_2_delay_13_14 <= io_A_Valid_2_delay_12_15;
    io_A_Valid_2_delay_14_13 <= io_A_Valid_2_delay_13_14;
    io_A_Valid_2_delay_15_12 <= io_A_Valid_2_delay_14_13;
    io_A_Valid_2_delay_16_11 <= io_A_Valid_2_delay_15_12;
    io_A_Valid_2_delay_17_10 <= io_A_Valid_2_delay_16_11;
    io_A_Valid_2_delay_18_9 <= io_A_Valid_2_delay_17_10;
    io_A_Valid_2_delay_19_8 <= io_A_Valid_2_delay_18_9;
    io_A_Valid_2_delay_20_7 <= io_A_Valid_2_delay_19_8;
    io_A_Valid_2_delay_21_6 <= io_A_Valid_2_delay_20_7;
    io_A_Valid_2_delay_22_5 <= io_A_Valid_2_delay_21_6;
    io_A_Valid_2_delay_23_4 <= io_A_Valid_2_delay_22_5;
    io_A_Valid_2_delay_24_3 <= io_A_Valid_2_delay_23_4;
    io_A_Valid_2_delay_25_2 <= io_A_Valid_2_delay_24_3;
    io_A_Valid_2_delay_26_1 <= io_A_Valid_2_delay_25_2;
    io_A_Valid_2_delay_27 <= io_A_Valid_2_delay_26_1;
    io_B_Valid_27_delay_1_1 <= io_B_Valid_27;
    io_B_Valid_27_delay_2 <= io_B_Valid_27_delay_1_1;
    io_A_Valid_2_delay_1_27 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_26 <= io_A_Valid_2_delay_1_27;
    io_A_Valid_2_delay_3_25 <= io_A_Valid_2_delay_2_26;
    io_A_Valid_2_delay_4_24 <= io_A_Valid_2_delay_3_25;
    io_A_Valid_2_delay_5_23 <= io_A_Valid_2_delay_4_24;
    io_A_Valid_2_delay_6_22 <= io_A_Valid_2_delay_5_23;
    io_A_Valid_2_delay_7_21 <= io_A_Valid_2_delay_6_22;
    io_A_Valid_2_delay_8_20 <= io_A_Valid_2_delay_7_21;
    io_A_Valid_2_delay_9_19 <= io_A_Valid_2_delay_8_20;
    io_A_Valid_2_delay_10_18 <= io_A_Valid_2_delay_9_19;
    io_A_Valid_2_delay_11_17 <= io_A_Valid_2_delay_10_18;
    io_A_Valid_2_delay_12_16 <= io_A_Valid_2_delay_11_17;
    io_A_Valid_2_delay_13_15 <= io_A_Valid_2_delay_12_16;
    io_A_Valid_2_delay_14_14 <= io_A_Valid_2_delay_13_15;
    io_A_Valid_2_delay_15_13 <= io_A_Valid_2_delay_14_14;
    io_A_Valid_2_delay_16_12 <= io_A_Valid_2_delay_15_13;
    io_A_Valid_2_delay_17_11 <= io_A_Valid_2_delay_16_12;
    io_A_Valid_2_delay_18_10 <= io_A_Valid_2_delay_17_11;
    io_A_Valid_2_delay_19_9 <= io_A_Valid_2_delay_18_10;
    io_A_Valid_2_delay_20_8 <= io_A_Valid_2_delay_19_9;
    io_A_Valid_2_delay_21_7 <= io_A_Valid_2_delay_20_8;
    io_A_Valid_2_delay_22_6 <= io_A_Valid_2_delay_21_7;
    io_A_Valid_2_delay_23_5 <= io_A_Valid_2_delay_22_6;
    io_A_Valid_2_delay_24_4 <= io_A_Valid_2_delay_23_5;
    io_A_Valid_2_delay_25_3 <= io_A_Valid_2_delay_24_4;
    io_A_Valid_2_delay_26_2 <= io_A_Valid_2_delay_25_3;
    io_A_Valid_2_delay_27_1 <= io_A_Valid_2_delay_26_2;
    io_A_Valid_2_delay_28 <= io_A_Valid_2_delay_27_1;
    io_B_Valid_28_delay_1_1 <= io_B_Valid_28;
    io_B_Valid_28_delay_2 <= io_B_Valid_28_delay_1_1;
    io_A_Valid_2_delay_1_28 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_27 <= io_A_Valid_2_delay_1_28;
    io_A_Valid_2_delay_3_26 <= io_A_Valid_2_delay_2_27;
    io_A_Valid_2_delay_4_25 <= io_A_Valid_2_delay_3_26;
    io_A_Valid_2_delay_5_24 <= io_A_Valid_2_delay_4_25;
    io_A_Valid_2_delay_6_23 <= io_A_Valid_2_delay_5_24;
    io_A_Valid_2_delay_7_22 <= io_A_Valid_2_delay_6_23;
    io_A_Valid_2_delay_8_21 <= io_A_Valid_2_delay_7_22;
    io_A_Valid_2_delay_9_20 <= io_A_Valid_2_delay_8_21;
    io_A_Valid_2_delay_10_19 <= io_A_Valid_2_delay_9_20;
    io_A_Valid_2_delay_11_18 <= io_A_Valid_2_delay_10_19;
    io_A_Valid_2_delay_12_17 <= io_A_Valid_2_delay_11_18;
    io_A_Valid_2_delay_13_16 <= io_A_Valid_2_delay_12_17;
    io_A_Valid_2_delay_14_15 <= io_A_Valid_2_delay_13_16;
    io_A_Valid_2_delay_15_14 <= io_A_Valid_2_delay_14_15;
    io_A_Valid_2_delay_16_13 <= io_A_Valid_2_delay_15_14;
    io_A_Valid_2_delay_17_12 <= io_A_Valid_2_delay_16_13;
    io_A_Valid_2_delay_18_11 <= io_A_Valid_2_delay_17_12;
    io_A_Valid_2_delay_19_10 <= io_A_Valid_2_delay_18_11;
    io_A_Valid_2_delay_20_9 <= io_A_Valid_2_delay_19_10;
    io_A_Valid_2_delay_21_8 <= io_A_Valid_2_delay_20_9;
    io_A_Valid_2_delay_22_7 <= io_A_Valid_2_delay_21_8;
    io_A_Valid_2_delay_23_6 <= io_A_Valid_2_delay_22_7;
    io_A_Valid_2_delay_24_5 <= io_A_Valid_2_delay_23_6;
    io_A_Valid_2_delay_25_4 <= io_A_Valid_2_delay_24_5;
    io_A_Valid_2_delay_26_3 <= io_A_Valid_2_delay_25_4;
    io_A_Valid_2_delay_27_2 <= io_A_Valid_2_delay_26_3;
    io_A_Valid_2_delay_28_1 <= io_A_Valid_2_delay_27_2;
    io_A_Valid_2_delay_29 <= io_A_Valid_2_delay_28_1;
    io_B_Valid_29_delay_1_1 <= io_B_Valid_29;
    io_B_Valid_29_delay_2 <= io_B_Valid_29_delay_1_1;
    io_A_Valid_2_delay_1_29 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_28 <= io_A_Valid_2_delay_1_29;
    io_A_Valid_2_delay_3_27 <= io_A_Valid_2_delay_2_28;
    io_A_Valid_2_delay_4_26 <= io_A_Valid_2_delay_3_27;
    io_A_Valid_2_delay_5_25 <= io_A_Valid_2_delay_4_26;
    io_A_Valid_2_delay_6_24 <= io_A_Valid_2_delay_5_25;
    io_A_Valid_2_delay_7_23 <= io_A_Valid_2_delay_6_24;
    io_A_Valid_2_delay_8_22 <= io_A_Valid_2_delay_7_23;
    io_A_Valid_2_delay_9_21 <= io_A_Valid_2_delay_8_22;
    io_A_Valid_2_delay_10_20 <= io_A_Valid_2_delay_9_21;
    io_A_Valid_2_delay_11_19 <= io_A_Valid_2_delay_10_20;
    io_A_Valid_2_delay_12_18 <= io_A_Valid_2_delay_11_19;
    io_A_Valid_2_delay_13_17 <= io_A_Valid_2_delay_12_18;
    io_A_Valid_2_delay_14_16 <= io_A_Valid_2_delay_13_17;
    io_A_Valid_2_delay_15_15 <= io_A_Valid_2_delay_14_16;
    io_A_Valid_2_delay_16_14 <= io_A_Valid_2_delay_15_15;
    io_A_Valid_2_delay_17_13 <= io_A_Valid_2_delay_16_14;
    io_A_Valid_2_delay_18_12 <= io_A_Valid_2_delay_17_13;
    io_A_Valid_2_delay_19_11 <= io_A_Valid_2_delay_18_12;
    io_A_Valid_2_delay_20_10 <= io_A_Valid_2_delay_19_11;
    io_A_Valid_2_delay_21_9 <= io_A_Valid_2_delay_20_10;
    io_A_Valid_2_delay_22_8 <= io_A_Valid_2_delay_21_9;
    io_A_Valid_2_delay_23_7 <= io_A_Valid_2_delay_22_8;
    io_A_Valid_2_delay_24_6 <= io_A_Valid_2_delay_23_7;
    io_A_Valid_2_delay_25_5 <= io_A_Valid_2_delay_24_6;
    io_A_Valid_2_delay_26_4 <= io_A_Valid_2_delay_25_5;
    io_A_Valid_2_delay_27_3 <= io_A_Valid_2_delay_26_4;
    io_A_Valid_2_delay_28_2 <= io_A_Valid_2_delay_27_3;
    io_A_Valid_2_delay_29_1 <= io_A_Valid_2_delay_28_2;
    io_A_Valid_2_delay_30 <= io_A_Valid_2_delay_29_1;
    io_B_Valid_30_delay_1_1 <= io_B_Valid_30;
    io_B_Valid_30_delay_2 <= io_B_Valid_30_delay_1_1;
    io_A_Valid_2_delay_1_30 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_29 <= io_A_Valid_2_delay_1_30;
    io_A_Valid_2_delay_3_28 <= io_A_Valid_2_delay_2_29;
    io_A_Valid_2_delay_4_27 <= io_A_Valid_2_delay_3_28;
    io_A_Valid_2_delay_5_26 <= io_A_Valid_2_delay_4_27;
    io_A_Valid_2_delay_6_25 <= io_A_Valid_2_delay_5_26;
    io_A_Valid_2_delay_7_24 <= io_A_Valid_2_delay_6_25;
    io_A_Valid_2_delay_8_23 <= io_A_Valid_2_delay_7_24;
    io_A_Valid_2_delay_9_22 <= io_A_Valid_2_delay_8_23;
    io_A_Valid_2_delay_10_21 <= io_A_Valid_2_delay_9_22;
    io_A_Valid_2_delay_11_20 <= io_A_Valid_2_delay_10_21;
    io_A_Valid_2_delay_12_19 <= io_A_Valid_2_delay_11_20;
    io_A_Valid_2_delay_13_18 <= io_A_Valid_2_delay_12_19;
    io_A_Valid_2_delay_14_17 <= io_A_Valid_2_delay_13_18;
    io_A_Valid_2_delay_15_16 <= io_A_Valid_2_delay_14_17;
    io_A_Valid_2_delay_16_15 <= io_A_Valid_2_delay_15_16;
    io_A_Valid_2_delay_17_14 <= io_A_Valid_2_delay_16_15;
    io_A_Valid_2_delay_18_13 <= io_A_Valid_2_delay_17_14;
    io_A_Valid_2_delay_19_12 <= io_A_Valid_2_delay_18_13;
    io_A_Valid_2_delay_20_11 <= io_A_Valid_2_delay_19_12;
    io_A_Valid_2_delay_21_10 <= io_A_Valid_2_delay_20_11;
    io_A_Valid_2_delay_22_9 <= io_A_Valid_2_delay_21_10;
    io_A_Valid_2_delay_23_8 <= io_A_Valid_2_delay_22_9;
    io_A_Valid_2_delay_24_7 <= io_A_Valid_2_delay_23_8;
    io_A_Valid_2_delay_25_6 <= io_A_Valid_2_delay_24_7;
    io_A_Valid_2_delay_26_5 <= io_A_Valid_2_delay_25_6;
    io_A_Valid_2_delay_27_4 <= io_A_Valid_2_delay_26_5;
    io_A_Valid_2_delay_28_3 <= io_A_Valid_2_delay_27_4;
    io_A_Valid_2_delay_29_2 <= io_A_Valid_2_delay_28_3;
    io_A_Valid_2_delay_30_1 <= io_A_Valid_2_delay_29_2;
    io_A_Valid_2_delay_31 <= io_A_Valid_2_delay_30_1;
    io_B_Valid_31_delay_1_1 <= io_B_Valid_31;
    io_B_Valid_31_delay_2 <= io_B_Valid_31_delay_1_1;
    io_A_Valid_2_delay_1_31 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_30 <= io_A_Valid_2_delay_1_31;
    io_A_Valid_2_delay_3_29 <= io_A_Valid_2_delay_2_30;
    io_A_Valid_2_delay_4_28 <= io_A_Valid_2_delay_3_29;
    io_A_Valid_2_delay_5_27 <= io_A_Valid_2_delay_4_28;
    io_A_Valid_2_delay_6_26 <= io_A_Valid_2_delay_5_27;
    io_A_Valid_2_delay_7_25 <= io_A_Valid_2_delay_6_26;
    io_A_Valid_2_delay_8_24 <= io_A_Valid_2_delay_7_25;
    io_A_Valid_2_delay_9_23 <= io_A_Valid_2_delay_8_24;
    io_A_Valid_2_delay_10_22 <= io_A_Valid_2_delay_9_23;
    io_A_Valid_2_delay_11_21 <= io_A_Valid_2_delay_10_22;
    io_A_Valid_2_delay_12_20 <= io_A_Valid_2_delay_11_21;
    io_A_Valid_2_delay_13_19 <= io_A_Valid_2_delay_12_20;
    io_A_Valid_2_delay_14_18 <= io_A_Valid_2_delay_13_19;
    io_A_Valid_2_delay_15_17 <= io_A_Valid_2_delay_14_18;
    io_A_Valid_2_delay_16_16 <= io_A_Valid_2_delay_15_17;
    io_A_Valid_2_delay_17_15 <= io_A_Valid_2_delay_16_16;
    io_A_Valid_2_delay_18_14 <= io_A_Valid_2_delay_17_15;
    io_A_Valid_2_delay_19_13 <= io_A_Valid_2_delay_18_14;
    io_A_Valid_2_delay_20_12 <= io_A_Valid_2_delay_19_13;
    io_A_Valid_2_delay_21_11 <= io_A_Valid_2_delay_20_12;
    io_A_Valid_2_delay_22_10 <= io_A_Valid_2_delay_21_11;
    io_A_Valid_2_delay_23_9 <= io_A_Valid_2_delay_22_10;
    io_A_Valid_2_delay_24_8 <= io_A_Valid_2_delay_23_9;
    io_A_Valid_2_delay_25_7 <= io_A_Valid_2_delay_24_8;
    io_A_Valid_2_delay_26_6 <= io_A_Valid_2_delay_25_7;
    io_A_Valid_2_delay_27_5 <= io_A_Valid_2_delay_26_6;
    io_A_Valid_2_delay_28_4 <= io_A_Valid_2_delay_27_5;
    io_A_Valid_2_delay_29_3 <= io_A_Valid_2_delay_28_4;
    io_A_Valid_2_delay_30_2 <= io_A_Valid_2_delay_29_3;
    io_A_Valid_2_delay_31_1 <= io_A_Valid_2_delay_30_2;
    io_A_Valid_2_delay_32 <= io_A_Valid_2_delay_31_1;
    io_B_Valid_32_delay_1_1 <= io_B_Valid_32;
    io_B_Valid_32_delay_2 <= io_B_Valid_32_delay_1_1;
    io_A_Valid_2_delay_1_32 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_31 <= io_A_Valid_2_delay_1_32;
    io_A_Valid_2_delay_3_30 <= io_A_Valid_2_delay_2_31;
    io_A_Valid_2_delay_4_29 <= io_A_Valid_2_delay_3_30;
    io_A_Valid_2_delay_5_28 <= io_A_Valid_2_delay_4_29;
    io_A_Valid_2_delay_6_27 <= io_A_Valid_2_delay_5_28;
    io_A_Valid_2_delay_7_26 <= io_A_Valid_2_delay_6_27;
    io_A_Valid_2_delay_8_25 <= io_A_Valid_2_delay_7_26;
    io_A_Valid_2_delay_9_24 <= io_A_Valid_2_delay_8_25;
    io_A_Valid_2_delay_10_23 <= io_A_Valid_2_delay_9_24;
    io_A_Valid_2_delay_11_22 <= io_A_Valid_2_delay_10_23;
    io_A_Valid_2_delay_12_21 <= io_A_Valid_2_delay_11_22;
    io_A_Valid_2_delay_13_20 <= io_A_Valid_2_delay_12_21;
    io_A_Valid_2_delay_14_19 <= io_A_Valid_2_delay_13_20;
    io_A_Valid_2_delay_15_18 <= io_A_Valid_2_delay_14_19;
    io_A_Valid_2_delay_16_17 <= io_A_Valid_2_delay_15_18;
    io_A_Valid_2_delay_17_16 <= io_A_Valid_2_delay_16_17;
    io_A_Valid_2_delay_18_15 <= io_A_Valid_2_delay_17_16;
    io_A_Valid_2_delay_19_14 <= io_A_Valid_2_delay_18_15;
    io_A_Valid_2_delay_20_13 <= io_A_Valid_2_delay_19_14;
    io_A_Valid_2_delay_21_12 <= io_A_Valid_2_delay_20_13;
    io_A_Valid_2_delay_22_11 <= io_A_Valid_2_delay_21_12;
    io_A_Valid_2_delay_23_10 <= io_A_Valid_2_delay_22_11;
    io_A_Valid_2_delay_24_9 <= io_A_Valid_2_delay_23_10;
    io_A_Valid_2_delay_25_8 <= io_A_Valid_2_delay_24_9;
    io_A_Valid_2_delay_26_7 <= io_A_Valid_2_delay_25_8;
    io_A_Valid_2_delay_27_6 <= io_A_Valid_2_delay_26_7;
    io_A_Valid_2_delay_28_5 <= io_A_Valid_2_delay_27_6;
    io_A_Valid_2_delay_29_4 <= io_A_Valid_2_delay_28_5;
    io_A_Valid_2_delay_30_3 <= io_A_Valid_2_delay_29_4;
    io_A_Valid_2_delay_31_2 <= io_A_Valid_2_delay_30_3;
    io_A_Valid_2_delay_32_1 <= io_A_Valid_2_delay_31_2;
    io_A_Valid_2_delay_33 <= io_A_Valid_2_delay_32_1;
    io_B_Valid_33_delay_1_1 <= io_B_Valid_33;
    io_B_Valid_33_delay_2 <= io_B_Valid_33_delay_1_1;
    io_A_Valid_2_delay_1_33 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_32 <= io_A_Valid_2_delay_1_33;
    io_A_Valid_2_delay_3_31 <= io_A_Valid_2_delay_2_32;
    io_A_Valid_2_delay_4_30 <= io_A_Valid_2_delay_3_31;
    io_A_Valid_2_delay_5_29 <= io_A_Valid_2_delay_4_30;
    io_A_Valid_2_delay_6_28 <= io_A_Valid_2_delay_5_29;
    io_A_Valid_2_delay_7_27 <= io_A_Valid_2_delay_6_28;
    io_A_Valid_2_delay_8_26 <= io_A_Valid_2_delay_7_27;
    io_A_Valid_2_delay_9_25 <= io_A_Valid_2_delay_8_26;
    io_A_Valid_2_delay_10_24 <= io_A_Valid_2_delay_9_25;
    io_A_Valid_2_delay_11_23 <= io_A_Valid_2_delay_10_24;
    io_A_Valid_2_delay_12_22 <= io_A_Valid_2_delay_11_23;
    io_A_Valid_2_delay_13_21 <= io_A_Valid_2_delay_12_22;
    io_A_Valid_2_delay_14_20 <= io_A_Valid_2_delay_13_21;
    io_A_Valid_2_delay_15_19 <= io_A_Valid_2_delay_14_20;
    io_A_Valid_2_delay_16_18 <= io_A_Valid_2_delay_15_19;
    io_A_Valid_2_delay_17_17 <= io_A_Valid_2_delay_16_18;
    io_A_Valid_2_delay_18_16 <= io_A_Valid_2_delay_17_17;
    io_A_Valid_2_delay_19_15 <= io_A_Valid_2_delay_18_16;
    io_A_Valid_2_delay_20_14 <= io_A_Valid_2_delay_19_15;
    io_A_Valid_2_delay_21_13 <= io_A_Valid_2_delay_20_14;
    io_A_Valid_2_delay_22_12 <= io_A_Valid_2_delay_21_13;
    io_A_Valid_2_delay_23_11 <= io_A_Valid_2_delay_22_12;
    io_A_Valid_2_delay_24_10 <= io_A_Valid_2_delay_23_11;
    io_A_Valid_2_delay_25_9 <= io_A_Valid_2_delay_24_10;
    io_A_Valid_2_delay_26_8 <= io_A_Valid_2_delay_25_9;
    io_A_Valid_2_delay_27_7 <= io_A_Valid_2_delay_26_8;
    io_A_Valid_2_delay_28_6 <= io_A_Valid_2_delay_27_7;
    io_A_Valid_2_delay_29_5 <= io_A_Valid_2_delay_28_6;
    io_A_Valid_2_delay_30_4 <= io_A_Valid_2_delay_29_5;
    io_A_Valid_2_delay_31_3 <= io_A_Valid_2_delay_30_4;
    io_A_Valid_2_delay_32_2 <= io_A_Valid_2_delay_31_3;
    io_A_Valid_2_delay_33_1 <= io_A_Valid_2_delay_32_2;
    io_A_Valid_2_delay_34 <= io_A_Valid_2_delay_33_1;
    io_B_Valid_34_delay_1_1 <= io_B_Valid_34;
    io_B_Valid_34_delay_2 <= io_B_Valid_34_delay_1_1;
    io_A_Valid_2_delay_1_34 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_33 <= io_A_Valid_2_delay_1_34;
    io_A_Valid_2_delay_3_32 <= io_A_Valid_2_delay_2_33;
    io_A_Valid_2_delay_4_31 <= io_A_Valid_2_delay_3_32;
    io_A_Valid_2_delay_5_30 <= io_A_Valid_2_delay_4_31;
    io_A_Valid_2_delay_6_29 <= io_A_Valid_2_delay_5_30;
    io_A_Valid_2_delay_7_28 <= io_A_Valid_2_delay_6_29;
    io_A_Valid_2_delay_8_27 <= io_A_Valid_2_delay_7_28;
    io_A_Valid_2_delay_9_26 <= io_A_Valid_2_delay_8_27;
    io_A_Valid_2_delay_10_25 <= io_A_Valid_2_delay_9_26;
    io_A_Valid_2_delay_11_24 <= io_A_Valid_2_delay_10_25;
    io_A_Valid_2_delay_12_23 <= io_A_Valid_2_delay_11_24;
    io_A_Valid_2_delay_13_22 <= io_A_Valid_2_delay_12_23;
    io_A_Valid_2_delay_14_21 <= io_A_Valid_2_delay_13_22;
    io_A_Valid_2_delay_15_20 <= io_A_Valid_2_delay_14_21;
    io_A_Valid_2_delay_16_19 <= io_A_Valid_2_delay_15_20;
    io_A_Valid_2_delay_17_18 <= io_A_Valid_2_delay_16_19;
    io_A_Valid_2_delay_18_17 <= io_A_Valid_2_delay_17_18;
    io_A_Valid_2_delay_19_16 <= io_A_Valid_2_delay_18_17;
    io_A_Valid_2_delay_20_15 <= io_A_Valid_2_delay_19_16;
    io_A_Valid_2_delay_21_14 <= io_A_Valid_2_delay_20_15;
    io_A_Valid_2_delay_22_13 <= io_A_Valid_2_delay_21_14;
    io_A_Valid_2_delay_23_12 <= io_A_Valid_2_delay_22_13;
    io_A_Valid_2_delay_24_11 <= io_A_Valid_2_delay_23_12;
    io_A_Valid_2_delay_25_10 <= io_A_Valid_2_delay_24_11;
    io_A_Valid_2_delay_26_9 <= io_A_Valid_2_delay_25_10;
    io_A_Valid_2_delay_27_8 <= io_A_Valid_2_delay_26_9;
    io_A_Valid_2_delay_28_7 <= io_A_Valid_2_delay_27_8;
    io_A_Valid_2_delay_29_6 <= io_A_Valid_2_delay_28_7;
    io_A_Valid_2_delay_30_5 <= io_A_Valid_2_delay_29_6;
    io_A_Valid_2_delay_31_4 <= io_A_Valid_2_delay_30_5;
    io_A_Valid_2_delay_32_3 <= io_A_Valid_2_delay_31_4;
    io_A_Valid_2_delay_33_2 <= io_A_Valid_2_delay_32_3;
    io_A_Valid_2_delay_34_1 <= io_A_Valid_2_delay_33_2;
    io_A_Valid_2_delay_35 <= io_A_Valid_2_delay_34_1;
    io_B_Valid_35_delay_1_1 <= io_B_Valid_35;
    io_B_Valid_35_delay_2 <= io_B_Valid_35_delay_1_1;
    io_A_Valid_2_delay_1_35 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_34 <= io_A_Valid_2_delay_1_35;
    io_A_Valid_2_delay_3_33 <= io_A_Valid_2_delay_2_34;
    io_A_Valid_2_delay_4_32 <= io_A_Valid_2_delay_3_33;
    io_A_Valid_2_delay_5_31 <= io_A_Valid_2_delay_4_32;
    io_A_Valid_2_delay_6_30 <= io_A_Valid_2_delay_5_31;
    io_A_Valid_2_delay_7_29 <= io_A_Valid_2_delay_6_30;
    io_A_Valid_2_delay_8_28 <= io_A_Valid_2_delay_7_29;
    io_A_Valid_2_delay_9_27 <= io_A_Valid_2_delay_8_28;
    io_A_Valid_2_delay_10_26 <= io_A_Valid_2_delay_9_27;
    io_A_Valid_2_delay_11_25 <= io_A_Valid_2_delay_10_26;
    io_A_Valid_2_delay_12_24 <= io_A_Valid_2_delay_11_25;
    io_A_Valid_2_delay_13_23 <= io_A_Valid_2_delay_12_24;
    io_A_Valid_2_delay_14_22 <= io_A_Valid_2_delay_13_23;
    io_A_Valid_2_delay_15_21 <= io_A_Valid_2_delay_14_22;
    io_A_Valid_2_delay_16_20 <= io_A_Valid_2_delay_15_21;
    io_A_Valid_2_delay_17_19 <= io_A_Valid_2_delay_16_20;
    io_A_Valid_2_delay_18_18 <= io_A_Valid_2_delay_17_19;
    io_A_Valid_2_delay_19_17 <= io_A_Valid_2_delay_18_18;
    io_A_Valid_2_delay_20_16 <= io_A_Valid_2_delay_19_17;
    io_A_Valid_2_delay_21_15 <= io_A_Valid_2_delay_20_16;
    io_A_Valid_2_delay_22_14 <= io_A_Valid_2_delay_21_15;
    io_A_Valid_2_delay_23_13 <= io_A_Valid_2_delay_22_14;
    io_A_Valid_2_delay_24_12 <= io_A_Valid_2_delay_23_13;
    io_A_Valid_2_delay_25_11 <= io_A_Valid_2_delay_24_12;
    io_A_Valid_2_delay_26_10 <= io_A_Valid_2_delay_25_11;
    io_A_Valid_2_delay_27_9 <= io_A_Valid_2_delay_26_10;
    io_A_Valid_2_delay_28_8 <= io_A_Valid_2_delay_27_9;
    io_A_Valid_2_delay_29_7 <= io_A_Valid_2_delay_28_8;
    io_A_Valid_2_delay_30_6 <= io_A_Valid_2_delay_29_7;
    io_A_Valid_2_delay_31_5 <= io_A_Valid_2_delay_30_6;
    io_A_Valid_2_delay_32_4 <= io_A_Valid_2_delay_31_5;
    io_A_Valid_2_delay_33_3 <= io_A_Valid_2_delay_32_4;
    io_A_Valid_2_delay_34_2 <= io_A_Valid_2_delay_33_3;
    io_A_Valid_2_delay_35_1 <= io_A_Valid_2_delay_34_2;
    io_A_Valid_2_delay_36 <= io_A_Valid_2_delay_35_1;
    io_B_Valid_36_delay_1_1 <= io_B_Valid_36;
    io_B_Valid_36_delay_2 <= io_B_Valid_36_delay_1_1;
    io_A_Valid_2_delay_1_36 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_35 <= io_A_Valid_2_delay_1_36;
    io_A_Valid_2_delay_3_34 <= io_A_Valid_2_delay_2_35;
    io_A_Valid_2_delay_4_33 <= io_A_Valid_2_delay_3_34;
    io_A_Valid_2_delay_5_32 <= io_A_Valid_2_delay_4_33;
    io_A_Valid_2_delay_6_31 <= io_A_Valid_2_delay_5_32;
    io_A_Valid_2_delay_7_30 <= io_A_Valid_2_delay_6_31;
    io_A_Valid_2_delay_8_29 <= io_A_Valid_2_delay_7_30;
    io_A_Valid_2_delay_9_28 <= io_A_Valid_2_delay_8_29;
    io_A_Valid_2_delay_10_27 <= io_A_Valid_2_delay_9_28;
    io_A_Valid_2_delay_11_26 <= io_A_Valid_2_delay_10_27;
    io_A_Valid_2_delay_12_25 <= io_A_Valid_2_delay_11_26;
    io_A_Valid_2_delay_13_24 <= io_A_Valid_2_delay_12_25;
    io_A_Valid_2_delay_14_23 <= io_A_Valid_2_delay_13_24;
    io_A_Valid_2_delay_15_22 <= io_A_Valid_2_delay_14_23;
    io_A_Valid_2_delay_16_21 <= io_A_Valid_2_delay_15_22;
    io_A_Valid_2_delay_17_20 <= io_A_Valid_2_delay_16_21;
    io_A_Valid_2_delay_18_19 <= io_A_Valid_2_delay_17_20;
    io_A_Valid_2_delay_19_18 <= io_A_Valid_2_delay_18_19;
    io_A_Valid_2_delay_20_17 <= io_A_Valid_2_delay_19_18;
    io_A_Valid_2_delay_21_16 <= io_A_Valid_2_delay_20_17;
    io_A_Valid_2_delay_22_15 <= io_A_Valid_2_delay_21_16;
    io_A_Valid_2_delay_23_14 <= io_A_Valid_2_delay_22_15;
    io_A_Valid_2_delay_24_13 <= io_A_Valid_2_delay_23_14;
    io_A_Valid_2_delay_25_12 <= io_A_Valid_2_delay_24_13;
    io_A_Valid_2_delay_26_11 <= io_A_Valid_2_delay_25_12;
    io_A_Valid_2_delay_27_10 <= io_A_Valid_2_delay_26_11;
    io_A_Valid_2_delay_28_9 <= io_A_Valid_2_delay_27_10;
    io_A_Valid_2_delay_29_8 <= io_A_Valid_2_delay_28_9;
    io_A_Valid_2_delay_30_7 <= io_A_Valid_2_delay_29_8;
    io_A_Valid_2_delay_31_6 <= io_A_Valid_2_delay_30_7;
    io_A_Valid_2_delay_32_5 <= io_A_Valid_2_delay_31_6;
    io_A_Valid_2_delay_33_4 <= io_A_Valid_2_delay_32_5;
    io_A_Valid_2_delay_34_3 <= io_A_Valid_2_delay_33_4;
    io_A_Valid_2_delay_35_2 <= io_A_Valid_2_delay_34_3;
    io_A_Valid_2_delay_36_1 <= io_A_Valid_2_delay_35_2;
    io_A_Valid_2_delay_37 <= io_A_Valid_2_delay_36_1;
    io_B_Valid_37_delay_1_1 <= io_B_Valid_37;
    io_B_Valid_37_delay_2 <= io_B_Valid_37_delay_1_1;
    io_A_Valid_2_delay_1_37 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_36 <= io_A_Valid_2_delay_1_37;
    io_A_Valid_2_delay_3_35 <= io_A_Valid_2_delay_2_36;
    io_A_Valid_2_delay_4_34 <= io_A_Valid_2_delay_3_35;
    io_A_Valid_2_delay_5_33 <= io_A_Valid_2_delay_4_34;
    io_A_Valid_2_delay_6_32 <= io_A_Valid_2_delay_5_33;
    io_A_Valid_2_delay_7_31 <= io_A_Valid_2_delay_6_32;
    io_A_Valid_2_delay_8_30 <= io_A_Valid_2_delay_7_31;
    io_A_Valid_2_delay_9_29 <= io_A_Valid_2_delay_8_30;
    io_A_Valid_2_delay_10_28 <= io_A_Valid_2_delay_9_29;
    io_A_Valid_2_delay_11_27 <= io_A_Valid_2_delay_10_28;
    io_A_Valid_2_delay_12_26 <= io_A_Valid_2_delay_11_27;
    io_A_Valid_2_delay_13_25 <= io_A_Valid_2_delay_12_26;
    io_A_Valid_2_delay_14_24 <= io_A_Valid_2_delay_13_25;
    io_A_Valid_2_delay_15_23 <= io_A_Valid_2_delay_14_24;
    io_A_Valid_2_delay_16_22 <= io_A_Valid_2_delay_15_23;
    io_A_Valid_2_delay_17_21 <= io_A_Valid_2_delay_16_22;
    io_A_Valid_2_delay_18_20 <= io_A_Valid_2_delay_17_21;
    io_A_Valid_2_delay_19_19 <= io_A_Valid_2_delay_18_20;
    io_A_Valid_2_delay_20_18 <= io_A_Valid_2_delay_19_19;
    io_A_Valid_2_delay_21_17 <= io_A_Valid_2_delay_20_18;
    io_A_Valid_2_delay_22_16 <= io_A_Valid_2_delay_21_17;
    io_A_Valid_2_delay_23_15 <= io_A_Valid_2_delay_22_16;
    io_A_Valid_2_delay_24_14 <= io_A_Valid_2_delay_23_15;
    io_A_Valid_2_delay_25_13 <= io_A_Valid_2_delay_24_14;
    io_A_Valid_2_delay_26_12 <= io_A_Valid_2_delay_25_13;
    io_A_Valid_2_delay_27_11 <= io_A_Valid_2_delay_26_12;
    io_A_Valid_2_delay_28_10 <= io_A_Valid_2_delay_27_11;
    io_A_Valid_2_delay_29_9 <= io_A_Valid_2_delay_28_10;
    io_A_Valid_2_delay_30_8 <= io_A_Valid_2_delay_29_9;
    io_A_Valid_2_delay_31_7 <= io_A_Valid_2_delay_30_8;
    io_A_Valid_2_delay_32_6 <= io_A_Valid_2_delay_31_7;
    io_A_Valid_2_delay_33_5 <= io_A_Valid_2_delay_32_6;
    io_A_Valid_2_delay_34_4 <= io_A_Valid_2_delay_33_5;
    io_A_Valid_2_delay_35_3 <= io_A_Valid_2_delay_34_4;
    io_A_Valid_2_delay_36_2 <= io_A_Valid_2_delay_35_3;
    io_A_Valid_2_delay_37_1 <= io_A_Valid_2_delay_36_2;
    io_A_Valid_2_delay_38 <= io_A_Valid_2_delay_37_1;
    io_B_Valid_38_delay_1_1 <= io_B_Valid_38;
    io_B_Valid_38_delay_2 <= io_B_Valid_38_delay_1_1;
    io_A_Valid_2_delay_1_38 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_37 <= io_A_Valid_2_delay_1_38;
    io_A_Valid_2_delay_3_36 <= io_A_Valid_2_delay_2_37;
    io_A_Valid_2_delay_4_35 <= io_A_Valid_2_delay_3_36;
    io_A_Valid_2_delay_5_34 <= io_A_Valid_2_delay_4_35;
    io_A_Valid_2_delay_6_33 <= io_A_Valid_2_delay_5_34;
    io_A_Valid_2_delay_7_32 <= io_A_Valid_2_delay_6_33;
    io_A_Valid_2_delay_8_31 <= io_A_Valid_2_delay_7_32;
    io_A_Valid_2_delay_9_30 <= io_A_Valid_2_delay_8_31;
    io_A_Valid_2_delay_10_29 <= io_A_Valid_2_delay_9_30;
    io_A_Valid_2_delay_11_28 <= io_A_Valid_2_delay_10_29;
    io_A_Valid_2_delay_12_27 <= io_A_Valid_2_delay_11_28;
    io_A_Valid_2_delay_13_26 <= io_A_Valid_2_delay_12_27;
    io_A_Valid_2_delay_14_25 <= io_A_Valid_2_delay_13_26;
    io_A_Valid_2_delay_15_24 <= io_A_Valid_2_delay_14_25;
    io_A_Valid_2_delay_16_23 <= io_A_Valid_2_delay_15_24;
    io_A_Valid_2_delay_17_22 <= io_A_Valid_2_delay_16_23;
    io_A_Valid_2_delay_18_21 <= io_A_Valid_2_delay_17_22;
    io_A_Valid_2_delay_19_20 <= io_A_Valid_2_delay_18_21;
    io_A_Valid_2_delay_20_19 <= io_A_Valid_2_delay_19_20;
    io_A_Valid_2_delay_21_18 <= io_A_Valid_2_delay_20_19;
    io_A_Valid_2_delay_22_17 <= io_A_Valid_2_delay_21_18;
    io_A_Valid_2_delay_23_16 <= io_A_Valid_2_delay_22_17;
    io_A_Valid_2_delay_24_15 <= io_A_Valid_2_delay_23_16;
    io_A_Valid_2_delay_25_14 <= io_A_Valid_2_delay_24_15;
    io_A_Valid_2_delay_26_13 <= io_A_Valid_2_delay_25_14;
    io_A_Valid_2_delay_27_12 <= io_A_Valid_2_delay_26_13;
    io_A_Valid_2_delay_28_11 <= io_A_Valid_2_delay_27_12;
    io_A_Valid_2_delay_29_10 <= io_A_Valid_2_delay_28_11;
    io_A_Valid_2_delay_30_9 <= io_A_Valid_2_delay_29_10;
    io_A_Valid_2_delay_31_8 <= io_A_Valid_2_delay_30_9;
    io_A_Valid_2_delay_32_7 <= io_A_Valid_2_delay_31_8;
    io_A_Valid_2_delay_33_6 <= io_A_Valid_2_delay_32_7;
    io_A_Valid_2_delay_34_5 <= io_A_Valid_2_delay_33_6;
    io_A_Valid_2_delay_35_4 <= io_A_Valid_2_delay_34_5;
    io_A_Valid_2_delay_36_3 <= io_A_Valid_2_delay_35_4;
    io_A_Valid_2_delay_37_2 <= io_A_Valid_2_delay_36_3;
    io_A_Valid_2_delay_38_1 <= io_A_Valid_2_delay_37_2;
    io_A_Valid_2_delay_39 <= io_A_Valid_2_delay_38_1;
    io_B_Valid_39_delay_1_1 <= io_B_Valid_39;
    io_B_Valid_39_delay_2 <= io_B_Valid_39_delay_1_1;
    io_A_Valid_2_delay_1_39 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_38 <= io_A_Valid_2_delay_1_39;
    io_A_Valid_2_delay_3_37 <= io_A_Valid_2_delay_2_38;
    io_A_Valid_2_delay_4_36 <= io_A_Valid_2_delay_3_37;
    io_A_Valid_2_delay_5_35 <= io_A_Valid_2_delay_4_36;
    io_A_Valid_2_delay_6_34 <= io_A_Valid_2_delay_5_35;
    io_A_Valid_2_delay_7_33 <= io_A_Valid_2_delay_6_34;
    io_A_Valid_2_delay_8_32 <= io_A_Valid_2_delay_7_33;
    io_A_Valid_2_delay_9_31 <= io_A_Valid_2_delay_8_32;
    io_A_Valid_2_delay_10_30 <= io_A_Valid_2_delay_9_31;
    io_A_Valid_2_delay_11_29 <= io_A_Valid_2_delay_10_30;
    io_A_Valid_2_delay_12_28 <= io_A_Valid_2_delay_11_29;
    io_A_Valid_2_delay_13_27 <= io_A_Valid_2_delay_12_28;
    io_A_Valid_2_delay_14_26 <= io_A_Valid_2_delay_13_27;
    io_A_Valid_2_delay_15_25 <= io_A_Valid_2_delay_14_26;
    io_A_Valid_2_delay_16_24 <= io_A_Valid_2_delay_15_25;
    io_A_Valid_2_delay_17_23 <= io_A_Valid_2_delay_16_24;
    io_A_Valid_2_delay_18_22 <= io_A_Valid_2_delay_17_23;
    io_A_Valid_2_delay_19_21 <= io_A_Valid_2_delay_18_22;
    io_A_Valid_2_delay_20_20 <= io_A_Valid_2_delay_19_21;
    io_A_Valid_2_delay_21_19 <= io_A_Valid_2_delay_20_20;
    io_A_Valid_2_delay_22_18 <= io_A_Valid_2_delay_21_19;
    io_A_Valid_2_delay_23_17 <= io_A_Valid_2_delay_22_18;
    io_A_Valid_2_delay_24_16 <= io_A_Valid_2_delay_23_17;
    io_A_Valid_2_delay_25_15 <= io_A_Valid_2_delay_24_16;
    io_A_Valid_2_delay_26_14 <= io_A_Valid_2_delay_25_15;
    io_A_Valid_2_delay_27_13 <= io_A_Valid_2_delay_26_14;
    io_A_Valid_2_delay_28_12 <= io_A_Valid_2_delay_27_13;
    io_A_Valid_2_delay_29_11 <= io_A_Valid_2_delay_28_12;
    io_A_Valid_2_delay_30_10 <= io_A_Valid_2_delay_29_11;
    io_A_Valid_2_delay_31_9 <= io_A_Valid_2_delay_30_10;
    io_A_Valid_2_delay_32_8 <= io_A_Valid_2_delay_31_9;
    io_A_Valid_2_delay_33_7 <= io_A_Valid_2_delay_32_8;
    io_A_Valid_2_delay_34_6 <= io_A_Valid_2_delay_33_7;
    io_A_Valid_2_delay_35_5 <= io_A_Valid_2_delay_34_6;
    io_A_Valid_2_delay_36_4 <= io_A_Valid_2_delay_35_5;
    io_A_Valid_2_delay_37_3 <= io_A_Valid_2_delay_36_4;
    io_A_Valid_2_delay_38_2 <= io_A_Valid_2_delay_37_3;
    io_A_Valid_2_delay_39_1 <= io_A_Valid_2_delay_38_2;
    io_A_Valid_2_delay_40 <= io_A_Valid_2_delay_39_1;
    io_B_Valid_40_delay_1_1 <= io_B_Valid_40;
    io_B_Valid_40_delay_2 <= io_B_Valid_40_delay_1_1;
    io_A_Valid_2_delay_1_40 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_39 <= io_A_Valid_2_delay_1_40;
    io_A_Valid_2_delay_3_38 <= io_A_Valid_2_delay_2_39;
    io_A_Valid_2_delay_4_37 <= io_A_Valid_2_delay_3_38;
    io_A_Valid_2_delay_5_36 <= io_A_Valid_2_delay_4_37;
    io_A_Valid_2_delay_6_35 <= io_A_Valid_2_delay_5_36;
    io_A_Valid_2_delay_7_34 <= io_A_Valid_2_delay_6_35;
    io_A_Valid_2_delay_8_33 <= io_A_Valid_2_delay_7_34;
    io_A_Valid_2_delay_9_32 <= io_A_Valid_2_delay_8_33;
    io_A_Valid_2_delay_10_31 <= io_A_Valid_2_delay_9_32;
    io_A_Valid_2_delay_11_30 <= io_A_Valid_2_delay_10_31;
    io_A_Valid_2_delay_12_29 <= io_A_Valid_2_delay_11_30;
    io_A_Valid_2_delay_13_28 <= io_A_Valid_2_delay_12_29;
    io_A_Valid_2_delay_14_27 <= io_A_Valid_2_delay_13_28;
    io_A_Valid_2_delay_15_26 <= io_A_Valid_2_delay_14_27;
    io_A_Valid_2_delay_16_25 <= io_A_Valid_2_delay_15_26;
    io_A_Valid_2_delay_17_24 <= io_A_Valid_2_delay_16_25;
    io_A_Valid_2_delay_18_23 <= io_A_Valid_2_delay_17_24;
    io_A_Valid_2_delay_19_22 <= io_A_Valid_2_delay_18_23;
    io_A_Valid_2_delay_20_21 <= io_A_Valid_2_delay_19_22;
    io_A_Valid_2_delay_21_20 <= io_A_Valid_2_delay_20_21;
    io_A_Valid_2_delay_22_19 <= io_A_Valid_2_delay_21_20;
    io_A_Valid_2_delay_23_18 <= io_A_Valid_2_delay_22_19;
    io_A_Valid_2_delay_24_17 <= io_A_Valid_2_delay_23_18;
    io_A_Valid_2_delay_25_16 <= io_A_Valid_2_delay_24_17;
    io_A_Valid_2_delay_26_15 <= io_A_Valid_2_delay_25_16;
    io_A_Valid_2_delay_27_14 <= io_A_Valid_2_delay_26_15;
    io_A_Valid_2_delay_28_13 <= io_A_Valid_2_delay_27_14;
    io_A_Valid_2_delay_29_12 <= io_A_Valid_2_delay_28_13;
    io_A_Valid_2_delay_30_11 <= io_A_Valid_2_delay_29_12;
    io_A_Valid_2_delay_31_10 <= io_A_Valid_2_delay_30_11;
    io_A_Valid_2_delay_32_9 <= io_A_Valid_2_delay_31_10;
    io_A_Valid_2_delay_33_8 <= io_A_Valid_2_delay_32_9;
    io_A_Valid_2_delay_34_7 <= io_A_Valid_2_delay_33_8;
    io_A_Valid_2_delay_35_6 <= io_A_Valid_2_delay_34_7;
    io_A_Valid_2_delay_36_5 <= io_A_Valid_2_delay_35_6;
    io_A_Valid_2_delay_37_4 <= io_A_Valid_2_delay_36_5;
    io_A_Valid_2_delay_38_3 <= io_A_Valid_2_delay_37_4;
    io_A_Valid_2_delay_39_2 <= io_A_Valid_2_delay_38_3;
    io_A_Valid_2_delay_40_1 <= io_A_Valid_2_delay_39_2;
    io_A_Valid_2_delay_41 <= io_A_Valid_2_delay_40_1;
    io_B_Valid_41_delay_1_1 <= io_B_Valid_41;
    io_B_Valid_41_delay_2 <= io_B_Valid_41_delay_1_1;
    io_A_Valid_2_delay_1_41 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_40 <= io_A_Valid_2_delay_1_41;
    io_A_Valid_2_delay_3_39 <= io_A_Valid_2_delay_2_40;
    io_A_Valid_2_delay_4_38 <= io_A_Valid_2_delay_3_39;
    io_A_Valid_2_delay_5_37 <= io_A_Valid_2_delay_4_38;
    io_A_Valid_2_delay_6_36 <= io_A_Valid_2_delay_5_37;
    io_A_Valid_2_delay_7_35 <= io_A_Valid_2_delay_6_36;
    io_A_Valid_2_delay_8_34 <= io_A_Valid_2_delay_7_35;
    io_A_Valid_2_delay_9_33 <= io_A_Valid_2_delay_8_34;
    io_A_Valid_2_delay_10_32 <= io_A_Valid_2_delay_9_33;
    io_A_Valid_2_delay_11_31 <= io_A_Valid_2_delay_10_32;
    io_A_Valid_2_delay_12_30 <= io_A_Valid_2_delay_11_31;
    io_A_Valid_2_delay_13_29 <= io_A_Valid_2_delay_12_30;
    io_A_Valid_2_delay_14_28 <= io_A_Valid_2_delay_13_29;
    io_A_Valid_2_delay_15_27 <= io_A_Valid_2_delay_14_28;
    io_A_Valid_2_delay_16_26 <= io_A_Valid_2_delay_15_27;
    io_A_Valid_2_delay_17_25 <= io_A_Valid_2_delay_16_26;
    io_A_Valid_2_delay_18_24 <= io_A_Valid_2_delay_17_25;
    io_A_Valid_2_delay_19_23 <= io_A_Valid_2_delay_18_24;
    io_A_Valid_2_delay_20_22 <= io_A_Valid_2_delay_19_23;
    io_A_Valid_2_delay_21_21 <= io_A_Valid_2_delay_20_22;
    io_A_Valid_2_delay_22_20 <= io_A_Valid_2_delay_21_21;
    io_A_Valid_2_delay_23_19 <= io_A_Valid_2_delay_22_20;
    io_A_Valid_2_delay_24_18 <= io_A_Valid_2_delay_23_19;
    io_A_Valid_2_delay_25_17 <= io_A_Valid_2_delay_24_18;
    io_A_Valid_2_delay_26_16 <= io_A_Valid_2_delay_25_17;
    io_A_Valid_2_delay_27_15 <= io_A_Valid_2_delay_26_16;
    io_A_Valid_2_delay_28_14 <= io_A_Valid_2_delay_27_15;
    io_A_Valid_2_delay_29_13 <= io_A_Valid_2_delay_28_14;
    io_A_Valid_2_delay_30_12 <= io_A_Valid_2_delay_29_13;
    io_A_Valid_2_delay_31_11 <= io_A_Valid_2_delay_30_12;
    io_A_Valid_2_delay_32_10 <= io_A_Valid_2_delay_31_11;
    io_A_Valid_2_delay_33_9 <= io_A_Valid_2_delay_32_10;
    io_A_Valid_2_delay_34_8 <= io_A_Valid_2_delay_33_9;
    io_A_Valid_2_delay_35_7 <= io_A_Valid_2_delay_34_8;
    io_A_Valid_2_delay_36_6 <= io_A_Valid_2_delay_35_7;
    io_A_Valid_2_delay_37_5 <= io_A_Valid_2_delay_36_6;
    io_A_Valid_2_delay_38_4 <= io_A_Valid_2_delay_37_5;
    io_A_Valid_2_delay_39_3 <= io_A_Valid_2_delay_38_4;
    io_A_Valid_2_delay_40_2 <= io_A_Valid_2_delay_39_3;
    io_A_Valid_2_delay_41_1 <= io_A_Valid_2_delay_40_2;
    io_A_Valid_2_delay_42 <= io_A_Valid_2_delay_41_1;
    io_B_Valid_42_delay_1_1 <= io_B_Valid_42;
    io_B_Valid_42_delay_2 <= io_B_Valid_42_delay_1_1;
    io_A_Valid_2_delay_1_42 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_41 <= io_A_Valid_2_delay_1_42;
    io_A_Valid_2_delay_3_40 <= io_A_Valid_2_delay_2_41;
    io_A_Valid_2_delay_4_39 <= io_A_Valid_2_delay_3_40;
    io_A_Valid_2_delay_5_38 <= io_A_Valid_2_delay_4_39;
    io_A_Valid_2_delay_6_37 <= io_A_Valid_2_delay_5_38;
    io_A_Valid_2_delay_7_36 <= io_A_Valid_2_delay_6_37;
    io_A_Valid_2_delay_8_35 <= io_A_Valid_2_delay_7_36;
    io_A_Valid_2_delay_9_34 <= io_A_Valid_2_delay_8_35;
    io_A_Valid_2_delay_10_33 <= io_A_Valid_2_delay_9_34;
    io_A_Valid_2_delay_11_32 <= io_A_Valid_2_delay_10_33;
    io_A_Valid_2_delay_12_31 <= io_A_Valid_2_delay_11_32;
    io_A_Valid_2_delay_13_30 <= io_A_Valid_2_delay_12_31;
    io_A_Valid_2_delay_14_29 <= io_A_Valid_2_delay_13_30;
    io_A_Valid_2_delay_15_28 <= io_A_Valid_2_delay_14_29;
    io_A_Valid_2_delay_16_27 <= io_A_Valid_2_delay_15_28;
    io_A_Valid_2_delay_17_26 <= io_A_Valid_2_delay_16_27;
    io_A_Valid_2_delay_18_25 <= io_A_Valid_2_delay_17_26;
    io_A_Valid_2_delay_19_24 <= io_A_Valid_2_delay_18_25;
    io_A_Valid_2_delay_20_23 <= io_A_Valid_2_delay_19_24;
    io_A_Valid_2_delay_21_22 <= io_A_Valid_2_delay_20_23;
    io_A_Valid_2_delay_22_21 <= io_A_Valid_2_delay_21_22;
    io_A_Valid_2_delay_23_20 <= io_A_Valid_2_delay_22_21;
    io_A_Valid_2_delay_24_19 <= io_A_Valid_2_delay_23_20;
    io_A_Valid_2_delay_25_18 <= io_A_Valid_2_delay_24_19;
    io_A_Valid_2_delay_26_17 <= io_A_Valid_2_delay_25_18;
    io_A_Valid_2_delay_27_16 <= io_A_Valid_2_delay_26_17;
    io_A_Valid_2_delay_28_15 <= io_A_Valid_2_delay_27_16;
    io_A_Valid_2_delay_29_14 <= io_A_Valid_2_delay_28_15;
    io_A_Valid_2_delay_30_13 <= io_A_Valid_2_delay_29_14;
    io_A_Valid_2_delay_31_12 <= io_A_Valid_2_delay_30_13;
    io_A_Valid_2_delay_32_11 <= io_A_Valid_2_delay_31_12;
    io_A_Valid_2_delay_33_10 <= io_A_Valid_2_delay_32_11;
    io_A_Valid_2_delay_34_9 <= io_A_Valid_2_delay_33_10;
    io_A_Valid_2_delay_35_8 <= io_A_Valid_2_delay_34_9;
    io_A_Valid_2_delay_36_7 <= io_A_Valid_2_delay_35_8;
    io_A_Valid_2_delay_37_6 <= io_A_Valid_2_delay_36_7;
    io_A_Valid_2_delay_38_5 <= io_A_Valid_2_delay_37_6;
    io_A_Valid_2_delay_39_4 <= io_A_Valid_2_delay_38_5;
    io_A_Valid_2_delay_40_3 <= io_A_Valid_2_delay_39_4;
    io_A_Valid_2_delay_41_2 <= io_A_Valid_2_delay_40_3;
    io_A_Valid_2_delay_42_1 <= io_A_Valid_2_delay_41_2;
    io_A_Valid_2_delay_43 <= io_A_Valid_2_delay_42_1;
    io_B_Valid_43_delay_1_1 <= io_B_Valid_43;
    io_B_Valid_43_delay_2 <= io_B_Valid_43_delay_1_1;
    io_A_Valid_2_delay_1_43 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_42 <= io_A_Valid_2_delay_1_43;
    io_A_Valid_2_delay_3_41 <= io_A_Valid_2_delay_2_42;
    io_A_Valid_2_delay_4_40 <= io_A_Valid_2_delay_3_41;
    io_A_Valid_2_delay_5_39 <= io_A_Valid_2_delay_4_40;
    io_A_Valid_2_delay_6_38 <= io_A_Valid_2_delay_5_39;
    io_A_Valid_2_delay_7_37 <= io_A_Valid_2_delay_6_38;
    io_A_Valid_2_delay_8_36 <= io_A_Valid_2_delay_7_37;
    io_A_Valid_2_delay_9_35 <= io_A_Valid_2_delay_8_36;
    io_A_Valid_2_delay_10_34 <= io_A_Valid_2_delay_9_35;
    io_A_Valid_2_delay_11_33 <= io_A_Valid_2_delay_10_34;
    io_A_Valid_2_delay_12_32 <= io_A_Valid_2_delay_11_33;
    io_A_Valid_2_delay_13_31 <= io_A_Valid_2_delay_12_32;
    io_A_Valid_2_delay_14_30 <= io_A_Valid_2_delay_13_31;
    io_A_Valid_2_delay_15_29 <= io_A_Valid_2_delay_14_30;
    io_A_Valid_2_delay_16_28 <= io_A_Valid_2_delay_15_29;
    io_A_Valid_2_delay_17_27 <= io_A_Valid_2_delay_16_28;
    io_A_Valid_2_delay_18_26 <= io_A_Valid_2_delay_17_27;
    io_A_Valid_2_delay_19_25 <= io_A_Valid_2_delay_18_26;
    io_A_Valid_2_delay_20_24 <= io_A_Valid_2_delay_19_25;
    io_A_Valid_2_delay_21_23 <= io_A_Valid_2_delay_20_24;
    io_A_Valid_2_delay_22_22 <= io_A_Valid_2_delay_21_23;
    io_A_Valid_2_delay_23_21 <= io_A_Valid_2_delay_22_22;
    io_A_Valid_2_delay_24_20 <= io_A_Valid_2_delay_23_21;
    io_A_Valid_2_delay_25_19 <= io_A_Valid_2_delay_24_20;
    io_A_Valid_2_delay_26_18 <= io_A_Valid_2_delay_25_19;
    io_A_Valid_2_delay_27_17 <= io_A_Valid_2_delay_26_18;
    io_A_Valid_2_delay_28_16 <= io_A_Valid_2_delay_27_17;
    io_A_Valid_2_delay_29_15 <= io_A_Valid_2_delay_28_16;
    io_A_Valid_2_delay_30_14 <= io_A_Valid_2_delay_29_15;
    io_A_Valid_2_delay_31_13 <= io_A_Valid_2_delay_30_14;
    io_A_Valid_2_delay_32_12 <= io_A_Valid_2_delay_31_13;
    io_A_Valid_2_delay_33_11 <= io_A_Valid_2_delay_32_12;
    io_A_Valid_2_delay_34_10 <= io_A_Valid_2_delay_33_11;
    io_A_Valid_2_delay_35_9 <= io_A_Valid_2_delay_34_10;
    io_A_Valid_2_delay_36_8 <= io_A_Valid_2_delay_35_9;
    io_A_Valid_2_delay_37_7 <= io_A_Valid_2_delay_36_8;
    io_A_Valid_2_delay_38_6 <= io_A_Valid_2_delay_37_7;
    io_A_Valid_2_delay_39_5 <= io_A_Valid_2_delay_38_6;
    io_A_Valid_2_delay_40_4 <= io_A_Valid_2_delay_39_5;
    io_A_Valid_2_delay_41_3 <= io_A_Valid_2_delay_40_4;
    io_A_Valid_2_delay_42_2 <= io_A_Valid_2_delay_41_3;
    io_A_Valid_2_delay_43_1 <= io_A_Valid_2_delay_42_2;
    io_A_Valid_2_delay_44 <= io_A_Valid_2_delay_43_1;
    io_B_Valid_44_delay_1_1 <= io_B_Valid_44;
    io_B_Valid_44_delay_2 <= io_B_Valid_44_delay_1_1;
    io_A_Valid_2_delay_1_44 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_43 <= io_A_Valid_2_delay_1_44;
    io_A_Valid_2_delay_3_42 <= io_A_Valid_2_delay_2_43;
    io_A_Valid_2_delay_4_41 <= io_A_Valid_2_delay_3_42;
    io_A_Valid_2_delay_5_40 <= io_A_Valid_2_delay_4_41;
    io_A_Valid_2_delay_6_39 <= io_A_Valid_2_delay_5_40;
    io_A_Valid_2_delay_7_38 <= io_A_Valid_2_delay_6_39;
    io_A_Valid_2_delay_8_37 <= io_A_Valid_2_delay_7_38;
    io_A_Valid_2_delay_9_36 <= io_A_Valid_2_delay_8_37;
    io_A_Valid_2_delay_10_35 <= io_A_Valid_2_delay_9_36;
    io_A_Valid_2_delay_11_34 <= io_A_Valid_2_delay_10_35;
    io_A_Valid_2_delay_12_33 <= io_A_Valid_2_delay_11_34;
    io_A_Valid_2_delay_13_32 <= io_A_Valid_2_delay_12_33;
    io_A_Valid_2_delay_14_31 <= io_A_Valid_2_delay_13_32;
    io_A_Valid_2_delay_15_30 <= io_A_Valid_2_delay_14_31;
    io_A_Valid_2_delay_16_29 <= io_A_Valid_2_delay_15_30;
    io_A_Valid_2_delay_17_28 <= io_A_Valid_2_delay_16_29;
    io_A_Valid_2_delay_18_27 <= io_A_Valid_2_delay_17_28;
    io_A_Valid_2_delay_19_26 <= io_A_Valid_2_delay_18_27;
    io_A_Valid_2_delay_20_25 <= io_A_Valid_2_delay_19_26;
    io_A_Valid_2_delay_21_24 <= io_A_Valid_2_delay_20_25;
    io_A_Valid_2_delay_22_23 <= io_A_Valid_2_delay_21_24;
    io_A_Valid_2_delay_23_22 <= io_A_Valid_2_delay_22_23;
    io_A_Valid_2_delay_24_21 <= io_A_Valid_2_delay_23_22;
    io_A_Valid_2_delay_25_20 <= io_A_Valid_2_delay_24_21;
    io_A_Valid_2_delay_26_19 <= io_A_Valid_2_delay_25_20;
    io_A_Valid_2_delay_27_18 <= io_A_Valid_2_delay_26_19;
    io_A_Valid_2_delay_28_17 <= io_A_Valid_2_delay_27_18;
    io_A_Valid_2_delay_29_16 <= io_A_Valid_2_delay_28_17;
    io_A_Valid_2_delay_30_15 <= io_A_Valid_2_delay_29_16;
    io_A_Valid_2_delay_31_14 <= io_A_Valid_2_delay_30_15;
    io_A_Valid_2_delay_32_13 <= io_A_Valid_2_delay_31_14;
    io_A_Valid_2_delay_33_12 <= io_A_Valid_2_delay_32_13;
    io_A_Valid_2_delay_34_11 <= io_A_Valid_2_delay_33_12;
    io_A_Valid_2_delay_35_10 <= io_A_Valid_2_delay_34_11;
    io_A_Valid_2_delay_36_9 <= io_A_Valid_2_delay_35_10;
    io_A_Valid_2_delay_37_8 <= io_A_Valid_2_delay_36_9;
    io_A_Valid_2_delay_38_7 <= io_A_Valid_2_delay_37_8;
    io_A_Valid_2_delay_39_6 <= io_A_Valid_2_delay_38_7;
    io_A_Valid_2_delay_40_5 <= io_A_Valid_2_delay_39_6;
    io_A_Valid_2_delay_41_4 <= io_A_Valid_2_delay_40_5;
    io_A_Valid_2_delay_42_3 <= io_A_Valid_2_delay_41_4;
    io_A_Valid_2_delay_43_2 <= io_A_Valid_2_delay_42_3;
    io_A_Valid_2_delay_44_1 <= io_A_Valid_2_delay_43_2;
    io_A_Valid_2_delay_45 <= io_A_Valid_2_delay_44_1;
    io_B_Valid_45_delay_1_1 <= io_B_Valid_45;
    io_B_Valid_45_delay_2 <= io_B_Valid_45_delay_1_1;
    io_A_Valid_2_delay_1_45 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_44 <= io_A_Valid_2_delay_1_45;
    io_A_Valid_2_delay_3_43 <= io_A_Valid_2_delay_2_44;
    io_A_Valid_2_delay_4_42 <= io_A_Valid_2_delay_3_43;
    io_A_Valid_2_delay_5_41 <= io_A_Valid_2_delay_4_42;
    io_A_Valid_2_delay_6_40 <= io_A_Valid_2_delay_5_41;
    io_A_Valid_2_delay_7_39 <= io_A_Valid_2_delay_6_40;
    io_A_Valid_2_delay_8_38 <= io_A_Valid_2_delay_7_39;
    io_A_Valid_2_delay_9_37 <= io_A_Valid_2_delay_8_38;
    io_A_Valid_2_delay_10_36 <= io_A_Valid_2_delay_9_37;
    io_A_Valid_2_delay_11_35 <= io_A_Valid_2_delay_10_36;
    io_A_Valid_2_delay_12_34 <= io_A_Valid_2_delay_11_35;
    io_A_Valid_2_delay_13_33 <= io_A_Valid_2_delay_12_34;
    io_A_Valid_2_delay_14_32 <= io_A_Valid_2_delay_13_33;
    io_A_Valid_2_delay_15_31 <= io_A_Valid_2_delay_14_32;
    io_A_Valid_2_delay_16_30 <= io_A_Valid_2_delay_15_31;
    io_A_Valid_2_delay_17_29 <= io_A_Valid_2_delay_16_30;
    io_A_Valid_2_delay_18_28 <= io_A_Valid_2_delay_17_29;
    io_A_Valid_2_delay_19_27 <= io_A_Valid_2_delay_18_28;
    io_A_Valid_2_delay_20_26 <= io_A_Valid_2_delay_19_27;
    io_A_Valid_2_delay_21_25 <= io_A_Valid_2_delay_20_26;
    io_A_Valid_2_delay_22_24 <= io_A_Valid_2_delay_21_25;
    io_A_Valid_2_delay_23_23 <= io_A_Valid_2_delay_22_24;
    io_A_Valid_2_delay_24_22 <= io_A_Valid_2_delay_23_23;
    io_A_Valid_2_delay_25_21 <= io_A_Valid_2_delay_24_22;
    io_A_Valid_2_delay_26_20 <= io_A_Valid_2_delay_25_21;
    io_A_Valid_2_delay_27_19 <= io_A_Valid_2_delay_26_20;
    io_A_Valid_2_delay_28_18 <= io_A_Valid_2_delay_27_19;
    io_A_Valid_2_delay_29_17 <= io_A_Valid_2_delay_28_18;
    io_A_Valid_2_delay_30_16 <= io_A_Valid_2_delay_29_17;
    io_A_Valid_2_delay_31_15 <= io_A_Valid_2_delay_30_16;
    io_A_Valid_2_delay_32_14 <= io_A_Valid_2_delay_31_15;
    io_A_Valid_2_delay_33_13 <= io_A_Valid_2_delay_32_14;
    io_A_Valid_2_delay_34_12 <= io_A_Valid_2_delay_33_13;
    io_A_Valid_2_delay_35_11 <= io_A_Valid_2_delay_34_12;
    io_A_Valid_2_delay_36_10 <= io_A_Valid_2_delay_35_11;
    io_A_Valid_2_delay_37_9 <= io_A_Valid_2_delay_36_10;
    io_A_Valid_2_delay_38_8 <= io_A_Valid_2_delay_37_9;
    io_A_Valid_2_delay_39_7 <= io_A_Valid_2_delay_38_8;
    io_A_Valid_2_delay_40_6 <= io_A_Valid_2_delay_39_7;
    io_A_Valid_2_delay_41_5 <= io_A_Valid_2_delay_40_6;
    io_A_Valid_2_delay_42_4 <= io_A_Valid_2_delay_41_5;
    io_A_Valid_2_delay_43_3 <= io_A_Valid_2_delay_42_4;
    io_A_Valid_2_delay_44_2 <= io_A_Valid_2_delay_43_3;
    io_A_Valid_2_delay_45_1 <= io_A_Valid_2_delay_44_2;
    io_A_Valid_2_delay_46 <= io_A_Valid_2_delay_45_1;
    io_B_Valid_46_delay_1_1 <= io_B_Valid_46;
    io_B_Valid_46_delay_2 <= io_B_Valid_46_delay_1_1;
    io_A_Valid_2_delay_1_46 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_45 <= io_A_Valid_2_delay_1_46;
    io_A_Valid_2_delay_3_44 <= io_A_Valid_2_delay_2_45;
    io_A_Valid_2_delay_4_43 <= io_A_Valid_2_delay_3_44;
    io_A_Valid_2_delay_5_42 <= io_A_Valid_2_delay_4_43;
    io_A_Valid_2_delay_6_41 <= io_A_Valid_2_delay_5_42;
    io_A_Valid_2_delay_7_40 <= io_A_Valid_2_delay_6_41;
    io_A_Valid_2_delay_8_39 <= io_A_Valid_2_delay_7_40;
    io_A_Valid_2_delay_9_38 <= io_A_Valid_2_delay_8_39;
    io_A_Valid_2_delay_10_37 <= io_A_Valid_2_delay_9_38;
    io_A_Valid_2_delay_11_36 <= io_A_Valid_2_delay_10_37;
    io_A_Valid_2_delay_12_35 <= io_A_Valid_2_delay_11_36;
    io_A_Valid_2_delay_13_34 <= io_A_Valid_2_delay_12_35;
    io_A_Valid_2_delay_14_33 <= io_A_Valid_2_delay_13_34;
    io_A_Valid_2_delay_15_32 <= io_A_Valid_2_delay_14_33;
    io_A_Valid_2_delay_16_31 <= io_A_Valid_2_delay_15_32;
    io_A_Valid_2_delay_17_30 <= io_A_Valid_2_delay_16_31;
    io_A_Valid_2_delay_18_29 <= io_A_Valid_2_delay_17_30;
    io_A_Valid_2_delay_19_28 <= io_A_Valid_2_delay_18_29;
    io_A_Valid_2_delay_20_27 <= io_A_Valid_2_delay_19_28;
    io_A_Valid_2_delay_21_26 <= io_A_Valid_2_delay_20_27;
    io_A_Valid_2_delay_22_25 <= io_A_Valid_2_delay_21_26;
    io_A_Valid_2_delay_23_24 <= io_A_Valid_2_delay_22_25;
    io_A_Valid_2_delay_24_23 <= io_A_Valid_2_delay_23_24;
    io_A_Valid_2_delay_25_22 <= io_A_Valid_2_delay_24_23;
    io_A_Valid_2_delay_26_21 <= io_A_Valid_2_delay_25_22;
    io_A_Valid_2_delay_27_20 <= io_A_Valid_2_delay_26_21;
    io_A_Valid_2_delay_28_19 <= io_A_Valid_2_delay_27_20;
    io_A_Valid_2_delay_29_18 <= io_A_Valid_2_delay_28_19;
    io_A_Valid_2_delay_30_17 <= io_A_Valid_2_delay_29_18;
    io_A_Valid_2_delay_31_16 <= io_A_Valid_2_delay_30_17;
    io_A_Valid_2_delay_32_15 <= io_A_Valid_2_delay_31_16;
    io_A_Valid_2_delay_33_14 <= io_A_Valid_2_delay_32_15;
    io_A_Valid_2_delay_34_13 <= io_A_Valid_2_delay_33_14;
    io_A_Valid_2_delay_35_12 <= io_A_Valid_2_delay_34_13;
    io_A_Valid_2_delay_36_11 <= io_A_Valid_2_delay_35_12;
    io_A_Valid_2_delay_37_10 <= io_A_Valid_2_delay_36_11;
    io_A_Valid_2_delay_38_9 <= io_A_Valid_2_delay_37_10;
    io_A_Valid_2_delay_39_8 <= io_A_Valid_2_delay_38_9;
    io_A_Valid_2_delay_40_7 <= io_A_Valid_2_delay_39_8;
    io_A_Valid_2_delay_41_6 <= io_A_Valid_2_delay_40_7;
    io_A_Valid_2_delay_42_5 <= io_A_Valid_2_delay_41_6;
    io_A_Valid_2_delay_43_4 <= io_A_Valid_2_delay_42_5;
    io_A_Valid_2_delay_44_3 <= io_A_Valid_2_delay_43_4;
    io_A_Valid_2_delay_45_2 <= io_A_Valid_2_delay_44_3;
    io_A_Valid_2_delay_46_1 <= io_A_Valid_2_delay_45_2;
    io_A_Valid_2_delay_47 <= io_A_Valid_2_delay_46_1;
    io_B_Valid_47_delay_1_1 <= io_B_Valid_47;
    io_B_Valid_47_delay_2 <= io_B_Valid_47_delay_1_1;
    io_A_Valid_2_delay_1_47 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_46 <= io_A_Valid_2_delay_1_47;
    io_A_Valid_2_delay_3_45 <= io_A_Valid_2_delay_2_46;
    io_A_Valid_2_delay_4_44 <= io_A_Valid_2_delay_3_45;
    io_A_Valid_2_delay_5_43 <= io_A_Valid_2_delay_4_44;
    io_A_Valid_2_delay_6_42 <= io_A_Valid_2_delay_5_43;
    io_A_Valid_2_delay_7_41 <= io_A_Valid_2_delay_6_42;
    io_A_Valid_2_delay_8_40 <= io_A_Valid_2_delay_7_41;
    io_A_Valid_2_delay_9_39 <= io_A_Valid_2_delay_8_40;
    io_A_Valid_2_delay_10_38 <= io_A_Valid_2_delay_9_39;
    io_A_Valid_2_delay_11_37 <= io_A_Valid_2_delay_10_38;
    io_A_Valid_2_delay_12_36 <= io_A_Valid_2_delay_11_37;
    io_A_Valid_2_delay_13_35 <= io_A_Valid_2_delay_12_36;
    io_A_Valid_2_delay_14_34 <= io_A_Valid_2_delay_13_35;
    io_A_Valid_2_delay_15_33 <= io_A_Valid_2_delay_14_34;
    io_A_Valid_2_delay_16_32 <= io_A_Valid_2_delay_15_33;
    io_A_Valid_2_delay_17_31 <= io_A_Valid_2_delay_16_32;
    io_A_Valid_2_delay_18_30 <= io_A_Valid_2_delay_17_31;
    io_A_Valid_2_delay_19_29 <= io_A_Valid_2_delay_18_30;
    io_A_Valid_2_delay_20_28 <= io_A_Valid_2_delay_19_29;
    io_A_Valid_2_delay_21_27 <= io_A_Valid_2_delay_20_28;
    io_A_Valid_2_delay_22_26 <= io_A_Valid_2_delay_21_27;
    io_A_Valid_2_delay_23_25 <= io_A_Valid_2_delay_22_26;
    io_A_Valid_2_delay_24_24 <= io_A_Valid_2_delay_23_25;
    io_A_Valid_2_delay_25_23 <= io_A_Valid_2_delay_24_24;
    io_A_Valid_2_delay_26_22 <= io_A_Valid_2_delay_25_23;
    io_A_Valid_2_delay_27_21 <= io_A_Valid_2_delay_26_22;
    io_A_Valid_2_delay_28_20 <= io_A_Valid_2_delay_27_21;
    io_A_Valid_2_delay_29_19 <= io_A_Valid_2_delay_28_20;
    io_A_Valid_2_delay_30_18 <= io_A_Valid_2_delay_29_19;
    io_A_Valid_2_delay_31_17 <= io_A_Valid_2_delay_30_18;
    io_A_Valid_2_delay_32_16 <= io_A_Valid_2_delay_31_17;
    io_A_Valid_2_delay_33_15 <= io_A_Valid_2_delay_32_16;
    io_A_Valid_2_delay_34_14 <= io_A_Valid_2_delay_33_15;
    io_A_Valid_2_delay_35_13 <= io_A_Valid_2_delay_34_14;
    io_A_Valid_2_delay_36_12 <= io_A_Valid_2_delay_35_13;
    io_A_Valid_2_delay_37_11 <= io_A_Valid_2_delay_36_12;
    io_A_Valid_2_delay_38_10 <= io_A_Valid_2_delay_37_11;
    io_A_Valid_2_delay_39_9 <= io_A_Valid_2_delay_38_10;
    io_A_Valid_2_delay_40_8 <= io_A_Valid_2_delay_39_9;
    io_A_Valid_2_delay_41_7 <= io_A_Valid_2_delay_40_8;
    io_A_Valid_2_delay_42_6 <= io_A_Valid_2_delay_41_7;
    io_A_Valid_2_delay_43_5 <= io_A_Valid_2_delay_42_6;
    io_A_Valid_2_delay_44_4 <= io_A_Valid_2_delay_43_5;
    io_A_Valid_2_delay_45_3 <= io_A_Valid_2_delay_44_4;
    io_A_Valid_2_delay_46_2 <= io_A_Valid_2_delay_45_3;
    io_A_Valid_2_delay_47_1 <= io_A_Valid_2_delay_46_2;
    io_A_Valid_2_delay_48 <= io_A_Valid_2_delay_47_1;
    io_B_Valid_48_delay_1_1 <= io_B_Valid_48;
    io_B_Valid_48_delay_2 <= io_B_Valid_48_delay_1_1;
    io_A_Valid_2_delay_1_48 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_47 <= io_A_Valid_2_delay_1_48;
    io_A_Valid_2_delay_3_46 <= io_A_Valid_2_delay_2_47;
    io_A_Valid_2_delay_4_45 <= io_A_Valid_2_delay_3_46;
    io_A_Valid_2_delay_5_44 <= io_A_Valid_2_delay_4_45;
    io_A_Valid_2_delay_6_43 <= io_A_Valid_2_delay_5_44;
    io_A_Valid_2_delay_7_42 <= io_A_Valid_2_delay_6_43;
    io_A_Valid_2_delay_8_41 <= io_A_Valid_2_delay_7_42;
    io_A_Valid_2_delay_9_40 <= io_A_Valid_2_delay_8_41;
    io_A_Valid_2_delay_10_39 <= io_A_Valid_2_delay_9_40;
    io_A_Valid_2_delay_11_38 <= io_A_Valid_2_delay_10_39;
    io_A_Valid_2_delay_12_37 <= io_A_Valid_2_delay_11_38;
    io_A_Valid_2_delay_13_36 <= io_A_Valid_2_delay_12_37;
    io_A_Valid_2_delay_14_35 <= io_A_Valid_2_delay_13_36;
    io_A_Valid_2_delay_15_34 <= io_A_Valid_2_delay_14_35;
    io_A_Valid_2_delay_16_33 <= io_A_Valid_2_delay_15_34;
    io_A_Valid_2_delay_17_32 <= io_A_Valid_2_delay_16_33;
    io_A_Valid_2_delay_18_31 <= io_A_Valid_2_delay_17_32;
    io_A_Valid_2_delay_19_30 <= io_A_Valid_2_delay_18_31;
    io_A_Valid_2_delay_20_29 <= io_A_Valid_2_delay_19_30;
    io_A_Valid_2_delay_21_28 <= io_A_Valid_2_delay_20_29;
    io_A_Valid_2_delay_22_27 <= io_A_Valid_2_delay_21_28;
    io_A_Valid_2_delay_23_26 <= io_A_Valid_2_delay_22_27;
    io_A_Valid_2_delay_24_25 <= io_A_Valid_2_delay_23_26;
    io_A_Valid_2_delay_25_24 <= io_A_Valid_2_delay_24_25;
    io_A_Valid_2_delay_26_23 <= io_A_Valid_2_delay_25_24;
    io_A_Valid_2_delay_27_22 <= io_A_Valid_2_delay_26_23;
    io_A_Valid_2_delay_28_21 <= io_A_Valid_2_delay_27_22;
    io_A_Valid_2_delay_29_20 <= io_A_Valid_2_delay_28_21;
    io_A_Valid_2_delay_30_19 <= io_A_Valid_2_delay_29_20;
    io_A_Valid_2_delay_31_18 <= io_A_Valid_2_delay_30_19;
    io_A_Valid_2_delay_32_17 <= io_A_Valid_2_delay_31_18;
    io_A_Valid_2_delay_33_16 <= io_A_Valid_2_delay_32_17;
    io_A_Valid_2_delay_34_15 <= io_A_Valid_2_delay_33_16;
    io_A_Valid_2_delay_35_14 <= io_A_Valid_2_delay_34_15;
    io_A_Valid_2_delay_36_13 <= io_A_Valid_2_delay_35_14;
    io_A_Valid_2_delay_37_12 <= io_A_Valid_2_delay_36_13;
    io_A_Valid_2_delay_38_11 <= io_A_Valid_2_delay_37_12;
    io_A_Valid_2_delay_39_10 <= io_A_Valid_2_delay_38_11;
    io_A_Valid_2_delay_40_9 <= io_A_Valid_2_delay_39_10;
    io_A_Valid_2_delay_41_8 <= io_A_Valid_2_delay_40_9;
    io_A_Valid_2_delay_42_7 <= io_A_Valid_2_delay_41_8;
    io_A_Valid_2_delay_43_6 <= io_A_Valid_2_delay_42_7;
    io_A_Valid_2_delay_44_5 <= io_A_Valid_2_delay_43_6;
    io_A_Valid_2_delay_45_4 <= io_A_Valid_2_delay_44_5;
    io_A_Valid_2_delay_46_3 <= io_A_Valid_2_delay_45_4;
    io_A_Valid_2_delay_47_2 <= io_A_Valid_2_delay_46_3;
    io_A_Valid_2_delay_48_1 <= io_A_Valid_2_delay_47_2;
    io_A_Valid_2_delay_49 <= io_A_Valid_2_delay_48_1;
    io_B_Valid_49_delay_1_1 <= io_B_Valid_49;
    io_B_Valid_49_delay_2 <= io_B_Valid_49_delay_1_1;
    io_A_Valid_2_delay_1_49 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_48 <= io_A_Valid_2_delay_1_49;
    io_A_Valid_2_delay_3_47 <= io_A_Valid_2_delay_2_48;
    io_A_Valid_2_delay_4_46 <= io_A_Valid_2_delay_3_47;
    io_A_Valid_2_delay_5_45 <= io_A_Valid_2_delay_4_46;
    io_A_Valid_2_delay_6_44 <= io_A_Valid_2_delay_5_45;
    io_A_Valid_2_delay_7_43 <= io_A_Valid_2_delay_6_44;
    io_A_Valid_2_delay_8_42 <= io_A_Valid_2_delay_7_43;
    io_A_Valid_2_delay_9_41 <= io_A_Valid_2_delay_8_42;
    io_A_Valid_2_delay_10_40 <= io_A_Valid_2_delay_9_41;
    io_A_Valid_2_delay_11_39 <= io_A_Valid_2_delay_10_40;
    io_A_Valid_2_delay_12_38 <= io_A_Valid_2_delay_11_39;
    io_A_Valid_2_delay_13_37 <= io_A_Valid_2_delay_12_38;
    io_A_Valid_2_delay_14_36 <= io_A_Valid_2_delay_13_37;
    io_A_Valid_2_delay_15_35 <= io_A_Valid_2_delay_14_36;
    io_A_Valid_2_delay_16_34 <= io_A_Valid_2_delay_15_35;
    io_A_Valid_2_delay_17_33 <= io_A_Valid_2_delay_16_34;
    io_A_Valid_2_delay_18_32 <= io_A_Valid_2_delay_17_33;
    io_A_Valid_2_delay_19_31 <= io_A_Valid_2_delay_18_32;
    io_A_Valid_2_delay_20_30 <= io_A_Valid_2_delay_19_31;
    io_A_Valid_2_delay_21_29 <= io_A_Valid_2_delay_20_30;
    io_A_Valid_2_delay_22_28 <= io_A_Valid_2_delay_21_29;
    io_A_Valid_2_delay_23_27 <= io_A_Valid_2_delay_22_28;
    io_A_Valid_2_delay_24_26 <= io_A_Valid_2_delay_23_27;
    io_A_Valid_2_delay_25_25 <= io_A_Valid_2_delay_24_26;
    io_A_Valid_2_delay_26_24 <= io_A_Valid_2_delay_25_25;
    io_A_Valid_2_delay_27_23 <= io_A_Valid_2_delay_26_24;
    io_A_Valid_2_delay_28_22 <= io_A_Valid_2_delay_27_23;
    io_A_Valid_2_delay_29_21 <= io_A_Valid_2_delay_28_22;
    io_A_Valid_2_delay_30_20 <= io_A_Valid_2_delay_29_21;
    io_A_Valid_2_delay_31_19 <= io_A_Valid_2_delay_30_20;
    io_A_Valid_2_delay_32_18 <= io_A_Valid_2_delay_31_19;
    io_A_Valid_2_delay_33_17 <= io_A_Valid_2_delay_32_18;
    io_A_Valid_2_delay_34_16 <= io_A_Valid_2_delay_33_17;
    io_A_Valid_2_delay_35_15 <= io_A_Valid_2_delay_34_16;
    io_A_Valid_2_delay_36_14 <= io_A_Valid_2_delay_35_15;
    io_A_Valid_2_delay_37_13 <= io_A_Valid_2_delay_36_14;
    io_A_Valid_2_delay_38_12 <= io_A_Valid_2_delay_37_13;
    io_A_Valid_2_delay_39_11 <= io_A_Valid_2_delay_38_12;
    io_A_Valid_2_delay_40_10 <= io_A_Valid_2_delay_39_11;
    io_A_Valid_2_delay_41_9 <= io_A_Valid_2_delay_40_10;
    io_A_Valid_2_delay_42_8 <= io_A_Valid_2_delay_41_9;
    io_A_Valid_2_delay_43_7 <= io_A_Valid_2_delay_42_8;
    io_A_Valid_2_delay_44_6 <= io_A_Valid_2_delay_43_7;
    io_A_Valid_2_delay_45_5 <= io_A_Valid_2_delay_44_6;
    io_A_Valid_2_delay_46_4 <= io_A_Valid_2_delay_45_5;
    io_A_Valid_2_delay_47_3 <= io_A_Valid_2_delay_46_4;
    io_A_Valid_2_delay_48_2 <= io_A_Valid_2_delay_47_3;
    io_A_Valid_2_delay_49_1 <= io_A_Valid_2_delay_48_2;
    io_A_Valid_2_delay_50 <= io_A_Valid_2_delay_49_1;
    io_B_Valid_50_delay_1_1 <= io_B_Valid_50;
    io_B_Valid_50_delay_2 <= io_B_Valid_50_delay_1_1;
    io_A_Valid_2_delay_1_50 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_49 <= io_A_Valid_2_delay_1_50;
    io_A_Valid_2_delay_3_48 <= io_A_Valid_2_delay_2_49;
    io_A_Valid_2_delay_4_47 <= io_A_Valid_2_delay_3_48;
    io_A_Valid_2_delay_5_46 <= io_A_Valid_2_delay_4_47;
    io_A_Valid_2_delay_6_45 <= io_A_Valid_2_delay_5_46;
    io_A_Valid_2_delay_7_44 <= io_A_Valid_2_delay_6_45;
    io_A_Valid_2_delay_8_43 <= io_A_Valid_2_delay_7_44;
    io_A_Valid_2_delay_9_42 <= io_A_Valid_2_delay_8_43;
    io_A_Valid_2_delay_10_41 <= io_A_Valid_2_delay_9_42;
    io_A_Valid_2_delay_11_40 <= io_A_Valid_2_delay_10_41;
    io_A_Valid_2_delay_12_39 <= io_A_Valid_2_delay_11_40;
    io_A_Valid_2_delay_13_38 <= io_A_Valid_2_delay_12_39;
    io_A_Valid_2_delay_14_37 <= io_A_Valid_2_delay_13_38;
    io_A_Valid_2_delay_15_36 <= io_A_Valid_2_delay_14_37;
    io_A_Valid_2_delay_16_35 <= io_A_Valid_2_delay_15_36;
    io_A_Valid_2_delay_17_34 <= io_A_Valid_2_delay_16_35;
    io_A_Valid_2_delay_18_33 <= io_A_Valid_2_delay_17_34;
    io_A_Valid_2_delay_19_32 <= io_A_Valid_2_delay_18_33;
    io_A_Valid_2_delay_20_31 <= io_A_Valid_2_delay_19_32;
    io_A_Valid_2_delay_21_30 <= io_A_Valid_2_delay_20_31;
    io_A_Valid_2_delay_22_29 <= io_A_Valid_2_delay_21_30;
    io_A_Valid_2_delay_23_28 <= io_A_Valid_2_delay_22_29;
    io_A_Valid_2_delay_24_27 <= io_A_Valid_2_delay_23_28;
    io_A_Valid_2_delay_25_26 <= io_A_Valid_2_delay_24_27;
    io_A_Valid_2_delay_26_25 <= io_A_Valid_2_delay_25_26;
    io_A_Valid_2_delay_27_24 <= io_A_Valid_2_delay_26_25;
    io_A_Valid_2_delay_28_23 <= io_A_Valid_2_delay_27_24;
    io_A_Valid_2_delay_29_22 <= io_A_Valid_2_delay_28_23;
    io_A_Valid_2_delay_30_21 <= io_A_Valid_2_delay_29_22;
    io_A_Valid_2_delay_31_20 <= io_A_Valid_2_delay_30_21;
    io_A_Valid_2_delay_32_19 <= io_A_Valid_2_delay_31_20;
    io_A_Valid_2_delay_33_18 <= io_A_Valid_2_delay_32_19;
    io_A_Valid_2_delay_34_17 <= io_A_Valid_2_delay_33_18;
    io_A_Valid_2_delay_35_16 <= io_A_Valid_2_delay_34_17;
    io_A_Valid_2_delay_36_15 <= io_A_Valid_2_delay_35_16;
    io_A_Valid_2_delay_37_14 <= io_A_Valid_2_delay_36_15;
    io_A_Valid_2_delay_38_13 <= io_A_Valid_2_delay_37_14;
    io_A_Valid_2_delay_39_12 <= io_A_Valid_2_delay_38_13;
    io_A_Valid_2_delay_40_11 <= io_A_Valid_2_delay_39_12;
    io_A_Valid_2_delay_41_10 <= io_A_Valid_2_delay_40_11;
    io_A_Valid_2_delay_42_9 <= io_A_Valid_2_delay_41_10;
    io_A_Valid_2_delay_43_8 <= io_A_Valid_2_delay_42_9;
    io_A_Valid_2_delay_44_7 <= io_A_Valid_2_delay_43_8;
    io_A_Valid_2_delay_45_6 <= io_A_Valid_2_delay_44_7;
    io_A_Valid_2_delay_46_5 <= io_A_Valid_2_delay_45_6;
    io_A_Valid_2_delay_47_4 <= io_A_Valid_2_delay_46_5;
    io_A_Valid_2_delay_48_3 <= io_A_Valid_2_delay_47_4;
    io_A_Valid_2_delay_49_2 <= io_A_Valid_2_delay_48_3;
    io_A_Valid_2_delay_50_1 <= io_A_Valid_2_delay_49_2;
    io_A_Valid_2_delay_51 <= io_A_Valid_2_delay_50_1;
    io_B_Valid_51_delay_1_1 <= io_B_Valid_51;
    io_B_Valid_51_delay_2 <= io_B_Valid_51_delay_1_1;
    io_A_Valid_2_delay_1_51 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_50 <= io_A_Valid_2_delay_1_51;
    io_A_Valid_2_delay_3_49 <= io_A_Valid_2_delay_2_50;
    io_A_Valid_2_delay_4_48 <= io_A_Valid_2_delay_3_49;
    io_A_Valid_2_delay_5_47 <= io_A_Valid_2_delay_4_48;
    io_A_Valid_2_delay_6_46 <= io_A_Valid_2_delay_5_47;
    io_A_Valid_2_delay_7_45 <= io_A_Valid_2_delay_6_46;
    io_A_Valid_2_delay_8_44 <= io_A_Valid_2_delay_7_45;
    io_A_Valid_2_delay_9_43 <= io_A_Valid_2_delay_8_44;
    io_A_Valid_2_delay_10_42 <= io_A_Valid_2_delay_9_43;
    io_A_Valid_2_delay_11_41 <= io_A_Valid_2_delay_10_42;
    io_A_Valid_2_delay_12_40 <= io_A_Valid_2_delay_11_41;
    io_A_Valid_2_delay_13_39 <= io_A_Valid_2_delay_12_40;
    io_A_Valid_2_delay_14_38 <= io_A_Valid_2_delay_13_39;
    io_A_Valid_2_delay_15_37 <= io_A_Valid_2_delay_14_38;
    io_A_Valid_2_delay_16_36 <= io_A_Valid_2_delay_15_37;
    io_A_Valid_2_delay_17_35 <= io_A_Valid_2_delay_16_36;
    io_A_Valid_2_delay_18_34 <= io_A_Valid_2_delay_17_35;
    io_A_Valid_2_delay_19_33 <= io_A_Valid_2_delay_18_34;
    io_A_Valid_2_delay_20_32 <= io_A_Valid_2_delay_19_33;
    io_A_Valid_2_delay_21_31 <= io_A_Valid_2_delay_20_32;
    io_A_Valid_2_delay_22_30 <= io_A_Valid_2_delay_21_31;
    io_A_Valid_2_delay_23_29 <= io_A_Valid_2_delay_22_30;
    io_A_Valid_2_delay_24_28 <= io_A_Valid_2_delay_23_29;
    io_A_Valid_2_delay_25_27 <= io_A_Valid_2_delay_24_28;
    io_A_Valid_2_delay_26_26 <= io_A_Valid_2_delay_25_27;
    io_A_Valid_2_delay_27_25 <= io_A_Valid_2_delay_26_26;
    io_A_Valid_2_delay_28_24 <= io_A_Valid_2_delay_27_25;
    io_A_Valid_2_delay_29_23 <= io_A_Valid_2_delay_28_24;
    io_A_Valid_2_delay_30_22 <= io_A_Valid_2_delay_29_23;
    io_A_Valid_2_delay_31_21 <= io_A_Valid_2_delay_30_22;
    io_A_Valid_2_delay_32_20 <= io_A_Valid_2_delay_31_21;
    io_A_Valid_2_delay_33_19 <= io_A_Valid_2_delay_32_20;
    io_A_Valid_2_delay_34_18 <= io_A_Valid_2_delay_33_19;
    io_A_Valid_2_delay_35_17 <= io_A_Valid_2_delay_34_18;
    io_A_Valid_2_delay_36_16 <= io_A_Valid_2_delay_35_17;
    io_A_Valid_2_delay_37_15 <= io_A_Valid_2_delay_36_16;
    io_A_Valid_2_delay_38_14 <= io_A_Valid_2_delay_37_15;
    io_A_Valid_2_delay_39_13 <= io_A_Valid_2_delay_38_14;
    io_A_Valid_2_delay_40_12 <= io_A_Valid_2_delay_39_13;
    io_A_Valid_2_delay_41_11 <= io_A_Valid_2_delay_40_12;
    io_A_Valid_2_delay_42_10 <= io_A_Valid_2_delay_41_11;
    io_A_Valid_2_delay_43_9 <= io_A_Valid_2_delay_42_10;
    io_A_Valid_2_delay_44_8 <= io_A_Valid_2_delay_43_9;
    io_A_Valid_2_delay_45_7 <= io_A_Valid_2_delay_44_8;
    io_A_Valid_2_delay_46_6 <= io_A_Valid_2_delay_45_7;
    io_A_Valid_2_delay_47_5 <= io_A_Valid_2_delay_46_6;
    io_A_Valid_2_delay_48_4 <= io_A_Valid_2_delay_47_5;
    io_A_Valid_2_delay_49_3 <= io_A_Valid_2_delay_48_4;
    io_A_Valid_2_delay_50_2 <= io_A_Valid_2_delay_49_3;
    io_A_Valid_2_delay_51_1 <= io_A_Valid_2_delay_50_2;
    io_A_Valid_2_delay_52 <= io_A_Valid_2_delay_51_1;
    io_B_Valid_52_delay_1_1 <= io_B_Valid_52;
    io_B_Valid_52_delay_2 <= io_B_Valid_52_delay_1_1;
    io_A_Valid_2_delay_1_52 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_51 <= io_A_Valid_2_delay_1_52;
    io_A_Valid_2_delay_3_50 <= io_A_Valid_2_delay_2_51;
    io_A_Valid_2_delay_4_49 <= io_A_Valid_2_delay_3_50;
    io_A_Valid_2_delay_5_48 <= io_A_Valid_2_delay_4_49;
    io_A_Valid_2_delay_6_47 <= io_A_Valid_2_delay_5_48;
    io_A_Valid_2_delay_7_46 <= io_A_Valid_2_delay_6_47;
    io_A_Valid_2_delay_8_45 <= io_A_Valid_2_delay_7_46;
    io_A_Valid_2_delay_9_44 <= io_A_Valid_2_delay_8_45;
    io_A_Valid_2_delay_10_43 <= io_A_Valid_2_delay_9_44;
    io_A_Valid_2_delay_11_42 <= io_A_Valid_2_delay_10_43;
    io_A_Valid_2_delay_12_41 <= io_A_Valid_2_delay_11_42;
    io_A_Valid_2_delay_13_40 <= io_A_Valid_2_delay_12_41;
    io_A_Valid_2_delay_14_39 <= io_A_Valid_2_delay_13_40;
    io_A_Valid_2_delay_15_38 <= io_A_Valid_2_delay_14_39;
    io_A_Valid_2_delay_16_37 <= io_A_Valid_2_delay_15_38;
    io_A_Valid_2_delay_17_36 <= io_A_Valid_2_delay_16_37;
    io_A_Valid_2_delay_18_35 <= io_A_Valid_2_delay_17_36;
    io_A_Valid_2_delay_19_34 <= io_A_Valid_2_delay_18_35;
    io_A_Valid_2_delay_20_33 <= io_A_Valid_2_delay_19_34;
    io_A_Valid_2_delay_21_32 <= io_A_Valid_2_delay_20_33;
    io_A_Valid_2_delay_22_31 <= io_A_Valid_2_delay_21_32;
    io_A_Valid_2_delay_23_30 <= io_A_Valid_2_delay_22_31;
    io_A_Valid_2_delay_24_29 <= io_A_Valid_2_delay_23_30;
    io_A_Valid_2_delay_25_28 <= io_A_Valid_2_delay_24_29;
    io_A_Valid_2_delay_26_27 <= io_A_Valid_2_delay_25_28;
    io_A_Valid_2_delay_27_26 <= io_A_Valid_2_delay_26_27;
    io_A_Valid_2_delay_28_25 <= io_A_Valid_2_delay_27_26;
    io_A_Valid_2_delay_29_24 <= io_A_Valid_2_delay_28_25;
    io_A_Valid_2_delay_30_23 <= io_A_Valid_2_delay_29_24;
    io_A_Valid_2_delay_31_22 <= io_A_Valid_2_delay_30_23;
    io_A_Valid_2_delay_32_21 <= io_A_Valid_2_delay_31_22;
    io_A_Valid_2_delay_33_20 <= io_A_Valid_2_delay_32_21;
    io_A_Valid_2_delay_34_19 <= io_A_Valid_2_delay_33_20;
    io_A_Valid_2_delay_35_18 <= io_A_Valid_2_delay_34_19;
    io_A_Valid_2_delay_36_17 <= io_A_Valid_2_delay_35_18;
    io_A_Valid_2_delay_37_16 <= io_A_Valid_2_delay_36_17;
    io_A_Valid_2_delay_38_15 <= io_A_Valid_2_delay_37_16;
    io_A_Valid_2_delay_39_14 <= io_A_Valid_2_delay_38_15;
    io_A_Valid_2_delay_40_13 <= io_A_Valid_2_delay_39_14;
    io_A_Valid_2_delay_41_12 <= io_A_Valid_2_delay_40_13;
    io_A_Valid_2_delay_42_11 <= io_A_Valid_2_delay_41_12;
    io_A_Valid_2_delay_43_10 <= io_A_Valid_2_delay_42_11;
    io_A_Valid_2_delay_44_9 <= io_A_Valid_2_delay_43_10;
    io_A_Valid_2_delay_45_8 <= io_A_Valid_2_delay_44_9;
    io_A_Valid_2_delay_46_7 <= io_A_Valid_2_delay_45_8;
    io_A_Valid_2_delay_47_6 <= io_A_Valid_2_delay_46_7;
    io_A_Valid_2_delay_48_5 <= io_A_Valid_2_delay_47_6;
    io_A_Valid_2_delay_49_4 <= io_A_Valid_2_delay_48_5;
    io_A_Valid_2_delay_50_3 <= io_A_Valid_2_delay_49_4;
    io_A_Valid_2_delay_51_2 <= io_A_Valid_2_delay_50_3;
    io_A_Valid_2_delay_52_1 <= io_A_Valid_2_delay_51_2;
    io_A_Valid_2_delay_53 <= io_A_Valid_2_delay_52_1;
    io_B_Valid_53_delay_1_1 <= io_B_Valid_53;
    io_B_Valid_53_delay_2 <= io_B_Valid_53_delay_1_1;
    io_A_Valid_2_delay_1_53 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_52 <= io_A_Valid_2_delay_1_53;
    io_A_Valid_2_delay_3_51 <= io_A_Valid_2_delay_2_52;
    io_A_Valid_2_delay_4_50 <= io_A_Valid_2_delay_3_51;
    io_A_Valid_2_delay_5_49 <= io_A_Valid_2_delay_4_50;
    io_A_Valid_2_delay_6_48 <= io_A_Valid_2_delay_5_49;
    io_A_Valid_2_delay_7_47 <= io_A_Valid_2_delay_6_48;
    io_A_Valid_2_delay_8_46 <= io_A_Valid_2_delay_7_47;
    io_A_Valid_2_delay_9_45 <= io_A_Valid_2_delay_8_46;
    io_A_Valid_2_delay_10_44 <= io_A_Valid_2_delay_9_45;
    io_A_Valid_2_delay_11_43 <= io_A_Valid_2_delay_10_44;
    io_A_Valid_2_delay_12_42 <= io_A_Valid_2_delay_11_43;
    io_A_Valid_2_delay_13_41 <= io_A_Valid_2_delay_12_42;
    io_A_Valid_2_delay_14_40 <= io_A_Valid_2_delay_13_41;
    io_A_Valid_2_delay_15_39 <= io_A_Valid_2_delay_14_40;
    io_A_Valid_2_delay_16_38 <= io_A_Valid_2_delay_15_39;
    io_A_Valid_2_delay_17_37 <= io_A_Valid_2_delay_16_38;
    io_A_Valid_2_delay_18_36 <= io_A_Valid_2_delay_17_37;
    io_A_Valid_2_delay_19_35 <= io_A_Valid_2_delay_18_36;
    io_A_Valid_2_delay_20_34 <= io_A_Valid_2_delay_19_35;
    io_A_Valid_2_delay_21_33 <= io_A_Valid_2_delay_20_34;
    io_A_Valid_2_delay_22_32 <= io_A_Valid_2_delay_21_33;
    io_A_Valid_2_delay_23_31 <= io_A_Valid_2_delay_22_32;
    io_A_Valid_2_delay_24_30 <= io_A_Valid_2_delay_23_31;
    io_A_Valid_2_delay_25_29 <= io_A_Valid_2_delay_24_30;
    io_A_Valid_2_delay_26_28 <= io_A_Valid_2_delay_25_29;
    io_A_Valid_2_delay_27_27 <= io_A_Valid_2_delay_26_28;
    io_A_Valid_2_delay_28_26 <= io_A_Valid_2_delay_27_27;
    io_A_Valid_2_delay_29_25 <= io_A_Valid_2_delay_28_26;
    io_A_Valid_2_delay_30_24 <= io_A_Valid_2_delay_29_25;
    io_A_Valid_2_delay_31_23 <= io_A_Valid_2_delay_30_24;
    io_A_Valid_2_delay_32_22 <= io_A_Valid_2_delay_31_23;
    io_A_Valid_2_delay_33_21 <= io_A_Valid_2_delay_32_22;
    io_A_Valid_2_delay_34_20 <= io_A_Valid_2_delay_33_21;
    io_A_Valid_2_delay_35_19 <= io_A_Valid_2_delay_34_20;
    io_A_Valid_2_delay_36_18 <= io_A_Valid_2_delay_35_19;
    io_A_Valid_2_delay_37_17 <= io_A_Valid_2_delay_36_18;
    io_A_Valid_2_delay_38_16 <= io_A_Valid_2_delay_37_17;
    io_A_Valid_2_delay_39_15 <= io_A_Valid_2_delay_38_16;
    io_A_Valid_2_delay_40_14 <= io_A_Valid_2_delay_39_15;
    io_A_Valid_2_delay_41_13 <= io_A_Valid_2_delay_40_14;
    io_A_Valid_2_delay_42_12 <= io_A_Valid_2_delay_41_13;
    io_A_Valid_2_delay_43_11 <= io_A_Valid_2_delay_42_12;
    io_A_Valid_2_delay_44_10 <= io_A_Valid_2_delay_43_11;
    io_A_Valid_2_delay_45_9 <= io_A_Valid_2_delay_44_10;
    io_A_Valid_2_delay_46_8 <= io_A_Valid_2_delay_45_9;
    io_A_Valid_2_delay_47_7 <= io_A_Valid_2_delay_46_8;
    io_A_Valid_2_delay_48_6 <= io_A_Valid_2_delay_47_7;
    io_A_Valid_2_delay_49_5 <= io_A_Valid_2_delay_48_6;
    io_A_Valid_2_delay_50_4 <= io_A_Valid_2_delay_49_5;
    io_A_Valid_2_delay_51_3 <= io_A_Valid_2_delay_50_4;
    io_A_Valid_2_delay_52_2 <= io_A_Valid_2_delay_51_3;
    io_A_Valid_2_delay_53_1 <= io_A_Valid_2_delay_52_2;
    io_A_Valid_2_delay_54 <= io_A_Valid_2_delay_53_1;
    io_B_Valid_54_delay_1_1 <= io_B_Valid_54;
    io_B_Valid_54_delay_2 <= io_B_Valid_54_delay_1_1;
    io_A_Valid_2_delay_1_54 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_53 <= io_A_Valid_2_delay_1_54;
    io_A_Valid_2_delay_3_52 <= io_A_Valid_2_delay_2_53;
    io_A_Valid_2_delay_4_51 <= io_A_Valid_2_delay_3_52;
    io_A_Valid_2_delay_5_50 <= io_A_Valid_2_delay_4_51;
    io_A_Valid_2_delay_6_49 <= io_A_Valid_2_delay_5_50;
    io_A_Valid_2_delay_7_48 <= io_A_Valid_2_delay_6_49;
    io_A_Valid_2_delay_8_47 <= io_A_Valid_2_delay_7_48;
    io_A_Valid_2_delay_9_46 <= io_A_Valid_2_delay_8_47;
    io_A_Valid_2_delay_10_45 <= io_A_Valid_2_delay_9_46;
    io_A_Valid_2_delay_11_44 <= io_A_Valid_2_delay_10_45;
    io_A_Valid_2_delay_12_43 <= io_A_Valid_2_delay_11_44;
    io_A_Valid_2_delay_13_42 <= io_A_Valid_2_delay_12_43;
    io_A_Valid_2_delay_14_41 <= io_A_Valid_2_delay_13_42;
    io_A_Valid_2_delay_15_40 <= io_A_Valid_2_delay_14_41;
    io_A_Valid_2_delay_16_39 <= io_A_Valid_2_delay_15_40;
    io_A_Valid_2_delay_17_38 <= io_A_Valid_2_delay_16_39;
    io_A_Valid_2_delay_18_37 <= io_A_Valid_2_delay_17_38;
    io_A_Valid_2_delay_19_36 <= io_A_Valid_2_delay_18_37;
    io_A_Valid_2_delay_20_35 <= io_A_Valid_2_delay_19_36;
    io_A_Valid_2_delay_21_34 <= io_A_Valid_2_delay_20_35;
    io_A_Valid_2_delay_22_33 <= io_A_Valid_2_delay_21_34;
    io_A_Valid_2_delay_23_32 <= io_A_Valid_2_delay_22_33;
    io_A_Valid_2_delay_24_31 <= io_A_Valid_2_delay_23_32;
    io_A_Valid_2_delay_25_30 <= io_A_Valid_2_delay_24_31;
    io_A_Valid_2_delay_26_29 <= io_A_Valid_2_delay_25_30;
    io_A_Valid_2_delay_27_28 <= io_A_Valid_2_delay_26_29;
    io_A_Valid_2_delay_28_27 <= io_A_Valid_2_delay_27_28;
    io_A_Valid_2_delay_29_26 <= io_A_Valid_2_delay_28_27;
    io_A_Valid_2_delay_30_25 <= io_A_Valid_2_delay_29_26;
    io_A_Valid_2_delay_31_24 <= io_A_Valid_2_delay_30_25;
    io_A_Valid_2_delay_32_23 <= io_A_Valid_2_delay_31_24;
    io_A_Valid_2_delay_33_22 <= io_A_Valid_2_delay_32_23;
    io_A_Valid_2_delay_34_21 <= io_A_Valid_2_delay_33_22;
    io_A_Valid_2_delay_35_20 <= io_A_Valid_2_delay_34_21;
    io_A_Valid_2_delay_36_19 <= io_A_Valid_2_delay_35_20;
    io_A_Valid_2_delay_37_18 <= io_A_Valid_2_delay_36_19;
    io_A_Valid_2_delay_38_17 <= io_A_Valid_2_delay_37_18;
    io_A_Valid_2_delay_39_16 <= io_A_Valid_2_delay_38_17;
    io_A_Valid_2_delay_40_15 <= io_A_Valid_2_delay_39_16;
    io_A_Valid_2_delay_41_14 <= io_A_Valid_2_delay_40_15;
    io_A_Valid_2_delay_42_13 <= io_A_Valid_2_delay_41_14;
    io_A_Valid_2_delay_43_12 <= io_A_Valid_2_delay_42_13;
    io_A_Valid_2_delay_44_11 <= io_A_Valid_2_delay_43_12;
    io_A_Valid_2_delay_45_10 <= io_A_Valid_2_delay_44_11;
    io_A_Valid_2_delay_46_9 <= io_A_Valid_2_delay_45_10;
    io_A_Valid_2_delay_47_8 <= io_A_Valid_2_delay_46_9;
    io_A_Valid_2_delay_48_7 <= io_A_Valid_2_delay_47_8;
    io_A_Valid_2_delay_49_6 <= io_A_Valid_2_delay_48_7;
    io_A_Valid_2_delay_50_5 <= io_A_Valid_2_delay_49_6;
    io_A_Valid_2_delay_51_4 <= io_A_Valid_2_delay_50_5;
    io_A_Valid_2_delay_52_3 <= io_A_Valid_2_delay_51_4;
    io_A_Valid_2_delay_53_2 <= io_A_Valid_2_delay_52_3;
    io_A_Valid_2_delay_54_1 <= io_A_Valid_2_delay_53_2;
    io_A_Valid_2_delay_55 <= io_A_Valid_2_delay_54_1;
    io_B_Valid_55_delay_1_1 <= io_B_Valid_55;
    io_B_Valid_55_delay_2 <= io_B_Valid_55_delay_1_1;
    io_A_Valid_2_delay_1_55 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_54 <= io_A_Valid_2_delay_1_55;
    io_A_Valid_2_delay_3_53 <= io_A_Valid_2_delay_2_54;
    io_A_Valid_2_delay_4_52 <= io_A_Valid_2_delay_3_53;
    io_A_Valid_2_delay_5_51 <= io_A_Valid_2_delay_4_52;
    io_A_Valid_2_delay_6_50 <= io_A_Valid_2_delay_5_51;
    io_A_Valid_2_delay_7_49 <= io_A_Valid_2_delay_6_50;
    io_A_Valid_2_delay_8_48 <= io_A_Valid_2_delay_7_49;
    io_A_Valid_2_delay_9_47 <= io_A_Valid_2_delay_8_48;
    io_A_Valid_2_delay_10_46 <= io_A_Valid_2_delay_9_47;
    io_A_Valid_2_delay_11_45 <= io_A_Valid_2_delay_10_46;
    io_A_Valid_2_delay_12_44 <= io_A_Valid_2_delay_11_45;
    io_A_Valid_2_delay_13_43 <= io_A_Valid_2_delay_12_44;
    io_A_Valid_2_delay_14_42 <= io_A_Valid_2_delay_13_43;
    io_A_Valid_2_delay_15_41 <= io_A_Valid_2_delay_14_42;
    io_A_Valid_2_delay_16_40 <= io_A_Valid_2_delay_15_41;
    io_A_Valid_2_delay_17_39 <= io_A_Valid_2_delay_16_40;
    io_A_Valid_2_delay_18_38 <= io_A_Valid_2_delay_17_39;
    io_A_Valid_2_delay_19_37 <= io_A_Valid_2_delay_18_38;
    io_A_Valid_2_delay_20_36 <= io_A_Valid_2_delay_19_37;
    io_A_Valid_2_delay_21_35 <= io_A_Valid_2_delay_20_36;
    io_A_Valid_2_delay_22_34 <= io_A_Valid_2_delay_21_35;
    io_A_Valid_2_delay_23_33 <= io_A_Valid_2_delay_22_34;
    io_A_Valid_2_delay_24_32 <= io_A_Valid_2_delay_23_33;
    io_A_Valid_2_delay_25_31 <= io_A_Valid_2_delay_24_32;
    io_A_Valid_2_delay_26_30 <= io_A_Valid_2_delay_25_31;
    io_A_Valid_2_delay_27_29 <= io_A_Valid_2_delay_26_30;
    io_A_Valid_2_delay_28_28 <= io_A_Valid_2_delay_27_29;
    io_A_Valid_2_delay_29_27 <= io_A_Valid_2_delay_28_28;
    io_A_Valid_2_delay_30_26 <= io_A_Valid_2_delay_29_27;
    io_A_Valid_2_delay_31_25 <= io_A_Valid_2_delay_30_26;
    io_A_Valid_2_delay_32_24 <= io_A_Valid_2_delay_31_25;
    io_A_Valid_2_delay_33_23 <= io_A_Valid_2_delay_32_24;
    io_A_Valid_2_delay_34_22 <= io_A_Valid_2_delay_33_23;
    io_A_Valid_2_delay_35_21 <= io_A_Valid_2_delay_34_22;
    io_A_Valid_2_delay_36_20 <= io_A_Valid_2_delay_35_21;
    io_A_Valid_2_delay_37_19 <= io_A_Valid_2_delay_36_20;
    io_A_Valid_2_delay_38_18 <= io_A_Valid_2_delay_37_19;
    io_A_Valid_2_delay_39_17 <= io_A_Valid_2_delay_38_18;
    io_A_Valid_2_delay_40_16 <= io_A_Valid_2_delay_39_17;
    io_A_Valid_2_delay_41_15 <= io_A_Valid_2_delay_40_16;
    io_A_Valid_2_delay_42_14 <= io_A_Valid_2_delay_41_15;
    io_A_Valid_2_delay_43_13 <= io_A_Valid_2_delay_42_14;
    io_A_Valid_2_delay_44_12 <= io_A_Valid_2_delay_43_13;
    io_A_Valid_2_delay_45_11 <= io_A_Valid_2_delay_44_12;
    io_A_Valid_2_delay_46_10 <= io_A_Valid_2_delay_45_11;
    io_A_Valid_2_delay_47_9 <= io_A_Valid_2_delay_46_10;
    io_A_Valid_2_delay_48_8 <= io_A_Valid_2_delay_47_9;
    io_A_Valid_2_delay_49_7 <= io_A_Valid_2_delay_48_8;
    io_A_Valid_2_delay_50_6 <= io_A_Valid_2_delay_49_7;
    io_A_Valid_2_delay_51_5 <= io_A_Valid_2_delay_50_6;
    io_A_Valid_2_delay_52_4 <= io_A_Valid_2_delay_51_5;
    io_A_Valid_2_delay_53_3 <= io_A_Valid_2_delay_52_4;
    io_A_Valid_2_delay_54_2 <= io_A_Valid_2_delay_53_3;
    io_A_Valid_2_delay_55_1 <= io_A_Valid_2_delay_54_2;
    io_A_Valid_2_delay_56 <= io_A_Valid_2_delay_55_1;
    io_B_Valid_56_delay_1_1 <= io_B_Valid_56;
    io_B_Valid_56_delay_2 <= io_B_Valid_56_delay_1_1;
    io_A_Valid_2_delay_1_56 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_55 <= io_A_Valid_2_delay_1_56;
    io_A_Valid_2_delay_3_54 <= io_A_Valid_2_delay_2_55;
    io_A_Valid_2_delay_4_53 <= io_A_Valid_2_delay_3_54;
    io_A_Valid_2_delay_5_52 <= io_A_Valid_2_delay_4_53;
    io_A_Valid_2_delay_6_51 <= io_A_Valid_2_delay_5_52;
    io_A_Valid_2_delay_7_50 <= io_A_Valid_2_delay_6_51;
    io_A_Valid_2_delay_8_49 <= io_A_Valid_2_delay_7_50;
    io_A_Valid_2_delay_9_48 <= io_A_Valid_2_delay_8_49;
    io_A_Valid_2_delay_10_47 <= io_A_Valid_2_delay_9_48;
    io_A_Valid_2_delay_11_46 <= io_A_Valid_2_delay_10_47;
    io_A_Valid_2_delay_12_45 <= io_A_Valid_2_delay_11_46;
    io_A_Valid_2_delay_13_44 <= io_A_Valid_2_delay_12_45;
    io_A_Valid_2_delay_14_43 <= io_A_Valid_2_delay_13_44;
    io_A_Valid_2_delay_15_42 <= io_A_Valid_2_delay_14_43;
    io_A_Valid_2_delay_16_41 <= io_A_Valid_2_delay_15_42;
    io_A_Valid_2_delay_17_40 <= io_A_Valid_2_delay_16_41;
    io_A_Valid_2_delay_18_39 <= io_A_Valid_2_delay_17_40;
    io_A_Valid_2_delay_19_38 <= io_A_Valid_2_delay_18_39;
    io_A_Valid_2_delay_20_37 <= io_A_Valid_2_delay_19_38;
    io_A_Valid_2_delay_21_36 <= io_A_Valid_2_delay_20_37;
    io_A_Valid_2_delay_22_35 <= io_A_Valid_2_delay_21_36;
    io_A_Valid_2_delay_23_34 <= io_A_Valid_2_delay_22_35;
    io_A_Valid_2_delay_24_33 <= io_A_Valid_2_delay_23_34;
    io_A_Valid_2_delay_25_32 <= io_A_Valid_2_delay_24_33;
    io_A_Valid_2_delay_26_31 <= io_A_Valid_2_delay_25_32;
    io_A_Valid_2_delay_27_30 <= io_A_Valid_2_delay_26_31;
    io_A_Valid_2_delay_28_29 <= io_A_Valid_2_delay_27_30;
    io_A_Valid_2_delay_29_28 <= io_A_Valid_2_delay_28_29;
    io_A_Valid_2_delay_30_27 <= io_A_Valid_2_delay_29_28;
    io_A_Valid_2_delay_31_26 <= io_A_Valid_2_delay_30_27;
    io_A_Valid_2_delay_32_25 <= io_A_Valid_2_delay_31_26;
    io_A_Valid_2_delay_33_24 <= io_A_Valid_2_delay_32_25;
    io_A_Valid_2_delay_34_23 <= io_A_Valid_2_delay_33_24;
    io_A_Valid_2_delay_35_22 <= io_A_Valid_2_delay_34_23;
    io_A_Valid_2_delay_36_21 <= io_A_Valid_2_delay_35_22;
    io_A_Valid_2_delay_37_20 <= io_A_Valid_2_delay_36_21;
    io_A_Valid_2_delay_38_19 <= io_A_Valid_2_delay_37_20;
    io_A_Valid_2_delay_39_18 <= io_A_Valid_2_delay_38_19;
    io_A_Valid_2_delay_40_17 <= io_A_Valid_2_delay_39_18;
    io_A_Valid_2_delay_41_16 <= io_A_Valid_2_delay_40_17;
    io_A_Valid_2_delay_42_15 <= io_A_Valid_2_delay_41_16;
    io_A_Valid_2_delay_43_14 <= io_A_Valid_2_delay_42_15;
    io_A_Valid_2_delay_44_13 <= io_A_Valid_2_delay_43_14;
    io_A_Valid_2_delay_45_12 <= io_A_Valid_2_delay_44_13;
    io_A_Valid_2_delay_46_11 <= io_A_Valid_2_delay_45_12;
    io_A_Valid_2_delay_47_10 <= io_A_Valid_2_delay_46_11;
    io_A_Valid_2_delay_48_9 <= io_A_Valid_2_delay_47_10;
    io_A_Valid_2_delay_49_8 <= io_A_Valid_2_delay_48_9;
    io_A_Valid_2_delay_50_7 <= io_A_Valid_2_delay_49_8;
    io_A_Valid_2_delay_51_6 <= io_A_Valid_2_delay_50_7;
    io_A_Valid_2_delay_52_5 <= io_A_Valid_2_delay_51_6;
    io_A_Valid_2_delay_53_4 <= io_A_Valid_2_delay_52_5;
    io_A_Valid_2_delay_54_3 <= io_A_Valid_2_delay_53_4;
    io_A_Valid_2_delay_55_2 <= io_A_Valid_2_delay_54_3;
    io_A_Valid_2_delay_56_1 <= io_A_Valid_2_delay_55_2;
    io_A_Valid_2_delay_57 <= io_A_Valid_2_delay_56_1;
    io_B_Valid_57_delay_1_1 <= io_B_Valid_57;
    io_B_Valid_57_delay_2 <= io_B_Valid_57_delay_1_1;
    io_A_Valid_2_delay_1_57 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_56 <= io_A_Valid_2_delay_1_57;
    io_A_Valid_2_delay_3_55 <= io_A_Valid_2_delay_2_56;
    io_A_Valid_2_delay_4_54 <= io_A_Valid_2_delay_3_55;
    io_A_Valid_2_delay_5_53 <= io_A_Valid_2_delay_4_54;
    io_A_Valid_2_delay_6_52 <= io_A_Valid_2_delay_5_53;
    io_A_Valid_2_delay_7_51 <= io_A_Valid_2_delay_6_52;
    io_A_Valid_2_delay_8_50 <= io_A_Valid_2_delay_7_51;
    io_A_Valid_2_delay_9_49 <= io_A_Valid_2_delay_8_50;
    io_A_Valid_2_delay_10_48 <= io_A_Valid_2_delay_9_49;
    io_A_Valid_2_delay_11_47 <= io_A_Valid_2_delay_10_48;
    io_A_Valid_2_delay_12_46 <= io_A_Valid_2_delay_11_47;
    io_A_Valid_2_delay_13_45 <= io_A_Valid_2_delay_12_46;
    io_A_Valid_2_delay_14_44 <= io_A_Valid_2_delay_13_45;
    io_A_Valid_2_delay_15_43 <= io_A_Valid_2_delay_14_44;
    io_A_Valid_2_delay_16_42 <= io_A_Valid_2_delay_15_43;
    io_A_Valid_2_delay_17_41 <= io_A_Valid_2_delay_16_42;
    io_A_Valid_2_delay_18_40 <= io_A_Valid_2_delay_17_41;
    io_A_Valid_2_delay_19_39 <= io_A_Valid_2_delay_18_40;
    io_A_Valid_2_delay_20_38 <= io_A_Valid_2_delay_19_39;
    io_A_Valid_2_delay_21_37 <= io_A_Valid_2_delay_20_38;
    io_A_Valid_2_delay_22_36 <= io_A_Valid_2_delay_21_37;
    io_A_Valid_2_delay_23_35 <= io_A_Valid_2_delay_22_36;
    io_A_Valid_2_delay_24_34 <= io_A_Valid_2_delay_23_35;
    io_A_Valid_2_delay_25_33 <= io_A_Valid_2_delay_24_34;
    io_A_Valid_2_delay_26_32 <= io_A_Valid_2_delay_25_33;
    io_A_Valid_2_delay_27_31 <= io_A_Valid_2_delay_26_32;
    io_A_Valid_2_delay_28_30 <= io_A_Valid_2_delay_27_31;
    io_A_Valid_2_delay_29_29 <= io_A_Valid_2_delay_28_30;
    io_A_Valid_2_delay_30_28 <= io_A_Valid_2_delay_29_29;
    io_A_Valid_2_delay_31_27 <= io_A_Valid_2_delay_30_28;
    io_A_Valid_2_delay_32_26 <= io_A_Valid_2_delay_31_27;
    io_A_Valid_2_delay_33_25 <= io_A_Valid_2_delay_32_26;
    io_A_Valid_2_delay_34_24 <= io_A_Valid_2_delay_33_25;
    io_A_Valid_2_delay_35_23 <= io_A_Valid_2_delay_34_24;
    io_A_Valid_2_delay_36_22 <= io_A_Valid_2_delay_35_23;
    io_A_Valid_2_delay_37_21 <= io_A_Valid_2_delay_36_22;
    io_A_Valid_2_delay_38_20 <= io_A_Valid_2_delay_37_21;
    io_A_Valid_2_delay_39_19 <= io_A_Valid_2_delay_38_20;
    io_A_Valid_2_delay_40_18 <= io_A_Valid_2_delay_39_19;
    io_A_Valid_2_delay_41_17 <= io_A_Valid_2_delay_40_18;
    io_A_Valid_2_delay_42_16 <= io_A_Valid_2_delay_41_17;
    io_A_Valid_2_delay_43_15 <= io_A_Valid_2_delay_42_16;
    io_A_Valid_2_delay_44_14 <= io_A_Valid_2_delay_43_15;
    io_A_Valid_2_delay_45_13 <= io_A_Valid_2_delay_44_14;
    io_A_Valid_2_delay_46_12 <= io_A_Valid_2_delay_45_13;
    io_A_Valid_2_delay_47_11 <= io_A_Valid_2_delay_46_12;
    io_A_Valid_2_delay_48_10 <= io_A_Valid_2_delay_47_11;
    io_A_Valid_2_delay_49_9 <= io_A_Valid_2_delay_48_10;
    io_A_Valid_2_delay_50_8 <= io_A_Valid_2_delay_49_9;
    io_A_Valid_2_delay_51_7 <= io_A_Valid_2_delay_50_8;
    io_A_Valid_2_delay_52_6 <= io_A_Valid_2_delay_51_7;
    io_A_Valid_2_delay_53_5 <= io_A_Valid_2_delay_52_6;
    io_A_Valid_2_delay_54_4 <= io_A_Valid_2_delay_53_5;
    io_A_Valid_2_delay_55_3 <= io_A_Valid_2_delay_54_4;
    io_A_Valid_2_delay_56_2 <= io_A_Valid_2_delay_55_3;
    io_A_Valid_2_delay_57_1 <= io_A_Valid_2_delay_56_2;
    io_A_Valid_2_delay_58 <= io_A_Valid_2_delay_57_1;
    io_B_Valid_58_delay_1_1 <= io_B_Valid_58;
    io_B_Valid_58_delay_2 <= io_B_Valid_58_delay_1_1;
    io_A_Valid_2_delay_1_58 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_57 <= io_A_Valid_2_delay_1_58;
    io_A_Valid_2_delay_3_56 <= io_A_Valid_2_delay_2_57;
    io_A_Valid_2_delay_4_55 <= io_A_Valid_2_delay_3_56;
    io_A_Valid_2_delay_5_54 <= io_A_Valid_2_delay_4_55;
    io_A_Valid_2_delay_6_53 <= io_A_Valid_2_delay_5_54;
    io_A_Valid_2_delay_7_52 <= io_A_Valid_2_delay_6_53;
    io_A_Valid_2_delay_8_51 <= io_A_Valid_2_delay_7_52;
    io_A_Valid_2_delay_9_50 <= io_A_Valid_2_delay_8_51;
    io_A_Valid_2_delay_10_49 <= io_A_Valid_2_delay_9_50;
    io_A_Valid_2_delay_11_48 <= io_A_Valid_2_delay_10_49;
    io_A_Valid_2_delay_12_47 <= io_A_Valid_2_delay_11_48;
    io_A_Valid_2_delay_13_46 <= io_A_Valid_2_delay_12_47;
    io_A_Valid_2_delay_14_45 <= io_A_Valid_2_delay_13_46;
    io_A_Valid_2_delay_15_44 <= io_A_Valid_2_delay_14_45;
    io_A_Valid_2_delay_16_43 <= io_A_Valid_2_delay_15_44;
    io_A_Valid_2_delay_17_42 <= io_A_Valid_2_delay_16_43;
    io_A_Valid_2_delay_18_41 <= io_A_Valid_2_delay_17_42;
    io_A_Valid_2_delay_19_40 <= io_A_Valid_2_delay_18_41;
    io_A_Valid_2_delay_20_39 <= io_A_Valid_2_delay_19_40;
    io_A_Valid_2_delay_21_38 <= io_A_Valid_2_delay_20_39;
    io_A_Valid_2_delay_22_37 <= io_A_Valid_2_delay_21_38;
    io_A_Valid_2_delay_23_36 <= io_A_Valid_2_delay_22_37;
    io_A_Valid_2_delay_24_35 <= io_A_Valid_2_delay_23_36;
    io_A_Valid_2_delay_25_34 <= io_A_Valid_2_delay_24_35;
    io_A_Valid_2_delay_26_33 <= io_A_Valid_2_delay_25_34;
    io_A_Valid_2_delay_27_32 <= io_A_Valid_2_delay_26_33;
    io_A_Valid_2_delay_28_31 <= io_A_Valid_2_delay_27_32;
    io_A_Valid_2_delay_29_30 <= io_A_Valid_2_delay_28_31;
    io_A_Valid_2_delay_30_29 <= io_A_Valid_2_delay_29_30;
    io_A_Valid_2_delay_31_28 <= io_A_Valid_2_delay_30_29;
    io_A_Valid_2_delay_32_27 <= io_A_Valid_2_delay_31_28;
    io_A_Valid_2_delay_33_26 <= io_A_Valid_2_delay_32_27;
    io_A_Valid_2_delay_34_25 <= io_A_Valid_2_delay_33_26;
    io_A_Valid_2_delay_35_24 <= io_A_Valid_2_delay_34_25;
    io_A_Valid_2_delay_36_23 <= io_A_Valid_2_delay_35_24;
    io_A_Valid_2_delay_37_22 <= io_A_Valid_2_delay_36_23;
    io_A_Valid_2_delay_38_21 <= io_A_Valid_2_delay_37_22;
    io_A_Valid_2_delay_39_20 <= io_A_Valid_2_delay_38_21;
    io_A_Valid_2_delay_40_19 <= io_A_Valid_2_delay_39_20;
    io_A_Valid_2_delay_41_18 <= io_A_Valid_2_delay_40_19;
    io_A_Valid_2_delay_42_17 <= io_A_Valid_2_delay_41_18;
    io_A_Valid_2_delay_43_16 <= io_A_Valid_2_delay_42_17;
    io_A_Valid_2_delay_44_15 <= io_A_Valid_2_delay_43_16;
    io_A_Valid_2_delay_45_14 <= io_A_Valid_2_delay_44_15;
    io_A_Valid_2_delay_46_13 <= io_A_Valid_2_delay_45_14;
    io_A_Valid_2_delay_47_12 <= io_A_Valid_2_delay_46_13;
    io_A_Valid_2_delay_48_11 <= io_A_Valid_2_delay_47_12;
    io_A_Valid_2_delay_49_10 <= io_A_Valid_2_delay_48_11;
    io_A_Valid_2_delay_50_9 <= io_A_Valid_2_delay_49_10;
    io_A_Valid_2_delay_51_8 <= io_A_Valid_2_delay_50_9;
    io_A_Valid_2_delay_52_7 <= io_A_Valid_2_delay_51_8;
    io_A_Valid_2_delay_53_6 <= io_A_Valid_2_delay_52_7;
    io_A_Valid_2_delay_54_5 <= io_A_Valid_2_delay_53_6;
    io_A_Valid_2_delay_55_4 <= io_A_Valid_2_delay_54_5;
    io_A_Valid_2_delay_56_3 <= io_A_Valid_2_delay_55_4;
    io_A_Valid_2_delay_57_2 <= io_A_Valid_2_delay_56_3;
    io_A_Valid_2_delay_58_1 <= io_A_Valid_2_delay_57_2;
    io_A_Valid_2_delay_59 <= io_A_Valid_2_delay_58_1;
    io_B_Valid_59_delay_1_1 <= io_B_Valid_59;
    io_B_Valid_59_delay_2 <= io_B_Valid_59_delay_1_1;
    io_A_Valid_2_delay_1_59 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_58 <= io_A_Valid_2_delay_1_59;
    io_A_Valid_2_delay_3_57 <= io_A_Valid_2_delay_2_58;
    io_A_Valid_2_delay_4_56 <= io_A_Valid_2_delay_3_57;
    io_A_Valid_2_delay_5_55 <= io_A_Valid_2_delay_4_56;
    io_A_Valid_2_delay_6_54 <= io_A_Valid_2_delay_5_55;
    io_A_Valid_2_delay_7_53 <= io_A_Valid_2_delay_6_54;
    io_A_Valid_2_delay_8_52 <= io_A_Valid_2_delay_7_53;
    io_A_Valid_2_delay_9_51 <= io_A_Valid_2_delay_8_52;
    io_A_Valid_2_delay_10_50 <= io_A_Valid_2_delay_9_51;
    io_A_Valid_2_delay_11_49 <= io_A_Valid_2_delay_10_50;
    io_A_Valid_2_delay_12_48 <= io_A_Valid_2_delay_11_49;
    io_A_Valid_2_delay_13_47 <= io_A_Valid_2_delay_12_48;
    io_A_Valid_2_delay_14_46 <= io_A_Valid_2_delay_13_47;
    io_A_Valid_2_delay_15_45 <= io_A_Valid_2_delay_14_46;
    io_A_Valid_2_delay_16_44 <= io_A_Valid_2_delay_15_45;
    io_A_Valid_2_delay_17_43 <= io_A_Valid_2_delay_16_44;
    io_A_Valid_2_delay_18_42 <= io_A_Valid_2_delay_17_43;
    io_A_Valid_2_delay_19_41 <= io_A_Valid_2_delay_18_42;
    io_A_Valid_2_delay_20_40 <= io_A_Valid_2_delay_19_41;
    io_A_Valid_2_delay_21_39 <= io_A_Valid_2_delay_20_40;
    io_A_Valid_2_delay_22_38 <= io_A_Valid_2_delay_21_39;
    io_A_Valid_2_delay_23_37 <= io_A_Valid_2_delay_22_38;
    io_A_Valid_2_delay_24_36 <= io_A_Valid_2_delay_23_37;
    io_A_Valid_2_delay_25_35 <= io_A_Valid_2_delay_24_36;
    io_A_Valid_2_delay_26_34 <= io_A_Valid_2_delay_25_35;
    io_A_Valid_2_delay_27_33 <= io_A_Valid_2_delay_26_34;
    io_A_Valid_2_delay_28_32 <= io_A_Valid_2_delay_27_33;
    io_A_Valid_2_delay_29_31 <= io_A_Valid_2_delay_28_32;
    io_A_Valid_2_delay_30_30 <= io_A_Valid_2_delay_29_31;
    io_A_Valid_2_delay_31_29 <= io_A_Valid_2_delay_30_30;
    io_A_Valid_2_delay_32_28 <= io_A_Valid_2_delay_31_29;
    io_A_Valid_2_delay_33_27 <= io_A_Valid_2_delay_32_28;
    io_A_Valid_2_delay_34_26 <= io_A_Valid_2_delay_33_27;
    io_A_Valid_2_delay_35_25 <= io_A_Valid_2_delay_34_26;
    io_A_Valid_2_delay_36_24 <= io_A_Valid_2_delay_35_25;
    io_A_Valid_2_delay_37_23 <= io_A_Valid_2_delay_36_24;
    io_A_Valid_2_delay_38_22 <= io_A_Valid_2_delay_37_23;
    io_A_Valid_2_delay_39_21 <= io_A_Valid_2_delay_38_22;
    io_A_Valid_2_delay_40_20 <= io_A_Valid_2_delay_39_21;
    io_A_Valid_2_delay_41_19 <= io_A_Valid_2_delay_40_20;
    io_A_Valid_2_delay_42_18 <= io_A_Valid_2_delay_41_19;
    io_A_Valid_2_delay_43_17 <= io_A_Valid_2_delay_42_18;
    io_A_Valid_2_delay_44_16 <= io_A_Valid_2_delay_43_17;
    io_A_Valid_2_delay_45_15 <= io_A_Valid_2_delay_44_16;
    io_A_Valid_2_delay_46_14 <= io_A_Valid_2_delay_45_15;
    io_A_Valid_2_delay_47_13 <= io_A_Valid_2_delay_46_14;
    io_A_Valid_2_delay_48_12 <= io_A_Valid_2_delay_47_13;
    io_A_Valid_2_delay_49_11 <= io_A_Valid_2_delay_48_12;
    io_A_Valid_2_delay_50_10 <= io_A_Valid_2_delay_49_11;
    io_A_Valid_2_delay_51_9 <= io_A_Valid_2_delay_50_10;
    io_A_Valid_2_delay_52_8 <= io_A_Valid_2_delay_51_9;
    io_A_Valid_2_delay_53_7 <= io_A_Valid_2_delay_52_8;
    io_A_Valid_2_delay_54_6 <= io_A_Valid_2_delay_53_7;
    io_A_Valid_2_delay_55_5 <= io_A_Valid_2_delay_54_6;
    io_A_Valid_2_delay_56_4 <= io_A_Valid_2_delay_55_5;
    io_A_Valid_2_delay_57_3 <= io_A_Valid_2_delay_56_4;
    io_A_Valid_2_delay_58_2 <= io_A_Valid_2_delay_57_3;
    io_A_Valid_2_delay_59_1 <= io_A_Valid_2_delay_58_2;
    io_A_Valid_2_delay_60 <= io_A_Valid_2_delay_59_1;
    io_B_Valid_60_delay_1_1 <= io_B_Valid_60;
    io_B_Valid_60_delay_2 <= io_B_Valid_60_delay_1_1;
    io_A_Valid_2_delay_1_60 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_59 <= io_A_Valid_2_delay_1_60;
    io_A_Valid_2_delay_3_58 <= io_A_Valid_2_delay_2_59;
    io_A_Valid_2_delay_4_57 <= io_A_Valid_2_delay_3_58;
    io_A_Valid_2_delay_5_56 <= io_A_Valid_2_delay_4_57;
    io_A_Valid_2_delay_6_55 <= io_A_Valid_2_delay_5_56;
    io_A_Valid_2_delay_7_54 <= io_A_Valid_2_delay_6_55;
    io_A_Valid_2_delay_8_53 <= io_A_Valid_2_delay_7_54;
    io_A_Valid_2_delay_9_52 <= io_A_Valid_2_delay_8_53;
    io_A_Valid_2_delay_10_51 <= io_A_Valid_2_delay_9_52;
    io_A_Valid_2_delay_11_50 <= io_A_Valid_2_delay_10_51;
    io_A_Valid_2_delay_12_49 <= io_A_Valid_2_delay_11_50;
    io_A_Valid_2_delay_13_48 <= io_A_Valid_2_delay_12_49;
    io_A_Valid_2_delay_14_47 <= io_A_Valid_2_delay_13_48;
    io_A_Valid_2_delay_15_46 <= io_A_Valid_2_delay_14_47;
    io_A_Valid_2_delay_16_45 <= io_A_Valid_2_delay_15_46;
    io_A_Valid_2_delay_17_44 <= io_A_Valid_2_delay_16_45;
    io_A_Valid_2_delay_18_43 <= io_A_Valid_2_delay_17_44;
    io_A_Valid_2_delay_19_42 <= io_A_Valid_2_delay_18_43;
    io_A_Valid_2_delay_20_41 <= io_A_Valid_2_delay_19_42;
    io_A_Valid_2_delay_21_40 <= io_A_Valid_2_delay_20_41;
    io_A_Valid_2_delay_22_39 <= io_A_Valid_2_delay_21_40;
    io_A_Valid_2_delay_23_38 <= io_A_Valid_2_delay_22_39;
    io_A_Valid_2_delay_24_37 <= io_A_Valid_2_delay_23_38;
    io_A_Valid_2_delay_25_36 <= io_A_Valid_2_delay_24_37;
    io_A_Valid_2_delay_26_35 <= io_A_Valid_2_delay_25_36;
    io_A_Valid_2_delay_27_34 <= io_A_Valid_2_delay_26_35;
    io_A_Valid_2_delay_28_33 <= io_A_Valid_2_delay_27_34;
    io_A_Valid_2_delay_29_32 <= io_A_Valid_2_delay_28_33;
    io_A_Valid_2_delay_30_31 <= io_A_Valid_2_delay_29_32;
    io_A_Valid_2_delay_31_30 <= io_A_Valid_2_delay_30_31;
    io_A_Valid_2_delay_32_29 <= io_A_Valid_2_delay_31_30;
    io_A_Valid_2_delay_33_28 <= io_A_Valid_2_delay_32_29;
    io_A_Valid_2_delay_34_27 <= io_A_Valid_2_delay_33_28;
    io_A_Valid_2_delay_35_26 <= io_A_Valid_2_delay_34_27;
    io_A_Valid_2_delay_36_25 <= io_A_Valid_2_delay_35_26;
    io_A_Valid_2_delay_37_24 <= io_A_Valid_2_delay_36_25;
    io_A_Valid_2_delay_38_23 <= io_A_Valid_2_delay_37_24;
    io_A_Valid_2_delay_39_22 <= io_A_Valid_2_delay_38_23;
    io_A_Valid_2_delay_40_21 <= io_A_Valid_2_delay_39_22;
    io_A_Valid_2_delay_41_20 <= io_A_Valid_2_delay_40_21;
    io_A_Valid_2_delay_42_19 <= io_A_Valid_2_delay_41_20;
    io_A_Valid_2_delay_43_18 <= io_A_Valid_2_delay_42_19;
    io_A_Valid_2_delay_44_17 <= io_A_Valid_2_delay_43_18;
    io_A_Valid_2_delay_45_16 <= io_A_Valid_2_delay_44_17;
    io_A_Valid_2_delay_46_15 <= io_A_Valid_2_delay_45_16;
    io_A_Valid_2_delay_47_14 <= io_A_Valid_2_delay_46_15;
    io_A_Valid_2_delay_48_13 <= io_A_Valid_2_delay_47_14;
    io_A_Valid_2_delay_49_12 <= io_A_Valid_2_delay_48_13;
    io_A_Valid_2_delay_50_11 <= io_A_Valid_2_delay_49_12;
    io_A_Valid_2_delay_51_10 <= io_A_Valid_2_delay_50_11;
    io_A_Valid_2_delay_52_9 <= io_A_Valid_2_delay_51_10;
    io_A_Valid_2_delay_53_8 <= io_A_Valid_2_delay_52_9;
    io_A_Valid_2_delay_54_7 <= io_A_Valid_2_delay_53_8;
    io_A_Valid_2_delay_55_6 <= io_A_Valid_2_delay_54_7;
    io_A_Valid_2_delay_56_5 <= io_A_Valid_2_delay_55_6;
    io_A_Valid_2_delay_57_4 <= io_A_Valid_2_delay_56_5;
    io_A_Valid_2_delay_58_3 <= io_A_Valid_2_delay_57_4;
    io_A_Valid_2_delay_59_2 <= io_A_Valid_2_delay_58_3;
    io_A_Valid_2_delay_60_1 <= io_A_Valid_2_delay_59_2;
    io_A_Valid_2_delay_61 <= io_A_Valid_2_delay_60_1;
    io_B_Valid_61_delay_1_1 <= io_B_Valid_61;
    io_B_Valid_61_delay_2 <= io_B_Valid_61_delay_1_1;
    io_A_Valid_2_delay_1_61 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_60 <= io_A_Valid_2_delay_1_61;
    io_A_Valid_2_delay_3_59 <= io_A_Valid_2_delay_2_60;
    io_A_Valid_2_delay_4_58 <= io_A_Valid_2_delay_3_59;
    io_A_Valid_2_delay_5_57 <= io_A_Valid_2_delay_4_58;
    io_A_Valid_2_delay_6_56 <= io_A_Valid_2_delay_5_57;
    io_A_Valid_2_delay_7_55 <= io_A_Valid_2_delay_6_56;
    io_A_Valid_2_delay_8_54 <= io_A_Valid_2_delay_7_55;
    io_A_Valid_2_delay_9_53 <= io_A_Valid_2_delay_8_54;
    io_A_Valid_2_delay_10_52 <= io_A_Valid_2_delay_9_53;
    io_A_Valid_2_delay_11_51 <= io_A_Valid_2_delay_10_52;
    io_A_Valid_2_delay_12_50 <= io_A_Valid_2_delay_11_51;
    io_A_Valid_2_delay_13_49 <= io_A_Valid_2_delay_12_50;
    io_A_Valid_2_delay_14_48 <= io_A_Valid_2_delay_13_49;
    io_A_Valid_2_delay_15_47 <= io_A_Valid_2_delay_14_48;
    io_A_Valid_2_delay_16_46 <= io_A_Valid_2_delay_15_47;
    io_A_Valid_2_delay_17_45 <= io_A_Valid_2_delay_16_46;
    io_A_Valid_2_delay_18_44 <= io_A_Valid_2_delay_17_45;
    io_A_Valid_2_delay_19_43 <= io_A_Valid_2_delay_18_44;
    io_A_Valid_2_delay_20_42 <= io_A_Valid_2_delay_19_43;
    io_A_Valid_2_delay_21_41 <= io_A_Valid_2_delay_20_42;
    io_A_Valid_2_delay_22_40 <= io_A_Valid_2_delay_21_41;
    io_A_Valid_2_delay_23_39 <= io_A_Valid_2_delay_22_40;
    io_A_Valid_2_delay_24_38 <= io_A_Valid_2_delay_23_39;
    io_A_Valid_2_delay_25_37 <= io_A_Valid_2_delay_24_38;
    io_A_Valid_2_delay_26_36 <= io_A_Valid_2_delay_25_37;
    io_A_Valid_2_delay_27_35 <= io_A_Valid_2_delay_26_36;
    io_A_Valid_2_delay_28_34 <= io_A_Valid_2_delay_27_35;
    io_A_Valid_2_delay_29_33 <= io_A_Valid_2_delay_28_34;
    io_A_Valid_2_delay_30_32 <= io_A_Valid_2_delay_29_33;
    io_A_Valid_2_delay_31_31 <= io_A_Valid_2_delay_30_32;
    io_A_Valid_2_delay_32_30 <= io_A_Valid_2_delay_31_31;
    io_A_Valid_2_delay_33_29 <= io_A_Valid_2_delay_32_30;
    io_A_Valid_2_delay_34_28 <= io_A_Valid_2_delay_33_29;
    io_A_Valid_2_delay_35_27 <= io_A_Valid_2_delay_34_28;
    io_A_Valid_2_delay_36_26 <= io_A_Valid_2_delay_35_27;
    io_A_Valid_2_delay_37_25 <= io_A_Valid_2_delay_36_26;
    io_A_Valid_2_delay_38_24 <= io_A_Valid_2_delay_37_25;
    io_A_Valid_2_delay_39_23 <= io_A_Valid_2_delay_38_24;
    io_A_Valid_2_delay_40_22 <= io_A_Valid_2_delay_39_23;
    io_A_Valid_2_delay_41_21 <= io_A_Valid_2_delay_40_22;
    io_A_Valid_2_delay_42_20 <= io_A_Valid_2_delay_41_21;
    io_A_Valid_2_delay_43_19 <= io_A_Valid_2_delay_42_20;
    io_A_Valid_2_delay_44_18 <= io_A_Valid_2_delay_43_19;
    io_A_Valid_2_delay_45_17 <= io_A_Valid_2_delay_44_18;
    io_A_Valid_2_delay_46_16 <= io_A_Valid_2_delay_45_17;
    io_A_Valid_2_delay_47_15 <= io_A_Valid_2_delay_46_16;
    io_A_Valid_2_delay_48_14 <= io_A_Valid_2_delay_47_15;
    io_A_Valid_2_delay_49_13 <= io_A_Valid_2_delay_48_14;
    io_A_Valid_2_delay_50_12 <= io_A_Valid_2_delay_49_13;
    io_A_Valid_2_delay_51_11 <= io_A_Valid_2_delay_50_12;
    io_A_Valid_2_delay_52_10 <= io_A_Valid_2_delay_51_11;
    io_A_Valid_2_delay_53_9 <= io_A_Valid_2_delay_52_10;
    io_A_Valid_2_delay_54_8 <= io_A_Valid_2_delay_53_9;
    io_A_Valid_2_delay_55_7 <= io_A_Valid_2_delay_54_8;
    io_A_Valid_2_delay_56_6 <= io_A_Valid_2_delay_55_7;
    io_A_Valid_2_delay_57_5 <= io_A_Valid_2_delay_56_6;
    io_A_Valid_2_delay_58_4 <= io_A_Valid_2_delay_57_5;
    io_A_Valid_2_delay_59_3 <= io_A_Valid_2_delay_58_4;
    io_A_Valid_2_delay_60_2 <= io_A_Valid_2_delay_59_3;
    io_A_Valid_2_delay_61_1 <= io_A_Valid_2_delay_60_2;
    io_A_Valid_2_delay_62 <= io_A_Valid_2_delay_61_1;
    io_B_Valid_62_delay_1_1 <= io_B_Valid_62;
    io_B_Valid_62_delay_2 <= io_B_Valid_62_delay_1_1;
    io_A_Valid_2_delay_1_62 <= io_A_Valid_2;
    io_A_Valid_2_delay_2_61 <= io_A_Valid_2_delay_1_62;
    io_A_Valid_2_delay_3_60 <= io_A_Valid_2_delay_2_61;
    io_A_Valid_2_delay_4_59 <= io_A_Valid_2_delay_3_60;
    io_A_Valid_2_delay_5_58 <= io_A_Valid_2_delay_4_59;
    io_A_Valid_2_delay_6_57 <= io_A_Valid_2_delay_5_58;
    io_A_Valid_2_delay_7_56 <= io_A_Valid_2_delay_6_57;
    io_A_Valid_2_delay_8_55 <= io_A_Valid_2_delay_7_56;
    io_A_Valid_2_delay_9_54 <= io_A_Valid_2_delay_8_55;
    io_A_Valid_2_delay_10_53 <= io_A_Valid_2_delay_9_54;
    io_A_Valid_2_delay_11_52 <= io_A_Valid_2_delay_10_53;
    io_A_Valid_2_delay_12_51 <= io_A_Valid_2_delay_11_52;
    io_A_Valid_2_delay_13_50 <= io_A_Valid_2_delay_12_51;
    io_A_Valid_2_delay_14_49 <= io_A_Valid_2_delay_13_50;
    io_A_Valid_2_delay_15_48 <= io_A_Valid_2_delay_14_49;
    io_A_Valid_2_delay_16_47 <= io_A_Valid_2_delay_15_48;
    io_A_Valid_2_delay_17_46 <= io_A_Valid_2_delay_16_47;
    io_A_Valid_2_delay_18_45 <= io_A_Valid_2_delay_17_46;
    io_A_Valid_2_delay_19_44 <= io_A_Valid_2_delay_18_45;
    io_A_Valid_2_delay_20_43 <= io_A_Valid_2_delay_19_44;
    io_A_Valid_2_delay_21_42 <= io_A_Valid_2_delay_20_43;
    io_A_Valid_2_delay_22_41 <= io_A_Valid_2_delay_21_42;
    io_A_Valid_2_delay_23_40 <= io_A_Valid_2_delay_22_41;
    io_A_Valid_2_delay_24_39 <= io_A_Valid_2_delay_23_40;
    io_A_Valid_2_delay_25_38 <= io_A_Valid_2_delay_24_39;
    io_A_Valid_2_delay_26_37 <= io_A_Valid_2_delay_25_38;
    io_A_Valid_2_delay_27_36 <= io_A_Valid_2_delay_26_37;
    io_A_Valid_2_delay_28_35 <= io_A_Valid_2_delay_27_36;
    io_A_Valid_2_delay_29_34 <= io_A_Valid_2_delay_28_35;
    io_A_Valid_2_delay_30_33 <= io_A_Valid_2_delay_29_34;
    io_A_Valid_2_delay_31_32 <= io_A_Valid_2_delay_30_33;
    io_A_Valid_2_delay_32_31 <= io_A_Valid_2_delay_31_32;
    io_A_Valid_2_delay_33_30 <= io_A_Valid_2_delay_32_31;
    io_A_Valid_2_delay_34_29 <= io_A_Valid_2_delay_33_30;
    io_A_Valid_2_delay_35_28 <= io_A_Valid_2_delay_34_29;
    io_A_Valid_2_delay_36_27 <= io_A_Valid_2_delay_35_28;
    io_A_Valid_2_delay_37_26 <= io_A_Valid_2_delay_36_27;
    io_A_Valid_2_delay_38_25 <= io_A_Valid_2_delay_37_26;
    io_A_Valid_2_delay_39_24 <= io_A_Valid_2_delay_38_25;
    io_A_Valid_2_delay_40_23 <= io_A_Valid_2_delay_39_24;
    io_A_Valid_2_delay_41_22 <= io_A_Valid_2_delay_40_23;
    io_A_Valid_2_delay_42_21 <= io_A_Valid_2_delay_41_22;
    io_A_Valid_2_delay_43_20 <= io_A_Valid_2_delay_42_21;
    io_A_Valid_2_delay_44_19 <= io_A_Valid_2_delay_43_20;
    io_A_Valid_2_delay_45_18 <= io_A_Valid_2_delay_44_19;
    io_A_Valid_2_delay_46_17 <= io_A_Valid_2_delay_45_18;
    io_A_Valid_2_delay_47_16 <= io_A_Valid_2_delay_46_17;
    io_A_Valid_2_delay_48_15 <= io_A_Valid_2_delay_47_16;
    io_A_Valid_2_delay_49_14 <= io_A_Valid_2_delay_48_15;
    io_A_Valid_2_delay_50_13 <= io_A_Valid_2_delay_49_14;
    io_A_Valid_2_delay_51_12 <= io_A_Valid_2_delay_50_13;
    io_A_Valid_2_delay_52_11 <= io_A_Valid_2_delay_51_12;
    io_A_Valid_2_delay_53_10 <= io_A_Valid_2_delay_52_11;
    io_A_Valid_2_delay_54_9 <= io_A_Valid_2_delay_53_10;
    io_A_Valid_2_delay_55_8 <= io_A_Valid_2_delay_54_9;
    io_A_Valid_2_delay_56_7 <= io_A_Valid_2_delay_55_8;
    io_A_Valid_2_delay_57_6 <= io_A_Valid_2_delay_56_7;
    io_A_Valid_2_delay_58_5 <= io_A_Valid_2_delay_57_6;
    io_A_Valid_2_delay_59_4 <= io_A_Valid_2_delay_58_5;
    io_A_Valid_2_delay_60_3 <= io_A_Valid_2_delay_59_4;
    io_A_Valid_2_delay_61_2 <= io_A_Valid_2_delay_60_3;
    io_A_Valid_2_delay_62_1 <= io_A_Valid_2_delay_61_2;
    io_A_Valid_2_delay_63 <= io_A_Valid_2_delay_62_1;
    io_B_Valid_63_delay_1_1 <= io_B_Valid_63;
    io_B_Valid_63_delay_2 <= io_B_Valid_63_delay_1_1;
    io_B_Valid_0_delay_1_2 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_1 <= io_B_Valid_0_delay_1_2;
    io_B_Valid_0_delay_3 <= io_B_Valid_0_delay_2_1;
    io_A_Valid_3_delay_1 <= io_A_Valid_3;
    io_B_Valid_1_delay_1_2 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_1 <= io_B_Valid_1_delay_1_2;
    io_B_Valid_1_delay_3 <= io_B_Valid_1_delay_2_1;
    io_A_Valid_3_delay_1_1 <= io_A_Valid_3;
    io_A_Valid_3_delay_2 <= io_A_Valid_3_delay_1_1;
    io_B_Valid_2_delay_1_2 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_1 <= io_B_Valid_2_delay_1_2;
    io_B_Valid_2_delay_3 <= io_B_Valid_2_delay_2_1;
    io_A_Valid_3_delay_1_2 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_1 <= io_A_Valid_3_delay_1_2;
    io_A_Valid_3_delay_3 <= io_A_Valid_3_delay_2_1;
    io_B_Valid_3_delay_1_2 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_1 <= io_B_Valid_3_delay_1_2;
    io_B_Valid_3_delay_3 <= io_B_Valid_3_delay_2_1;
    io_A_Valid_3_delay_1_3 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_2 <= io_A_Valid_3_delay_1_3;
    io_A_Valid_3_delay_3_1 <= io_A_Valid_3_delay_2_2;
    io_A_Valid_3_delay_4 <= io_A_Valid_3_delay_3_1;
    io_B_Valid_4_delay_1_2 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_1 <= io_B_Valid_4_delay_1_2;
    io_B_Valid_4_delay_3 <= io_B_Valid_4_delay_2_1;
    io_A_Valid_3_delay_1_4 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_3 <= io_A_Valid_3_delay_1_4;
    io_A_Valid_3_delay_3_2 <= io_A_Valid_3_delay_2_3;
    io_A_Valid_3_delay_4_1 <= io_A_Valid_3_delay_3_2;
    io_A_Valid_3_delay_5 <= io_A_Valid_3_delay_4_1;
    io_B_Valid_5_delay_1_2 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_1 <= io_B_Valid_5_delay_1_2;
    io_B_Valid_5_delay_3 <= io_B_Valid_5_delay_2_1;
    io_A_Valid_3_delay_1_5 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_4 <= io_A_Valid_3_delay_1_5;
    io_A_Valid_3_delay_3_3 <= io_A_Valid_3_delay_2_4;
    io_A_Valid_3_delay_4_2 <= io_A_Valid_3_delay_3_3;
    io_A_Valid_3_delay_5_1 <= io_A_Valid_3_delay_4_2;
    io_A_Valid_3_delay_6 <= io_A_Valid_3_delay_5_1;
    io_B_Valid_6_delay_1_2 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_1 <= io_B_Valid_6_delay_1_2;
    io_B_Valid_6_delay_3 <= io_B_Valid_6_delay_2_1;
    io_A_Valid_3_delay_1_6 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_5 <= io_A_Valid_3_delay_1_6;
    io_A_Valid_3_delay_3_4 <= io_A_Valid_3_delay_2_5;
    io_A_Valid_3_delay_4_3 <= io_A_Valid_3_delay_3_4;
    io_A_Valid_3_delay_5_2 <= io_A_Valid_3_delay_4_3;
    io_A_Valid_3_delay_6_1 <= io_A_Valid_3_delay_5_2;
    io_A_Valid_3_delay_7 <= io_A_Valid_3_delay_6_1;
    io_B_Valid_7_delay_1_2 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_1 <= io_B_Valid_7_delay_1_2;
    io_B_Valid_7_delay_3 <= io_B_Valid_7_delay_2_1;
    io_A_Valid_3_delay_1_7 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_6 <= io_A_Valid_3_delay_1_7;
    io_A_Valid_3_delay_3_5 <= io_A_Valid_3_delay_2_6;
    io_A_Valid_3_delay_4_4 <= io_A_Valid_3_delay_3_5;
    io_A_Valid_3_delay_5_3 <= io_A_Valid_3_delay_4_4;
    io_A_Valid_3_delay_6_2 <= io_A_Valid_3_delay_5_3;
    io_A_Valid_3_delay_7_1 <= io_A_Valid_3_delay_6_2;
    io_A_Valid_3_delay_8 <= io_A_Valid_3_delay_7_1;
    io_B_Valid_8_delay_1_2 <= io_B_Valid_8;
    io_B_Valid_8_delay_2_1 <= io_B_Valid_8_delay_1_2;
    io_B_Valid_8_delay_3 <= io_B_Valid_8_delay_2_1;
    io_A_Valid_3_delay_1_8 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_7 <= io_A_Valid_3_delay_1_8;
    io_A_Valid_3_delay_3_6 <= io_A_Valid_3_delay_2_7;
    io_A_Valid_3_delay_4_5 <= io_A_Valid_3_delay_3_6;
    io_A_Valid_3_delay_5_4 <= io_A_Valid_3_delay_4_5;
    io_A_Valid_3_delay_6_3 <= io_A_Valid_3_delay_5_4;
    io_A_Valid_3_delay_7_2 <= io_A_Valid_3_delay_6_3;
    io_A_Valid_3_delay_8_1 <= io_A_Valid_3_delay_7_2;
    io_A_Valid_3_delay_9 <= io_A_Valid_3_delay_8_1;
    io_B_Valid_9_delay_1_2 <= io_B_Valid_9;
    io_B_Valid_9_delay_2_1 <= io_B_Valid_9_delay_1_2;
    io_B_Valid_9_delay_3 <= io_B_Valid_9_delay_2_1;
    io_A_Valid_3_delay_1_9 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_8 <= io_A_Valid_3_delay_1_9;
    io_A_Valid_3_delay_3_7 <= io_A_Valid_3_delay_2_8;
    io_A_Valid_3_delay_4_6 <= io_A_Valid_3_delay_3_7;
    io_A_Valid_3_delay_5_5 <= io_A_Valid_3_delay_4_6;
    io_A_Valid_3_delay_6_4 <= io_A_Valid_3_delay_5_5;
    io_A_Valid_3_delay_7_3 <= io_A_Valid_3_delay_6_4;
    io_A_Valid_3_delay_8_2 <= io_A_Valid_3_delay_7_3;
    io_A_Valid_3_delay_9_1 <= io_A_Valid_3_delay_8_2;
    io_A_Valid_3_delay_10 <= io_A_Valid_3_delay_9_1;
    io_B_Valid_10_delay_1_2 <= io_B_Valid_10;
    io_B_Valid_10_delay_2_1 <= io_B_Valid_10_delay_1_2;
    io_B_Valid_10_delay_3 <= io_B_Valid_10_delay_2_1;
    io_A_Valid_3_delay_1_10 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_9 <= io_A_Valid_3_delay_1_10;
    io_A_Valid_3_delay_3_8 <= io_A_Valid_3_delay_2_9;
    io_A_Valid_3_delay_4_7 <= io_A_Valid_3_delay_3_8;
    io_A_Valid_3_delay_5_6 <= io_A_Valid_3_delay_4_7;
    io_A_Valid_3_delay_6_5 <= io_A_Valid_3_delay_5_6;
    io_A_Valid_3_delay_7_4 <= io_A_Valid_3_delay_6_5;
    io_A_Valid_3_delay_8_3 <= io_A_Valid_3_delay_7_4;
    io_A_Valid_3_delay_9_2 <= io_A_Valid_3_delay_8_3;
    io_A_Valid_3_delay_10_1 <= io_A_Valid_3_delay_9_2;
    io_A_Valid_3_delay_11 <= io_A_Valid_3_delay_10_1;
    io_B_Valid_11_delay_1_2 <= io_B_Valid_11;
    io_B_Valid_11_delay_2_1 <= io_B_Valid_11_delay_1_2;
    io_B_Valid_11_delay_3 <= io_B_Valid_11_delay_2_1;
    io_A_Valid_3_delay_1_11 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_10 <= io_A_Valid_3_delay_1_11;
    io_A_Valid_3_delay_3_9 <= io_A_Valid_3_delay_2_10;
    io_A_Valid_3_delay_4_8 <= io_A_Valid_3_delay_3_9;
    io_A_Valid_3_delay_5_7 <= io_A_Valid_3_delay_4_8;
    io_A_Valid_3_delay_6_6 <= io_A_Valid_3_delay_5_7;
    io_A_Valid_3_delay_7_5 <= io_A_Valid_3_delay_6_6;
    io_A_Valid_3_delay_8_4 <= io_A_Valid_3_delay_7_5;
    io_A_Valid_3_delay_9_3 <= io_A_Valid_3_delay_8_4;
    io_A_Valid_3_delay_10_2 <= io_A_Valid_3_delay_9_3;
    io_A_Valid_3_delay_11_1 <= io_A_Valid_3_delay_10_2;
    io_A_Valid_3_delay_12 <= io_A_Valid_3_delay_11_1;
    io_B_Valid_12_delay_1_2 <= io_B_Valid_12;
    io_B_Valid_12_delay_2_1 <= io_B_Valid_12_delay_1_2;
    io_B_Valid_12_delay_3 <= io_B_Valid_12_delay_2_1;
    io_A_Valid_3_delay_1_12 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_11 <= io_A_Valid_3_delay_1_12;
    io_A_Valid_3_delay_3_10 <= io_A_Valid_3_delay_2_11;
    io_A_Valid_3_delay_4_9 <= io_A_Valid_3_delay_3_10;
    io_A_Valid_3_delay_5_8 <= io_A_Valid_3_delay_4_9;
    io_A_Valid_3_delay_6_7 <= io_A_Valid_3_delay_5_8;
    io_A_Valid_3_delay_7_6 <= io_A_Valid_3_delay_6_7;
    io_A_Valid_3_delay_8_5 <= io_A_Valid_3_delay_7_6;
    io_A_Valid_3_delay_9_4 <= io_A_Valid_3_delay_8_5;
    io_A_Valid_3_delay_10_3 <= io_A_Valid_3_delay_9_4;
    io_A_Valid_3_delay_11_2 <= io_A_Valid_3_delay_10_3;
    io_A_Valid_3_delay_12_1 <= io_A_Valid_3_delay_11_2;
    io_A_Valid_3_delay_13 <= io_A_Valid_3_delay_12_1;
    io_B_Valid_13_delay_1_2 <= io_B_Valid_13;
    io_B_Valid_13_delay_2_1 <= io_B_Valid_13_delay_1_2;
    io_B_Valid_13_delay_3 <= io_B_Valid_13_delay_2_1;
    io_A_Valid_3_delay_1_13 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_12 <= io_A_Valid_3_delay_1_13;
    io_A_Valid_3_delay_3_11 <= io_A_Valid_3_delay_2_12;
    io_A_Valid_3_delay_4_10 <= io_A_Valid_3_delay_3_11;
    io_A_Valid_3_delay_5_9 <= io_A_Valid_3_delay_4_10;
    io_A_Valid_3_delay_6_8 <= io_A_Valid_3_delay_5_9;
    io_A_Valid_3_delay_7_7 <= io_A_Valid_3_delay_6_8;
    io_A_Valid_3_delay_8_6 <= io_A_Valid_3_delay_7_7;
    io_A_Valid_3_delay_9_5 <= io_A_Valid_3_delay_8_6;
    io_A_Valid_3_delay_10_4 <= io_A_Valid_3_delay_9_5;
    io_A_Valid_3_delay_11_3 <= io_A_Valid_3_delay_10_4;
    io_A_Valid_3_delay_12_2 <= io_A_Valid_3_delay_11_3;
    io_A_Valid_3_delay_13_1 <= io_A_Valid_3_delay_12_2;
    io_A_Valid_3_delay_14 <= io_A_Valid_3_delay_13_1;
    io_B_Valid_14_delay_1_2 <= io_B_Valid_14;
    io_B_Valid_14_delay_2_1 <= io_B_Valid_14_delay_1_2;
    io_B_Valid_14_delay_3 <= io_B_Valid_14_delay_2_1;
    io_A_Valid_3_delay_1_14 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_13 <= io_A_Valid_3_delay_1_14;
    io_A_Valid_3_delay_3_12 <= io_A_Valid_3_delay_2_13;
    io_A_Valid_3_delay_4_11 <= io_A_Valid_3_delay_3_12;
    io_A_Valid_3_delay_5_10 <= io_A_Valid_3_delay_4_11;
    io_A_Valid_3_delay_6_9 <= io_A_Valid_3_delay_5_10;
    io_A_Valid_3_delay_7_8 <= io_A_Valid_3_delay_6_9;
    io_A_Valid_3_delay_8_7 <= io_A_Valid_3_delay_7_8;
    io_A_Valid_3_delay_9_6 <= io_A_Valid_3_delay_8_7;
    io_A_Valid_3_delay_10_5 <= io_A_Valid_3_delay_9_6;
    io_A_Valid_3_delay_11_4 <= io_A_Valid_3_delay_10_5;
    io_A_Valid_3_delay_12_3 <= io_A_Valid_3_delay_11_4;
    io_A_Valid_3_delay_13_2 <= io_A_Valid_3_delay_12_3;
    io_A_Valid_3_delay_14_1 <= io_A_Valid_3_delay_13_2;
    io_A_Valid_3_delay_15 <= io_A_Valid_3_delay_14_1;
    io_B_Valid_15_delay_1_2 <= io_B_Valid_15;
    io_B_Valid_15_delay_2_1 <= io_B_Valid_15_delay_1_2;
    io_B_Valid_15_delay_3 <= io_B_Valid_15_delay_2_1;
    io_A_Valid_3_delay_1_15 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_14 <= io_A_Valid_3_delay_1_15;
    io_A_Valid_3_delay_3_13 <= io_A_Valid_3_delay_2_14;
    io_A_Valid_3_delay_4_12 <= io_A_Valid_3_delay_3_13;
    io_A_Valid_3_delay_5_11 <= io_A_Valid_3_delay_4_12;
    io_A_Valid_3_delay_6_10 <= io_A_Valid_3_delay_5_11;
    io_A_Valid_3_delay_7_9 <= io_A_Valid_3_delay_6_10;
    io_A_Valid_3_delay_8_8 <= io_A_Valid_3_delay_7_9;
    io_A_Valid_3_delay_9_7 <= io_A_Valid_3_delay_8_8;
    io_A_Valid_3_delay_10_6 <= io_A_Valid_3_delay_9_7;
    io_A_Valid_3_delay_11_5 <= io_A_Valid_3_delay_10_6;
    io_A_Valid_3_delay_12_4 <= io_A_Valid_3_delay_11_5;
    io_A_Valid_3_delay_13_3 <= io_A_Valid_3_delay_12_4;
    io_A_Valid_3_delay_14_2 <= io_A_Valid_3_delay_13_3;
    io_A_Valid_3_delay_15_1 <= io_A_Valid_3_delay_14_2;
    io_A_Valid_3_delay_16 <= io_A_Valid_3_delay_15_1;
    io_B_Valid_16_delay_1_2 <= io_B_Valid_16;
    io_B_Valid_16_delay_2_1 <= io_B_Valid_16_delay_1_2;
    io_B_Valid_16_delay_3 <= io_B_Valid_16_delay_2_1;
    io_A_Valid_3_delay_1_16 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_15 <= io_A_Valid_3_delay_1_16;
    io_A_Valid_3_delay_3_14 <= io_A_Valid_3_delay_2_15;
    io_A_Valid_3_delay_4_13 <= io_A_Valid_3_delay_3_14;
    io_A_Valid_3_delay_5_12 <= io_A_Valid_3_delay_4_13;
    io_A_Valid_3_delay_6_11 <= io_A_Valid_3_delay_5_12;
    io_A_Valid_3_delay_7_10 <= io_A_Valid_3_delay_6_11;
    io_A_Valid_3_delay_8_9 <= io_A_Valid_3_delay_7_10;
    io_A_Valid_3_delay_9_8 <= io_A_Valid_3_delay_8_9;
    io_A_Valid_3_delay_10_7 <= io_A_Valid_3_delay_9_8;
    io_A_Valid_3_delay_11_6 <= io_A_Valid_3_delay_10_7;
    io_A_Valid_3_delay_12_5 <= io_A_Valid_3_delay_11_6;
    io_A_Valid_3_delay_13_4 <= io_A_Valid_3_delay_12_5;
    io_A_Valid_3_delay_14_3 <= io_A_Valid_3_delay_13_4;
    io_A_Valid_3_delay_15_2 <= io_A_Valid_3_delay_14_3;
    io_A_Valid_3_delay_16_1 <= io_A_Valid_3_delay_15_2;
    io_A_Valid_3_delay_17 <= io_A_Valid_3_delay_16_1;
    io_B_Valid_17_delay_1_2 <= io_B_Valid_17;
    io_B_Valid_17_delay_2_1 <= io_B_Valid_17_delay_1_2;
    io_B_Valid_17_delay_3 <= io_B_Valid_17_delay_2_1;
    io_A_Valid_3_delay_1_17 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_16 <= io_A_Valid_3_delay_1_17;
    io_A_Valid_3_delay_3_15 <= io_A_Valid_3_delay_2_16;
    io_A_Valid_3_delay_4_14 <= io_A_Valid_3_delay_3_15;
    io_A_Valid_3_delay_5_13 <= io_A_Valid_3_delay_4_14;
    io_A_Valid_3_delay_6_12 <= io_A_Valid_3_delay_5_13;
    io_A_Valid_3_delay_7_11 <= io_A_Valid_3_delay_6_12;
    io_A_Valid_3_delay_8_10 <= io_A_Valid_3_delay_7_11;
    io_A_Valid_3_delay_9_9 <= io_A_Valid_3_delay_8_10;
    io_A_Valid_3_delay_10_8 <= io_A_Valid_3_delay_9_9;
    io_A_Valid_3_delay_11_7 <= io_A_Valid_3_delay_10_8;
    io_A_Valid_3_delay_12_6 <= io_A_Valid_3_delay_11_7;
    io_A_Valid_3_delay_13_5 <= io_A_Valid_3_delay_12_6;
    io_A_Valid_3_delay_14_4 <= io_A_Valid_3_delay_13_5;
    io_A_Valid_3_delay_15_3 <= io_A_Valid_3_delay_14_4;
    io_A_Valid_3_delay_16_2 <= io_A_Valid_3_delay_15_3;
    io_A_Valid_3_delay_17_1 <= io_A_Valid_3_delay_16_2;
    io_A_Valid_3_delay_18 <= io_A_Valid_3_delay_17_1;
    io_B_Valid_18_delay_1_2 <= io_B_Valid_18;
    io_B_Valid_18_delay_2_1 <= io_B_Valid_18_delay_1_2;
    io_B_Valid_18_delay_3 <= io_B_Valid_18_delay_2_1;
    io_A_Valid_3_delay_1_18 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_17 <= io_A_Valid_3_delay_1_18;
    io_A_Valid_3_delay_3_16 <= io_A_Valid_3_delay_2_17;
    io_A_Valid_3_delay_4_15 <= io_A_Valid_3_delay_3_16;
    io_A_Valid_3_delay_5_14 <= io_A_Valid_3_delay_4_15;
    io_A_Valid_3_delay_6_13 <= io_A_Valid_3_delay_5_14;
    io_A_Valid_3_delay_7_12 <= io_A_Valid_3_delay_6_13;
    io_A_Valid_3_delay_8_11 <= io_A_Valid_3_delay_7_12;
    io_A_Valid_3_delay_9_10 <= io_A_Valid_3_delay_8_11;
    io_A_Valid_3_delay_10_9 <= io_A_Valid_3_delay_9_10;
    io_A_Valid_3_delay_11_8 <= io_A_Valid_3_delay_10_9;
    io_A_Valid_3_delay_12_7 <= io_A_Valid_3_delay_11_8;
    io_A_Valid_3_delay_13_6 <= io_A_Valid_3_delay_12_7;
    io_A_Valid_3_delay_14_5 <= io_A_Valid_3_delay_13_6;
    io_A_Valid_3_delay_15_4 <= io_A_Valid_3_delay_14_5;
    io_A_Valid_3_delay_16_3 <= io_A_Valid_3_delay_15_4;
    io_A_Valid_3_delay_17_2 <= io_A_Valid_3_delay_16_3;
    io_A_Valid_3_delay_18_1 <= io_A_Valid_3_delay_17_2;
    io_A_Valid_3_delay_19 <= io_A_Valid_3_delay_18_1;
    io_B_Valid_19_delay_1_2 <= io_B_Valid_19;
    io_B_Valid_19_delay_2_1 <= io_B_Valid_19_delay_1_2;
    io_B_Valid_19_delay_3 <= io_B_Valid_19_delay_2_1;
    io_A_Valid_3_delay_1_19 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_18 <= io_A_Valid_3_delay_1_19;
    io_A_Valid_3_delay_3_17 <= io_A_Valid_3_delay_2_18;
    io_A_Valid_3_delay_4_16 <= io_A_Valid_3_delay_3_17;
    io_A_Valid_3_delay_5_15 <= io_A_Valid_3_delay_4_16;
    io_A_Valid_3_delay_6_14 <= io_A_Valid_3_delay_5_15;
    io_A_Valid_3_delay_7_13 <= io_A_Valid_3_delay_6_14;
    io_A_Valid_3_delay_8_12 <= io_A_Valid_3_delay_7_13;
    io_A_Valid_3_delay_9_11 <= io_A_Valid_3_delay_8_12;
    io_A_Valid_3_delay_10_10 <= io_A_Valid_3_delay_9_11;
    io_A_Valid_3_delay_11_9 <= io_A_Valid_3_delay_10_10;
    io_A_Valid_3_delay_12_8 <= io_A_Valid_3_delay_11_9;
    io_A_Valid_3_delay_13_7 <= io_A_Valid_3_delay_12_8;
    io_A_Valid_3_delay_14_6 <= io_A_Valid_3_delay_13_7;
    io_A_Valid_3_delay_15_5 <= io_A_Valid_3_delay_14_6;
    io_A_Valid_3_delay_16_4 <= io_A_Valid_3_delay_15_5;
    io_A_Valid_3_delay_17_3 <= io_A_Valid_3_delay_16_4;
    io_A_Valid_3_delay_18_2 <= io_A_Valid_3_delay_17_3;
    io_A_Valid_3_delay_19_1 <= io_A_Valid_3_delay_18_2;
    io_A_Valid_3_delay_20 <= io_A_Valid_3_delay_19_1;
    io_B_Valid_20_delay_1_2 <= io_B_Valid_20;
    io_B_Valid_20_delay_2_1 <= io_B_Valid_20_delay_1_2;
    io_B_Valid_20_delay_3 <= io_B_Valid_20_delay_2_1;
    io_A_Valid_3_delay_1_20 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_19 <= io_A_Valid_3_delay_1_20;
    io_A_Valid_3_delay_3_18 <= io_A_Valid_3_delay_2_19;
    io_A_Valid_3_delay_4_17 <= io_A_Valid_3_delay_3_18;
    io_A_Valid_3_delay_5_16 <= io_A_Valid_3_delay_4_17;
    io_A_Valid_3_delay_6_15 <= io_A_Valid_3_delay_5_16;
    io_A_Valid_3_delay_7_14 <= io_A_Valid_3_delay_6_15;
    io_A_Valid_3_delay_8_13 <= io_A_Valid_3_delay_7_14;
    io_A_Valid_3_delay_9_12 <= io_A_Valid_3_delay_8_13;
    io_A_Valid_3_delay_10_11 <= io_A_Valid_3_delay_9_12;
    io_A_Valid_3_delay_11_10 <= io_A_Valid_3_delay_10_11;
    io_A_Valid_3_delay_12_9 <= io_A_Valid_3_delay_11_10;
    io_A_Valid_3_delay_13_8 <= io_A_Valid_3_delay_12_9;
    io_A_Valid_3_delay_14_7 <= io_A_Valid_3_delay_13_8;
    io_A_Valid_3_delay_15_6 <= io_A_Valid_3_delay_14_7;
    io_A_Valid_3_delay_16_5 <= io_A_Valid_3_delay_15_6;
    io_A_Valid_3_delay_17_4 <= io_A_Valid_3_delay_16_5;
    io_A_Valid_3_delay_18_3 <= io_A_Valid_3_delay_17_4;
    io_A_Valid_3_delay_19_2 <= io_A_Valid_3_delay_18_3;
    io_A_Valid_3_delay_20_1 <= io_A_Valid_3_delay_19_2;
    io_A_Valid_3_delay_21 <= io_A_Valid_3_delay_20_1;
    io_B_Valid_21_delay_1_2 <= io_B_Valid_21;
    io_B_Valid_21_delay_2_1 <= io_B_Valid_21_delay_1_2;
    io_B_Valid_21_delay_3 <= io_B_Valid_21_delay_2_1;
    io_A_Valid_3_delay_1_21 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_20 <= io_A_Valid_3_delay_1_21;
    io_A_Valid_3_delay_3_19 <= io_A_Valid_3_delay_2_20;
    io_A_Valid_3_delay_4_18 <= io_A_Valid_3_delay_3_19;
    io_A_Valid_3_delay_5_17 <= io_A_Valid_3_delay_4_18;
    io_A_Valid_3_delay_6_16 <= io_A_Valid_3_delay_5_17;
    io_A_Valid_3_delay_7_15 <= io_A_Valid_3_delay_6_16;
    io_A_Valid_3_delay_8_14 <= io_A_Valid_3_delay_7_15;
    io_A_Valid_3_delay_9_13 <= io_A_Valid_3_delay_8_14;
    io_A_Valid_3_delay_10_12 <= io_A_Valid_3_delay_9_13;
    io_A_Valid_3_delay_11_11 <= io_A_Valid_3_delay_10_12;
    io_A_Valid_3_delay_12_10 <= io_A_Valid_3_delay_11_11;
    io_A_Valid_3_delay_13_9 <= io_A_Valid_3_delay_12_10;
    io_A_Valid_3_delay_14_8 <= io_A_Valid_3_delay_13_9;
    io_A_Valid_3_delay_15_7 <= io_A_Valid_3_delay_14_8;
    io_A_Valid_3_delay_16_6 <= io_A_Valid_3_delay_15_7;
    io_A_Valid_3_delay_17_5 <= io_A_Valid_3_delay_16_6;
    io_A_Valid_3_delay_18_4 <= io_A_Valid_3_delay_17_5;
    io_A_Valid_3_delay_19_3 <= io_A_Valid_3_delay_18_4;
    io_A_Valid_3_delay_20_2 <= io_A_Valid_3_delay_19_3;
    io_A_Valid_3_delay_21_1 <= io_A_Valid_3_delay_20_2;
    io_A_Valid_3_delay_22 <= io_A_Valid_3_delay_21_1;
    io_B_Valid_22_delay_1_2 <= io_B_Valid_22;
    io_B_Valid_22_delay_2_1 <= io_B_Valid_22_delay_1_2;
    io_B_Valid_22_delay_3 <= io_B_Valid_22_delay_2_1;
    io_A_Valid_3_delay_1_22 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_21 <= io_A_Valid_3_delay_1_22;
    io_A_Valid_3_delay_3_20 <= io_A_Valid_3_delay_2_21;
    io_A_Valid_3_delay_4_19 <= io_A_Valid_3_delay_3_20;
    io_A_Valid_3_delay_5_18 <= io_A_Valid_3_delay_4_19;
    io_A_Valid_3_delay_6_17 <= io_A_Valid_3_delay_5_18;
    io_A_Valid_3_delay_7_16 <= io_A_Valid_3_delay_6_17;
    io_A_Valid_3_delay_8_15 <= io_A_Valid_3_delay_7_16;
    io_A_Valid_3_delay_9_14 <= io_A_Valid_3_delay_8_15;
    io_A_Valid_3_delay_10_13 <= io_A_Valid_3_delay_9_14;
    io_A_Valid_3_delay_11_12 <= io_A_Valid_3_delay_10_13;
    io_A_Valid_3_delay_12_11 <= io_A_Valid_3_delay_11_12;
    io_A_Valid_3_delay_13_10 <= io_A_Valid_3_delay_12_11;
    io_A_Valid_3_delay_14_9 <= io_A_Valid_3_delay_13_10;
    io_A_Valid_3_delay_15_8 <= io_A_Valid_3_delay_14_9;
    io_A_Valid_3_delay_16_7 <= io_A_Valid_3_delay_15_8;
    io_A_Valid_3_delay_17_6 <= io_A_Valid_3_delay_16_7;
    io_A_Valid_3_delay_18_5 <= io_A_Valid_3_delay_17_6;
    io_A_Valid_3_delay_19_4 <= io_A_Valid_3_delay_18_5;
    io_A_Valid_3_delay_20_3 <= io_A_Valid_3_delay_19_4;
    io_A_Valid_3_delay_21_2 <= io_A_Valid_3_delay_20_3;
    io_A_Valid_3_delay_22_1 <= io_A_Valid_3_delay_21_2;
    io_A_Valid_3_delay_23 <= io_A_Valid_3_delay_22_1;
    io_B_Valid_23_delay_1_2 <= io_B_Valid_23;
    io_B_Valid_23_delay_2_1 <= io_B_Valid_23_delay_1_2;
    io_B_Valid_23_delay_3 <= io_B_Valid_23_delay_2_1;
    io_A_Valid_3_delay_1_23 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_22 <= io_A_Valid_3_delay_1_23;
    io_A_Valid_3_delay_3_21 <= io_A_Valid_3_delay_2_22;
    io_A_Valid_3_delay_4_20 <= io_A_Valid_3_delay_3_21;
    io_A_Valid_3_delay_5_19 <= io_A_Valid_3_delay_4_20;
    io_A_Valid_3_delay_6_18 <= io_A_Valid_3_delay_5_19;
    io_A_Valid_3_delay_7_17 <= io_A_Valid_3_delay_6_18;
    io_A_Valid_3_delay_8_16 <= io_A_Valid_3_delay_7_17;
    io_A_Valid_3_delay_9_15 <= io_A_Valid_3_delay_8_16;
    io_A_Valid_3_delay_10_14 <= io_A_Valid_3_delay_9_15;
    io_A_Valid_3_delay_11_13 <= io_A_Valid_3_delay_10_14;
    io_A_Valid_3_delay_12_12 <= io_A_Valid_3_delay_11_13;
    io_A_Valid_3_delay_13_11 <= io_A_Valid_3_delay_12_12;
    io_A_Valid_3_delay_14_10 <= io_A_Valid_3_delay_13_11;
    io_A_Valid_3_delay_15_9 <= io_A_Valid_3_delay_14_10;
    io_A_Valid_3_delay_16_8 <= io_A_Valid_3_delay_15_9;
    io_A_Valid_3_delay_17_7 <= io_A_Valid_3_delay_16_8;
    io_A_Valid_3_delay_18_6 <= io_A_Valid_3_delay_17_7;
    io_A_Valid_3_delay_19_5 <= io_A_Valid_3_delay_18_6;
    io_A_Valid_3_delay_20_4 <= io_A_Valid_3_delay_19_5;
    io_A_Valid_3_delay_21_3 <= io_A_Valid_3_delay_20_4;
    io_A_Valid_3_delay_22_2 <= io_A_Valid_3_delay_21_3;
    io_A_Valid_3_delay_23_1 <= io_A_Valid_3_delay_22_2;
    io_A_Valid_3_delay_24 <= io_A_Valid_3_delay_23_1;
    io_B_Valid_24_delay_1_2 <= io_B_Valid_24;
    io_B_Valid_24_delay_2_1 <= io_B_Valid_24_delay_1_2;
    io_B_Valid_24_delay_3 <= io_B_Valid_24_delay_2_1;
    io_A_Valid_3_delay_1_24 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_23 <= io_A_Valid_3_delay_1_24;
    io_A_Valid_3_delay_3_22 <= io_A_Valid_3_delay_2_23;
    io_A_Valid_3_delay_4_21 <= io_A_Valid_3_delay_3_22;
    io_A_Valid_3_delay_5_20 <= io_A_Valid_3_delay_4_21;
    io_A_Valid_3_delay_6_19 <= io_A_Valid_3_delay_5_20;
    io_A_Valid_3_delay_7_18 <= io_A_Valid_3_delay_6_19;
    io_A_Valid_3_delay_8_17 <= io_A_Valid_3_delay_7_18;
    io_A_Valid_3_delay_9_16 <= io_A_Valid_3_delay_8_17;
    io_A_Valid_3_delay_10_15 <= io_A_Valid_3_delay_9_16;
    io_A_Valid_3_delay_11_14 <= io_A_Valid_3_delay_10_15;
    io_A_Valid_3_delay_12_13 <= io_A_Valid_3_delay_11_14;
    io_A_Valid_3_delay_13_12 <= io_A_Valid_3_delay_12_13;
    io_A_Valid_3_delay_14_11 <= io_A_Valid_3_delay_13_12;
    io_A_Valid_3_delay_15_10 <= io_A_Valid_3_delay_14_11;
    io_A_Valid_3_delay_16_9 <= io_A_Valid_3_delay_15_10;
    io_A_Valid_3_delay_17_8 <= io_A_Valid_3_delay_16_9;
    io_A_Valid_3_delay_18_7 <= io_A_Valid_3_delay_17_8;
    io_A_Valid_3_delay_19_6 <= io_A_Valid_3_delay_18_7;
    io_A_Valid_3_delay_20_5 <= io_A_Valid_3_delay_19_6;
    io_A_Valid_3_delay_21_4 <= io_A_Valid_3_delay_20_5;
    io_A_Valid_3_delay_22_3 <= io_A_Valid_3_delay_21_4;
    io_A_Valid_3_delay_23_2 <= io_A_Valid_3_delay_22_3;
    io_A_Valid_3_delay_24_1 <= io_A_Valid_3_delay_23_2;
    io_A_Valid_3_delay_25 <= io_A_Valid_3_delay_24_1;
    io_B_Valid_25_delay_1_2 <= io_B_Valid_25;
    io_B_Valid_25_delay_2_1 <= io_B_Valid_25_delay_1_2;
    io_B_Valid_25_delay_3 <= io_B_Valid_25_delay_2_1;
    io_A_Valid_3_delay_1_25 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_24 <= io_A_Valid_3_delay_1_25;
    io_A_Valid_3_delay_3_23 <= io_A_Valid_3_delay_2_24;
    io_A_Valid_3_delay_4_22 <= io_A_Valid_3_delay_3_23;
    io_A_Valid_3_delay_5_21 <= io_A_Valid_3_delay_4_22;
    io_A_Valid_3_delay_6_20 <= io_A_Valid_3_delay_5_21;
    io_A_Valid_3_delay_7_19 <= io_A_Valid_3_delay_6_20;
    io_A_Valid_3_delay_8_18 <= io_A_Valid_3_delay_7_19;
    io_A_Valid_3_delay_9_17 <= io_A_Valid_3_delay_8_18;
    io_A_Valid_3_delay_10_16 <= io_A_Valid_3_delay_9_17;
    io_A_Valid_3_delay_11_15 <= io_A_Valid_3_delay_10_16;
    io_A_Valid_3_delay_12_14 <= io_A_Valid_3_delay_11_15;
    io_A_Valid_3_delay_13_13 <= io_A_Valid_3_delay_12_14;
    io_A_Valid_3_delay_14_12 <= io_A_Valid_3_delay_13_13;
    io_A_Valid_3_delay_15_11 <= io_A_Valid_3_delay_14_12;
    io_A_Valid_3_delay_16_10 <= io_A_Valid_3_delay_15_11;
    io_A_Valid_3_delay_17_9 <= io_A_Valid_3_delay_16_10;
    io_A_Valid_3_delay_18_8 <= io_A_Valid_3_delay_17_9;
    io_A_Valid_3_delay_19_7 <= io_A_Valid_3_delay_18_8;
    io_A_Valid_3_delay_20_6 <= io_A_Valid_3_delay_19_7;
    io_A_Valid_3_delay_21_5 <= io_A_Valid_3_delay_20_6;
    io_A_Valid_3_delay_22_4 <= io_A_Valid_3_delay_21_5;
    io_A_Valid_3_delay_23_3 <= io_A_Valid_3_delay_22_4;
    io_A_Valid_3_delay_24_2 <= io_A_Valid_3_delay_23_3;
    io_A_Valid_3_delay_25_1 <= io_A_Valid_3_delay_24_2;
    io_A_Valid_3_delay_26 <= io_A_Valid_3_delay_25_1;
    io_B_Valid_26_delay_1_2 <= io_B_Valid_26;
    io_B_Valid_26_delay_2_1 <= io_B_Valid_26_delay_1_2;
    io_B_Valid_26_delay_3 <= io_B_Valid_26_delay_2_1;
    io_A_Valid_3_delay_1_26 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_25 <= io_A_Valid_3_delay_1_26;
    io_A_Valid_3_delay_3_24 <= io_A_Valid_3_delay_2_25;
    io_A_Valid_3_delay_4_23 <= io_A_Valid_3_delay_3_24;
    io_A_Valid_3_delay_5_22 <= io_A_Valid_3_delay_4_23;
    io_A_Valid_3_delay_6_21 <= io_A_Valid_3_delay_5_22;
    io_A_Valid_3_delay_7_20 <= io_A_Valid_3_delay_6_21;
    io_A_Valid_3_delay_8_19 <= io_A_Valid_3_delay_7_20;
    io_A_Valid_3_delay_9_18 <= io_A_Valid_3_delay_8_19;
    io_A_Valid_3_delay_10_17 <= io_A_Valid_3_delay_9_18;
    io_A_Valid_3_delay_11_16 <= io_A_Valid_3_delay_10_17;
    io_A_Valid_3_delay_12_15 <= io_A_Valid_3_delay_11_16;
    io_A_Valid_3_delay_13_14 <= io_A_Valid_3_delay_12_15;
    io_A_Valid_3_delay_14_13 <= io_A_Valid_3_delay_13_14;
    io_A_Valid_3_delay_15_12 <= io_A_Valid_3_delay_14_13;
    io_A_Valid_3_delay_16_11 <= io_A_Valid_3_delay_15_12;
    io_A_Valid_3_delay_17_10 <= io_A_Valid_3_delay_16_11;
    io_A_Valid_3_delay_18_9 <= io_A_Valid_3_delay_17_10;
    io_A_Valid_3_delay_19_8 <= io_A_Valid_3_delay_18_9;
    io_A_Valid_3_delay_20_7 <= io_A_Valid_3_delay_19_8;
    io_A_Valid_3_delay_21_6 <= io_A_Valid_3_delay_20_7;
    io_A_Valid_3_delay_22_5 <= io_A_Valid_3_delay_21_6;
    io_A_Valid_3_delay_23_4 <= io_A_Valid_3_delay_22_5;
    io_A_Valid_3_delay_24_3 <= io_A_Valid_3_delay_23_4;
    io_A_Valid_3_delay_25_2 <= io_A_Valid_3_delay_24_3;
    io_A_Valid_3_delay_26_1 <= io_A_Valid_3_delay_25_2;
    io_A_Valid_3_delay_27 <= io_A_Valid_3_delay_26_1;
    io_B_Valid_27_delay_1_2 <= io_B_Valid_27;
    io_B_Valid_27_delay_2_1 <= io_B_Valid_27_delay_1_2;
    io_B_Valid_27_delay_3 <= io_B_Valid_27_delay_2_1;
    io_A_Valid_3_delay_1_27 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_26 <= io_A_Valid_3_delay_1_27;
    io_A_Valid_3_delay_3_25 <= io_A_Valid_3_delay_2_26;
    io_A_Valid_3_delay_4_24 <= io_A_Valid_3_delay_3_25;
    io_A_Valid_3_delay_5_23 <= io_A_Valid_3_delay_4_24;
    io_A_Valid_3_delay_6_22 <= io_A_Valid_3_delay_5_23;
    io_A_Valid_3_delay_7_21 <= io_A_Valid_3_delay_6_22;
    io_A_Valid_3_delay_8_20 <= io_A_Valid_3_delay_7_21;
    io_A_Valid_3_delay_9_19 <= io_A_Valid_3_delay_8_20;
    io_A_Valid_3_delay_10_18 <= io_A_Valid_3_delay_9_19;
    io_A_Valid_3_delay_11_17 <= io_A_Valid_3_delay_10_18;
    io_A_Valid_3_delay_12_16 <= io_A_Valid_3_delay_11_17;
    io_A_Valid_3_delay_13_15 <= io_A_Valid_3_delay_12_16;
    io_A_Valid_3_delay_14_14 <= io_A_Valid_3_delay_13_15;
    io_A_Valid_3_delay_15_13 <= io_A_Valid_3_delay_14_14;
    io_A_Valid_3_delay_16_12 <= io_A_Valid_3_delay_15_13;
    io_A_Valid_3_delay_17_11 <= io_A_Valid_3_delay_16_12;
    io_A_Valid_3_delay_18_10 <= io_A_Valid_3_delay_17_11;
    io_A_Valid_3_delay_19_9 <= io_A_Valid_3_delay_18_10;
    io_A_Valid_3_delay_20_8 <= io_A_Valid_3_delay_19_9;
    io_A_Valid_3_delay_21_7 <= io_A_Valid_3_delay_20_8;
    io_A_Valid_3_delay_22_6 <= io_A_Valid_3_delay_21_7;
    io_A_Valid_3_delay_23_5 <= io_A_Valid_3_delay_22_6;
    io_A_Valid_3_delay_24_4 <= io_A_Valid_3_delay_23_5;
    io_A_Valid_3_delay_25_3 <= io_A_Valid_3_delay_24_4;
    io_A_Valid_3_delay_26_2 <= io_A_Valid_3_delay_25_3;
    io_A_Valid_3_delay_27_1 <= io_A_Valid_3_delay_26_2;
    io_A_Valid_3_delay_28 <= io_A_Valid_3_delay_27_1;
    io_B_Valid_28_delay_1_2 <= io_B_Valid_28;
    io_B_Valid_28_delay_2_1 <= io_B_Valid_28_delay_1_2;
    io_B_Valid_28_delay_3 <= io_B_Valid_28_delay_2_1;
    io_A_Valid_3_delay_1_28 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_27 <= io_A_Valid_3_delay_1_28;
    io_A_Valid_3_delay_3_26 <= io_A_Valid_3_delay_2_27;
    io_A_Valid_3_delay_4_25 <= io_A_Valid_3_delay_3_26;
    io_A_Valid_3_delay_5_24 <= io_A_Valid_3_delay_4_25;
    io_A_Valid_3_delay_6_23 <= io_A_Valid_3_delay_5_24;
    io_A_Valid_3_delay_7_22 <= io_A_Valid_3_delay_6_23;
    io_A_Valid_3_delay_8_21 <= io_A_Valid_3_delay_7_22;
    io_A_Valid_3_delay_9_20 <= io_A_Valid_3_delay_8_21;
    io_A_Valid_3_delay_10_19 <= io_A_Valid_3_delay_9_20;
    io_A_Valid_3_delay_11_18 <= io_A_Valid_3_delay_10_19;
    io_A_Valid_3_delay_12_17 <= io_A_Valid_3_delay_11_18;
    io_A_Valid_3_delay_13_16 <= io_A_Valid_3_delay_12_17;
    io_A_Valid_3_delay_14_15 <= io_A_Valid_3_delay_13_16;
    io_A_Valid_3_delay_15_14 <= io_A_Valid_3_delay_14_15;
    io_A_Valid_3_delay_16_13 <= io_A_Valid_3_delay_15_14;
    io_A_Valid_3_delay_17_12 <= io_A_Valid_3_delay_16_13;
    io_A_Valid_3_delay_18_11 <= io_A_Valid_3_delay_17_12;
    io_A_Valid_3_delay_19_10 <= io_A_Valid_3_delay_18_11;
    io_A_Valid_3_delay_20_9 <= io_A_Valid_3_delay_19_10;
    io_A_Valid_3_delay_21_8 <= io_A_Valid_3_delay_20_9;
    io_A_Valid_3_delay_22_7 <= io_A_Valid_3_delay_21_8;
    io_A_Valid_3_delay_23_6 <= io_A_Valid_3_delay_22_7;
    io_A_Valid_3_delay_24_5 <= io_A_Valid_3_delay_23_6;
    io_A_Valid_3_delay_25_4 <= io_A_Valid_3_delay_24_5;
    io_A_Valid_3_delay_26_3 <= io_A_Valid_3_delay_25_4;
    io_A_Valid_3_delay_27_2 <= io_A_Valid_3_delay_26_3;
    io_A_Valid_3_delay_28_1 <= io_A_Valid_3_delay_27_2;
    io_A_Valid_3_delay_29 <= io_A_Valid_3_delay_28_1;
    io_B_Valid_29_delay_1_2 <= io_B_Valid_29;
    io_B_Valid_29_delay_2_1 <= io_B_Valid_29_delay_1_2;
    io_B_Valid_29_delay_3 <= io_B_Valid_29_delay_2_1;
    io_A_Valid_3_delay_1_29 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_28 <= io_A_Valid_3_delay_1_29;
    io_A_Valid_3_delay_3_27 <= io_A_Valid_3_delay_2_28;
    io_A_Valid_3_delay_4_26 <= io_A_Valid_3_delay_3_27;
    io_A_Valid_3_delay_5_25 <= io_A_Valid_3_delay_4_26;
    io_A_Valid_3_delay_6_24 <= io_A_Valid_3_delay_5_25;
    io_A_Valid_3_delay_7_23 <= io_A_Valid_3_delay_6_24;
    io_A_Valid_3_delay_8_22 <= io_A_Valid_3_delay_7_23;
    io_A_Valid_3_delay_9_21 <= io_A_Valid_3_delay_8_22;
    io_A_Valid_3_delay_10_20 <= io_A_Valid_3_delay_9_21;
    io_A_Valid_3_delay_11_19 <= io_A_Valid_3_delay_10_20;
    io_A_Valid_3_delay_12_18 <= io_A_Valid_3_delay_11_19;
    io_A_Valid_3_delay_13_17 <= io_A_Valid_3_delay_12_18;
    io_A_Valid_3_delay_14_16 <= io_A_Valid_3_delay_13_17;
    io_A_Valid_3_delay_15_15 <= io_A_Valid_3_delay_14_16;
    io_A_Valid_3_delay_16_14 <= io_A_Valid_3_delay_15_15;
    io_A_Valid_3_delay_17_13 <= io_A_Valid_3_delay_16_14;
    io_A_Valid_3_delay_18_12 <= io_A_Valid_3_delay_17_13;
    io_A_Valid_3_delay_19_11 <= io_A_Valid_3_delay_18_12;
    io_A_Valid_3_delay_20_10 <= io_A_Valid_3_delay_19_11;
    io_A_Valid_3_delay_21_9 <= io_A_Valid_3_delay_20_10;
    io_A_Valid_3_delay_22_8 <= io_A_Valid_3_delay_21_9;
    io_A_Valid_3_delay_23_7 <= io_A_Valid_3_delay_22_8;
    io_A_Valid_3_delay_24_6 <= io_A_Valid_3_delay_23_7;
    io_A_Valid_3_delay_25_5 <= io_A_Valid_3_delay_24_6;
    io_A_Valid_3_delay_26_4 <= io_A_Valid_3_delay_25_5;
    io_A_Valid_3_delay_27_3 <= io_A_Valid_3_delay_26_4;
    io_A_Valid_3_delay_28_2 <= io_A_Valid_3_delay_27_3;
    io_A_Valid_3_delay_29_1 <= io_A_Valid_3_delay_28_2;
    io_A_Valid_3_delay_30 <= io_A_Valid_3_delay_29_1;
    io_B_Valid_30_delay_1_2 <= io_B_Valid_30;
    io_B_Valid_30_delay_2_1 <= io_B_Valid_30_delay_1_2;
    io_B_Valid_30_delay_3 <= io_B_Valid_30_delay_2_1;
    io_A_Valid_3_delay_1_30 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_29 <= io_A_Valid_3_delay_1_30;
    io_A_Valid_3_delay_3_28 <= io_A_Valid_3_delay_2_29;
    io_A_Valid_3_delay_4_27 <= io_A_Valid_3_delay_3_28;
    io_A_Valid_3_delay_5_26 <= io_A_Valid_3_delay_4_27;
    io_A_Valid_3_delay_6_25 <= io_A_Valid_3_delay_5_26;
    io_A_Valid_3_delay_7_24 <= io_A_Valid_3_delay_6_25;
    io_A_Valid_3_delay_8_23 <= io_A_Valid_3_delay_7_24;
    io_A_Valid_3_delay_9_22 <= io_A_Valid_3_delay_8_23;
    io_A_Valid_3_delay_10_21 <= io_A_Valid_3_delay_9_22;
    io_A_Valid_3_delay_11_20 <= io_A_Valid_3_delay_10_21;
    io_A_Valid_3_delay_12_19 <= io_A_Valid_3_delay_11_20;
    io_A_Valid_3_delay_13_18 <= io_A_Valid_3_delay_12_19;
    io_A_Valid_3_delay_14_17 <= io_A_Valid_3_delay_13_18;
    io_A_Valid_3_delay_15_16 <= io_A_Valid_3_delay_14_17;
    io_A_Valid_3_delay_16_15 <= io_A_Valid_3_delay_15_16;
    io_A_Valid_3_delay_17_14 <= io_A_Valid_3_delay_16_15;
    io_A_Valid_3_delay_18_13 <= io_A_Valid_3_delay_17_14;
    io_A_Valid_3_delay_19_12 <= io_A_Valid_3_delay_18_13;
    io_A_Valid_3_delay_20_11 <= io_A_Valid_3_delay_19_12;
    io_A_Valid_3_delay_21_10 <= io_A_Valid_3_delay_20_11;
    io_A_Valid_3_delay_22_9 <= io_A_Valid_3_delay_21_10;
    io_A_Valid_3_delay_23_8 <= io_A_Valid_3_delay_22_9;
    io_A_Valid_3_delay_24_7 <= io_A_Valid_3_delay_23_8;
    io_A_Valid_3_delay_25_6 <= io_A_Valid_3_delay_24_7;
    io_A_Valid_3_delay_26_5 <= io_A_Valid_3_delay_25_6;
    io_A_Valid_3_delay_27_4 <= io_A_Valid_3_delay_26_5;
    io_A_Valid_3_delay_28_3 <= io_A_Valid_3_delay_27_4;
    io_A_Valid_3_delay_29_2 <= io_A_Valid_3_delay_28_3;
    io_A_Valid_3_delay_30_1 <= io_A_Valid_3_delay_29_2;
    io_A_Valid_3_delay_31 <= io_A_Valid_3_delay_30_1;
    io_B_Valid_31_delay_1_2 <= io_B_Valid_31;
    io_B_Valid_31_delay_2_1 <= io_B_Valid_31_delay_1_2;
    io_B_Valid_31_delay_3 <= io_B_Valid_31_delay_2_1;
    io_A_Valid_3_delay_1_31 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_30 <= io_A_Valid_3_delay_1_31;
    io_A_Valid_3_delay_3_29 <= io_A_Valid_3_delay_2_30;
    io_A_Valid_3_delay_4_28 <= io_A_Valid_3_delay_3_29;
    io_A_Valid_3_delay_5_27 <= io_A_Valid_3_delay_4_28;
    io_A_Valid_3_delay_6_26 <= io_A_Valid_3_delay_5_27;
    io_A_Valid_3_delay_7_25 <= io_A_Valid_3_delay_6_26;
    io_A_Valid_3_delay_8_24 <= io_A_Valid_3_delay_7_25;
    io_A_Valid_3_delay_9_23 <= io_A_Valid_3_delay_8_24;
    io_A_Valid_3_delay_10_22 <= io_A_Valid_3_delay_9_23;
    io_A_Valid_3_delay_11_21 <= io_A_Valid_3_delay_10_22;
    io_A_Valid_3_delay_12_20 <= io_A_Valid_3_delay_11_21;
    io_A_Valid_3_delay_13_19 <= io_A_Valid_3_delay_12_20;
    io_A_Valid_3_delay_14_18 <= io_A_Valid_3_delay_13_19;
    io_A_Valid_3_delay_15_17 <= io_A_Valid_3_delay_14_18;
    io_A_Valid_3_delay_16_16 <= io_A_Valid_3_delay_15_17;
    io_A_Valid_3_delay_17_15 <= io_A_Valid_3_delay_16_16;
    io_A_Valid_3_delay_18_14 <= io_A_Valid_3_delay_17_15;
    io_A_Valid_3_delay_19_13 <= io_A_Valid_3_delay_18_14;
    io_A_Valid_3_delay_20_12 <= io_A_Valid_3_delay_19_13;
    io_A_Valid_3_delay_21_11 <= io_A_Valid_3_delay_20_12;
    io_A_Valid_3_delay_22_10 <= io_A_Valid_3_delay_21_11;
    io_A_Valid_3_delay_23_9 <= io_A_Valid_3_delay_22_10;
    io_A_Valid_3_delay_24_8 <= io_A_Valid_3_delay_23_9;
    io_A_Valid_3_delay_25_7 <= io_A_Valid_3_delay_24_8;
    io_A_Valid_3_delay_26_6 <= io_A_Valid_3_delay_25_7;
    io_A_Valid_3_delay_27_5 <= io_A_Valid_3_delay_26_6;
    io_A_Valid_3_delay_28_4 <= io_A_Valid_3_delay_27_5;
    io_A_Valid_3_delay_29_3 <= io_A_Valid_3_delay_28_4;
    io_A_Valid_3_delay_30_2 <= io_A_Valid_3_delay_29_3;
    io_A_Valid_3_delay_31_1 <= io_A_Valid_3_delay_30_2;
    io_A_Valid_3_delay_32 <= io_A_Valid_3_delay_31_1;
    io_B_Valid_32_delay_1_2 <= io_B_Valid_32;
    io_B_Valid_32_delay_2_1 <= io_B_Valid_32_delay_1_2;
    io_B_Valid_32_delay_3 <= io_B_Valid_32_delay_2_1;
    io_A_Valid_3_delay_1_32 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_31 <= io_A_Valid_3_delay_1_32;
    io_A_Valid_3_delay_3_30 <= io_A_Valid_3_delay_2_31;
    io_A_Valid_3_delay_4_29 <= io_A_Valid_3_delay_3_30;
    io_A_Valid_3_delay_5_28 <= io_A_Valid_3_delay_4_29;
    io_A_Valid_3_delay_6_27 <= io_A_Valid_3_delay_5_28;
    io_A_Valid_3_delay_7_26 <= io_A_Valid_3_delay_6_27;
    io_A_Valid_3_delay_8_25 <= io_A_Valid_3_delay_7_26;
    io_A_Valid_3_delay_9_24 <= io_A_Valid_3_delay_8_25;
    io_A_Valid_3_delay_10_23 <= io_A_Valid_3_delay_9_24;
    io_A_Valid_3_delay_11_22 <= io_A_Valid_3_delay_10_23;
    io_A_Valid_3_delay_12_21 <= io_A_Valid_3_delay_11_22;
    io_A_Valid_3_delay_13_20 <= io_A_Valid_3_delay_12_21;
    io_A_Valid_3_delay_14_19 <= io_A_Valid_3_delay_13_20;
    io_A_Valid_3_delay_15_18 <= io_A_Valid_3_delay_14_19;
    io_A_Valid_3_delay_16_17 <= io_A_Valid_3_delay_15_18;
    io_A_Valid_3_delay_17_16 <= io_A_Valid_3_delay_16_17;
    io_A_Valid_3_delay_18_15 <= io_A_Valid_3_delay_17_16;
    io_A_Valid_3_delay_19_14 <= io_A_Valid_3_delay_18_15;
    io_A_Valid_3_delay_20_13 <= io_A_Valid_3_delay_19_14;
    io_A_Valid_3_delay_21_12 <= io_A_Valid_3_delay_20_13;
    io_A_Valid_3_delay_22_11 <= io_A_Valid_3_delay_21_12;
    io_A_Valid_3_delay_23_10 <= io_A_Valid_3_delay_22_11;
    io_A_Valid_3_delay_24_9 <= io_A_Valid_3_delay_23_10;
    io_A_Valid_3_delay_25_8 <= io_A_Valid_3_delay_24_9;
    io_A_Valid_3_delay_26_7 <= io_A_Valid_3_delay_25_8;
    io_A_Valid_3_delay_27_6 <= io_A_Valid_3_delay_26_7;
    io_A_Valid_3_delay_28_5 <= io_A_Valid_3_delay_27_6;
    io_A_Valid_3_delay_29_4 <= io_A_Valid_3_delay_28_5;
    io_A_Valid_3_delay_30_3 <= io_A_Valid_3_delay_29_4;
    io_A_Valid_3_delay_31_2 <= io_A_Valid_3_delay_30_3;
    io_A_Valid_3_delay_32_1 <= io_A_Valid_3_delay_31_2;
    io_A_Valid_3_delay_33 <= io_A_Valid_3_delay_32_1;
    io_B_Valid_33_delay_1_2 <= io_B_Valid_33;
    io_B_Valid_33_delay_2_1 <= io_B_Valid_33_delay_1_2;
    io_B_Valid_33_delay_3 <= io_B_Valid_33_delay_2_1;
    io_A_Valid_3_delay_1_33 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_32 <= io_A_Valid_3_delay_1_33;
    io_A_Valid_3_delay_3_31 <= io_A_Valid_3_delay_2_32;
    io_A_Valid_3_delay_4_30 <= io_A_Valid_3_delay_3_31;
    io_A_Valid_3_delay_5_29 <= io_A_Valid_3_delay_4_30;
    io_A_Valid_3_delay_6_28 <= io_A_Valid_3_delay_5_29;
    io_A_Valid_3_delay_7_27 <= io_A_Valid_3_delay_6_28;
    io_A_Valid_3_delay_8_26 <= io_A_Valid_3_delay_7_27;
    io_A_Valid_3_delay_9_25 <= io_A_Valid_3_delay_8_26;
    io_A_Valid_3_delay_10_24 <= io_A_Valid_3_delay_9_25;
    io_A_Valid_3_delay_11_23 <= io_A_Valid_3_delay_10_24;
    io_A_Valid_3_delay_12_22 <= io_A_Valid_3_delay_11_23;
    io_A_Valid_3_delay_13_21 <= io_A_Valid_3_delay_12_22;
    io_A_Valid_3_delay_14_20 <= io_A_Valid_3_delay_13_21;
    io_A_Valid_3_delay_15_19 <= io_A_Valid_3_delay_14_20;
    io_A_Valid_3_delay_16_18 <= io_A_Valid_3_delay_15_19;
    io_A_Valid_3_delay_17_17 <= io_A_Valid_3_delay_16_18;
    io_A_Valid_3_delay_18_16 <= io_A_Valid_3_delay_17_17;
    io_A_Valid_3_delay_19_15 <= io_A_Valid_3_delay_18_16;
    io_A_Valid_3_delay_20_14 <= io_A_Valid_3_delay_19_15;
    io_A_Valid_3_delay_21_13 <= io_A_Valid_3_delay_20_14;
    io_A_Valid_3_delay_22_12 <= io_A_Valid_3_delay_21_13;
    io_A_Valid_3_delay_23_11 <= io_A_Valid_3_delay_22_12;
    io_A_Valid_3_delay_24_10 <= io_A_Valid_3_delay_23_11;
    io_A_Valid_3_delay_25_9 <= io_A_Valid_3_delay_24_10;
    io_A_Valid_3_delay_26_8 <= io_A_Valid_3_delay_25_9;
    io_A_Valid_3_delay_27_7 <= io_A_Valid_3_delay_26_8;
    io_A_Valid_3_delay_28_6 <= io_A_Valid_3_delay_27_7;
    io_A_Valid_3_delay_29_5 <= io_A_Valid_3_delay_28_6;
    io_A_Valid_3_delay_30_4 <= io_A_Valid_3_delay_29_5;
    io_A_Valid_3_delay_31_3 <= io_A_Valid_3_delay_30_4;
    io_A_Valid_3_delay_32_2 <= io_A_Valid_3_delay_31_3;
    io_A_Valid_3_delay_33_1 <= io_A_Valid_3_delay_32_2;
    io_A_Valid_3_delay_34 <= io_A_Valid_3_delay_33_1;
    io_B_Valid_34_delay_1_2 <= io_B_Valid_34;
    io_B_Valid_34_delay_2_1 <= io_B_Valid_34_delay_1_2;
    io_B_Valid_34_delay_3 <= io_B_Valid_34_delay_2_1;
    io_A_Valid_3_delay_1_34 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_33 <= io_A_Valid_3_delay_1_34;
    io_A_Valid_3_delay_3_32 <= io_A_Valid_3_delay_2_33;
    io_A_Valid_3_delay_4_31 <= io_A_Valid_3_delay_3_32;
    io_A_Valid_3_delay_5_30 <= io_A_Valid_3_delay_4_31;
    io_A_Valid_3_delay_6_29 <= io_A_Valid_3_delay_5_30;
    io_A_Valid_3_delay_7_28 <= io_A_Valid_3_delay_6_29;
    io_A_Valid_3_delay_8_27 <= io_A_Valid_3_delay_7_28;
    io_A_Valid_3_delay_9_26 <= io_A_Valid_3_delay_8_27;
    io_A_Valid_3_delay_10_25 <= io_A_Valid_3_delay_9_26;
    io_A_Valid_3_delay_11_24 <= io_A_Valid_3_delay_10_25;
    io_A_Valid_3_delay_12_23 <= io_A_Valid_3_delay_11_24;
    io_A_Valid_3_delay_13_22 <= io_A_Valid_3_delay_12_23;
    io_A_Valid_3_delay_14_21 <= io_A_Valid_3_delay_13_22;
    io_A_Valid_3_delay_15_20 <= io_A_Valid_3_delay_14_21;
    io_A_Valid_3_delay_16_19 <= io_A_Valid_3_delay_15_20;
    io_A_Valid_3_delay_17_18 <= io_A_Valid_3_delay_16_19;
    io_A_Valid_3_delay_18_17 <= io_A_Valid_3_delay_17_18;
    io_A_Valid_3_delay_19_16 <= io_A_Valid_3_delay_18_17;
    io_A_Valid_3_delay_20_15 <= io_A_Valid_3_delay_19_16;
    io_A_Valid_3_delay_21_14 <= io_A_Valid_3_delay_20_15;
    io_A_Valid_3_delay_22_13 <= io_A_Valid_3_delay_21_14;
    io_A_Valid_3_delay_23_12 <= io_A_Valid_3_delay_22_13;
    io_A_Valid_3_delay_24_11 <= io_A_Valid_3_delay_23_12;
    io_A_Valid_3_delay_25_10 <= io_A_Valid_3_delay_24_11;
    io_A_Valid_3_delay_26_9 <= io_A_Valid_3_delay_25_10;
    io_A_Valid_3_delay_27_8 <= io_A_Valid_3_delay_26_9;
    io_A_Valid_3_delay_28_7 <= io_A_Valid_3_delay_27_8;
    io_A_Valid_3_delay_29_6 <= io_A_Valid_3_delay_28_7;
    io_A_Valid_3_delay_30_5 <= io_A_Valid_3_delay_29_6;
    io_A_Valid_3_delay_31_4 <= io_A_Valid_3_delay_30_5;
    io_A_Valid_3_delay_32_3 <= io_A_Valid_3_delay_31_4;
    io_A_Valid_3_delay_33_2 <= io_A_Valid_3_delay_32_3;
    io_A_Valid_3_delay_34_1 <= io_A_Valid_3_delay_33_2;
    io_A_Valid_3_delay_35 <= io_A_Valid_3_delay_34_1;
    io_B_Valid_35_delay_1_2 <= io_B_Valid_35;
    io_B_Valid_35_delay_2_1 <= io_B_Valid_35_delay_1_2;
    io_B_Valid_35_delay_3 <= io_B_Valid_35_delay_2_1;
    io_A_Valid_3_delay_1_35 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_34 <= io_A_Valid_3_delay_1_35;
    io_A_Valid_3_delay_3_33 <= io_A_Valid_3_delay_2_34;
    io_A_Valid_3_delay_4_32 <= io_A_Valid_3_delay_3_33;
    io_A_Valid_3_delay_5_31 <= io_A_Valid_3_delay_4_32;
    io_A_Valid_3_delay_6_30 <= io_A_Valid_3_delay_5_31;
    io_A_Valid_3_delay_7_29 <= io_A_Valid_3_delay_6_30;
    io_A_Valid_3_delay_8_28 <= io_A_Valid_3_delay_7_29;
    io_A_Valid_3_delay_9_27 <= io_A_Valid_3_delay_8_28;
    io_A_Valid_3_delay_10_26 <= io_A_Valid_3_delay_9_27;
    io_A_Valid_3_delay_11_25 <= io_A_Valid_3_delay_10_26;
    io_A_Valid_3_delay_12_24 <= io_A_Valid_3_delay_11_25;
    io_A_Valid_3_delay_13_23 <= io_A_Valid_3_delay_12_24;
    io_A_Valid_3_delay_14_22 <= io_A_Valid_3_delay_13_23;
    io_A_Valid_3_delay_15_21 <= io_A_Valid_3_delay_14_22;
    io_A_Valid_3_delay_16_20 <= io_A_Valid_3_delay_15_21;
    io_A_Valid_3_delay_17_19 <= io_A_Valid_3_delay_16_20;
    io_A_Valid_3_delay_18_18 <= io_A_Valid_3_delay_17_19;
    io_A_Valid_3_delay_19_17 <= io_A_Valid_3_delay_18_18;
    io_A_Valid_3_delay_20_16 <= io_A_Valid_3_delay_19_17;
    io_A_Valid_3_delay_21_15 <= io_A_Valid_3_delay_20_16;
    io_A_Valid_3_delay_22_14 <= io_A_Valid_3_delay_21_15;
    io_A_Valid_3_delay_23_13 <= io_A_Valid_3_delay_22_14;
    io_A_Valid_3_delay_24_12 <= io_A_Valid_3_delay_23_13;
    io_A_Valid_3_delay_25_11 <= io_A_Valid_3_delay_24_12;
    io_A_Valid_3_delay_26_10 <= io_A_Valid_3_delay_25_11;
    io_A_Valid_3_delay_27_9 <= io_A_Valid_3_delay_26_10;
    io_A_Valid_3_delay_28_8 <= io_A_Valid_3_delay_27_9;
    io_A_Valid_3_delay_29_7 <= io_A_Valid_3_delay_28_8;
    io_A_Valid_3_delay_30_6 <= io_A_Valid_3_delay_29_7;
    io_A_Valid_3_delay_31_5 <= io_A_Valid_3_delay_30_6;
    io_A_Valid_3_delay_32_4 <= io_A_Valid_3_delay_31_5;
    io_A_Valid_3_delay_33_3 <= io_A_Valid_3_delay_32_4;
    io_A_Valid_3_delay_34_2 <= io_A_Valid_3_delay_33_3;
    io_A_Valid_3_delay_35_1 <= io_A_Valid_3_delay_34_2;
    io_A_Valid_3_delay_36 <= io_A_Valid_3_delay_35_1;
    io_B_Valid_36_delay_1_2 <= io_B_Valid_36;
    io_B_Valid_36_delay_2_1 <= io_B_Valid_36_delay_1_2;
    io_B_Valid_36_delay_3 <= io_B_Valid_36_delay_2_1;
    io_A_Valid_3_delay_1_36 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_35 <= io_A_Valid_3_delay_1_36;
    io_A_Valid_3_delay_3_34 <= io_A_Valid_3_delay_2_35;
    io_A_Valid_3_delay_4_33 <= io_A_Valid_3_delay_3_34;
    io_A_Valid_3_delay_5_32 <= io_A_Valid_3_delay_4_33;
    io_A_Valid_3_delay_6_31 <= io_A_Valid_3_delay_5_32;
    io_A_Valid_3_delay_7_30 <= io_A_Valid_3_delay_6_31;
    io_A_Valid_3_delay_8_29 <= io_A_Valid_3_delay_7_30;
    io_A_Valid_3_delay_9_28 <= io_A_Valid_3_delay_8_29;
    io_A_Valid_3_delay_10_27 <= io_A_Valid_3_delay_9_28;
    io_A_Valid_3_delay_11_26 <= io_A_Valid_3_delay_10_27;
    io_A_Valid_3_delay_12_25 <= io_A_Valid_3_delay_11_26;
    io_A_Valid_3_delay_13_24 <= io_A_Valid_3_delay_12_25;
    io_A_Valid_3_delay_14_23 <= io_A_Valid_3_delay_13_24;
    io_A_Valid_3_delay_15_22 <= io_A_Valid_3_delay_14_23;
    io_A_Valid_3_delay_16_21 <= io_A_Valid_3_delay_15_22;
    io_A_Valid_3_delay_17_20 <= io_A_Valid_3_delay_16_21;
    io_A_Valid_3_delay_18_19 <= io_A_Valid_3_delay_17_20;
    io_A_Valid_3_delay_19_18 <= io_A_Valid_3_delay_18_19;
    io_A_Valid_3_delay_20_17 <= io_A_Valid_3_delay_19_18;
    io_A_Valid_3_delay_21_16 <= io_A_Valid_3_delay_20_17;
    io_A_Valid_3_delay_22_15 <= io_A_Valid_3_delay_21_16;
    io_A_Valid_3_delay_23_14 <= io_A_Valid_3_delay_22_15;
    io_A_Valid_3_delay_24_13 <= io_A_Valid_3_delay_23_14;
    io_A_Valid_3_delay_25_12 <= io_A_Valid_3_delay_24_13;
    io_A_Valid_3_delay_26_11 <= io_A_Valid_3_delay_25_12;
    io_A_Valid_3_delay_27_10 <= io_A_Valid_3_delay_26_11;
    io_A_Valid_3_delay_28_9 <= io_A_Valid_3_delay_27_10;
    io_A_Valid_3_delay_29_8 <= io_A_Valid_3_delay_28_9;
    io_A_Valid_3_delay_30_7 <= io_A_Valid_3_delay_29_8;
    io_A_Valid_3_delay_31_6 <= io_A_Valid_3_delay_30_7;
    io_A_Valid_3_delay_32_5 <= io_A_Valid_3_delay_31_6;
    io_A_Valid_3_delay_33_4 <= io_A_Valid_3_delay_32_5;
    io_A_Valid_3_delay_34_3 <= io_A_Valid_3_delay_33_4;
    io_A_Valid_3_delay_35_2 <= io_A_Valid_3_delay_34_3;
    io_A_Valid_3_delay_36_1 <= io_A_Valid_3_delay_35_2;
    io_A_Valid_3_delay_37 <= io_A_Valid_3_delay_36_1;
    io_B_Valid_37_delay_1_2 <= io_B_Valid_37;
    io_B_Valid_37_delay_2_1 <= io_B_Valid_37_delay_1_2;
    io_B_Valid_37_delay_3 <= io_B_Valid_37_delay_2_1;
    io_A_Valid_3_delay_1_37 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_36 <= io_A_Valid_3_delay_1_37;
    io_A_Valid_3_delay_3_35 <= io_A_Valid_3_delay_2_36;
    io_A_Valid_3_delay_4_34 <= io_A_Valid_3_delay_3_35;
    io_A_Valid_3_delay_5_33 <= io_A_Valid_3_delay_4_34;
    io_A_Valid_3_delay_6_32 <= io_A_Valid_3_delay_5_33;
    io_A_Valid_3_delay_7_31 <= io_A_Valid_3_delay_6_32;
    io_A_Valid_3_delay_8_30 <= io_A_Valid_3_delay_7_31;
    io_A_Valid_3_delay_9_29 <= io_A_Valid_3_delay_8_30;
    io_A_Valid_3_delay_10_28 <= io_A_Valid_3_delay_9_29;
    io_A_Valid_3_delay_11_27 <= io_A_Valid_3_delay_10_28;
    io_A_Valid_3_delay_12_26 <= io_A_Valid_3_delay_11_27;
    io_A_Valid_3_delay_13_25 <= io_A_Valid_3_delay_12_26;
    io_A_Valid_3_delay_14_24 <= io_A_Valid_3_delay_13_25;
    io_A_Valid_3_delay_15_23 <= io_A_Valid_3_delay_14_24;
    io_A_Valid_3_delay_16_22 <= io_A_Valid_3_delay_15_23;
    io_A_Valid_3_delay_17_21 <= io_A_Valid_3_delay_16_22;
    io_A_Valid_3_delay_18_20 <= io_A_Valid_3_delay_17_21;
    io_A_Valid_3_delay_19_19 <= io_A_Valid_3_delay_18_20;
    io_A_Valid_3_delay_20_18 <= io_A_Valid_3_delay_19_19;
    io_A_Valid_3_delay_21_17 <= io_A_Valid_3_delay_20_18;
    io_A_Valid_3_delay_22_16 <= io_A_Valid_3_delay_21_17;
    io_A_Valid_3_delay_23_15 <= io_A_Valid_3_delay_22_16;
    io_A_Valid_3_delay_24_14 <= io_A_Valid_3_delay_23_15;
    io_A_Valid_3_delay_25_13 <= io_A_Valid_3_delay_24_14;
    io_A_Valid_3_delay_26_12 <= io_A_Valid_3_delay_25_13;
    io_A_Valid_3_delay_27_11 <= io_A_Valid_3_delay_26_12;
    io_A_Valid_3_delay_28_10 <= io_A_Valid_3_delay_27_11;
    io_A_Valid_3_delay_29_9 <= io_A_Valid_3_delay_28_10;
    io_A_Valid_3_delay_30_8 <= io_A_Valid_3_delay_29_9;
    io_A_Valid_3_delay_31_7 <= io_A_Valid_3_delay_30_8;
    io_A_Valid_3_delay_32_6 <= io_A_Valid_3_delay_31_7;
    io_A_Valid_3_delay_33_5 <= io_A_Valid_3_delay_32_6;
    io_A_Valid_3_delay_34_4 <= io_A_Valid_3_delay_33_5;
    io_A_Valid_3_delay_35_3 <= io_A_Valid_3_delay_34_4;
    io_A_Valid_3_delay_36_2 <= io_A_Valid_3_delay_35_3;
    io_A_Valid_3_delay_37_1 <= io_A_Valid_3_delay_36_2;
    io_A_Valid_3_delay_38 <= io_A_Valid_3_delay_37_1;
    io_B_Valid_38_delay_1_2 <= io_B_Valid_38;
    io_B_Valid_38_delay_2_1 <= io_B_Valid_38_delay_1_2;
    io_B_Valid_38_delay_3 <= io_B_Valid_38_delay_2_1;
    io_A_Valid_3_delay_1_38 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_37 <= io_A_Valid_3_delay_1_38;
    io_A_Valid_3_delay_3_36 <= io_A_Valid_3_delay_2_37;
    io_A_Valid_3_delay_4_35 <= io_A_Valid_3_delay_3_36;
    io_A_Valid_3_delay_5_34 <= io_A_Valid_3_delay_4_35;
    io_A_Valid_3_delay_6_33 <= io_A_Valid_3_delay_5_34;
    io_A_Valid_3_delay_7_32 <= io_A_Valid_3_delay_6_33;
    io_A_Valid_3_delay_8_31 <= io_A_Valid_3_delay_7_32;
    io_A_Valid_3_delay_9_30 <= io_A_Valid_3_delay_8_31;
    io_A_Valid_3_delay_10_29 <= io_A_Valid_3_delay_9_30;
    io_A_Valid_3_delay_11_28 <= io_A_Valid_3_delay_10_29;
    io_A_Valid_3_delay_12_27 <= io_A_Valid_3_delay_11_28;
    io_A_Valid_3_delay_13_26 <= io_A_Valid_3_delay_12_27;
    io_A_Valid_3_delay_14_25 <= io_A_Valid_3_delay_13_26;
    io_A_Valid_3_delay_15_24 <= io_A_Valid_3_delay_14_25;
    io_A_Valid_3_delay_16_23 <= io_A_Valid_3_delay_15_24;
    io_A_Valid_3_delay_17_22 <= io_A_Valid_3_delay_16_23;
    io_A_Valid_3_delay_18_21 <= io_A_Valid_3_delay_17_22;
    io_A_Valid_3_delay_19_20 <= io_A_Valid_3_delay_18_21;
    io_A_Valid_3_delay_20_19 <= io_A_Valid_3_delay_19_20;
    io_A_Valid_3_delay_21_18 <= io_A_Valid_3_delay_20_19;
    io_A_Valid_3_delay_22_17 <= io_A_Valid_3_delay_21_18;
    io_A_Valid_3_delay_23_16 <= io_A_Valid_3_delay_22_17;
    io_A_Valid_3_delay_24_15 <= io_A_Valid_3_delay_23_16;
    io_A_Valid_3_delay_25_14 <= io_A_Valid_3_delay_24_15;
    io_A_Valid_3_delay_26_13 <= io_A_Valid_3_delay_25_14;
    io_A_Valid_3_delay_27_12 <= io_A_Valid_3_delay_26_13;
    io_A_Valid_3_delay_28_11 <= io_A_Valid_3_delay_27_12;
    io_A_Valid_3_delay_29_10 <= io_A_Valid_3_delay_28_11;
    io_A_Valid_3_delay_30_9 <= io_A_Valid_3_delay_29_10;
    io_A_Valid_3_delay_31_8 <= io_A_Valid_3_delay_30_9;
    io_A_Valid_3_delay_32_7 <= io_A_Valid_3_delay_31_8;
    io_A_Valid_3_delay_33_6 <= io_A_Valid_3_delay_32_7;
    io_A_Valid_3_delay_34_5 <= io_A_Valid_3_delay_33_6;
    io_A_Valid_3_delay_35_4 <= io_A_Valid_3_delay_34_5;
    io_A_Valid_3_delay_36_3 <= io_A_Valid_3_delay_35_4;
    io_A_Valid_3_delay_37_2 <= io_A_Valid_3_delay_36_3;
    io_A_Valid_3_delay_38_1 <= io_A_Valid_3_delay_37_2;
    io_A_Valid_3_delay_39 <= io_A_Valid_3_delay_38_1;
    io_B_Valid_39_delay_1_2 <= io_B_Valid_39;
    io_B_Valid_39_delay_2_1 <= io_B_Valid_39_delay_1_2;
    io_B_Valid_39_delay_3 <= io_B_Valid_39_delay_2_1;
    io_A_Valid_3_delay_1_39 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_38 <= io_A_Valid_3_delay_1_39;
    io_A_Valid_3_delay_3_37 <= io_A_Valid_3_delay_2_38;
    io_A_Valid_3_delay_4_36 <= io_A_Valid_3_delay_3_37;
    io_A_Valid_3_delay_5_35 <= io_A_Valid_3_delay_4_36;
    io_A_Valid_3_delay_6_34 <= io_A_Valid_3_delay_5_35;
    io_A_Valid_3_delay_7_33 <= io_A_Valid_3_delay_6_34;
    io_A_Valid_3_delay_8_32 <= io_A_Valid_3_delay_7_33;
    io_A_Valid_3_delay_9_31 <= io_A_Valid_3_delay_8_32;
    io_A_Valid_3_delay_10_30 <= io_A_Valid_3_delay_9_31;
    io_A_Valid_3_delay_11_29 <= io_A_Valid_3_delay_10_30;
    io_A_Valid_3_delay_12_28 <= io_A_Valid_3_delay_11_29;
    io_A_Valid_3_delay_13_27 <= io_A_Valid_3_delay_12_28;
    io_A_Valid_3_delay_14_26 <= io_A_Valid_3_delay_13_27;
    io_A_Valid_3_delay_15_25 <= io_A_Valid_3_delay_14_26;
    io_A_Valid_3_delay_16_24 <= io_A_Valid_3_delay_15_25;
    io_A_Valid_3_delay_17_23 <= io_A_Valid_3_delay_16_24;
    io_A_Valid_3_delay_18_22 <= io_A_Valid_3_delay_17_23;
    io_A_Valid_3_delay_19_21 <= io_A_Valid_3_delay_18_22;
    io_A_Valid_3_delay_20_20 <= io_A_Valid_3_delay_19_21;
    io_A_Valid_3_delay_21_19 <= io_A_Valid_3_delay_20_20;
    io_A_Valid_3_delay_22_18 <= io_A_Valid_3_delay_21_19;
    io_A_Valid_3_delay_23_17 <= io_A_Valid_3_delay_22_18;
    io_A_Valid_3_delay_24_16 <= io_A_Valid_3_delay_23_17;
    io_A_Valid_3_delay_25_15 <= io_A_Valid_3_delay_24_16;
    io_A_Valid_3_delay_26_14 <= io_A_Valid_3_delay_25_15;
    io_A_Valid_3_delay_27_13 <= io_A_Valid_3_delay_26_14;
    io_A_Valid_3_delay_28_12 <= io_A_Valid_3_delay_27_13;
    io_A_Valid_3_delay_29_11 <= io_A_Valid_3_delay_28_12;
    io_A_Valid_3_delay_30_10 <= io_A_Valid_3_delay_29_11;
    io_A_Valid_3_delay_31_9 <= io_A_Valid_3_delay_30_10;
    io_A_Valid_3_delay_32_8 <= io_A_Valid_3_delay_31_9;
    io_A_Valid_3_delay_33_7 <= io_A_Valid_3_delay_32_8;
    io_A_Valid_3_delay_34_6 <= io_A_Valid_3_delay_33_7;
    io_A_Valid_3_delay_35_5 <= io_A_Valid_3_delay_34_6;
    io_A_Valid_3_delay_36_4 <= io_A_Valid_3_delay_35_5;
    io_A_Valid_3_delay_37_3 <= io_A_Valid_3_delay_36_4;
    io_A_Valid_3_delay_38_2 <= io_A_Valid_3_delay_37_3;
    io_A_Valid_3_delay_39_1 <= io_A_Valid_3_delay_38_2;
    io_A_Valid_3_delay_40 <= io_A_Valid_3_delay_39_1;
    io_B_Valid_40_delay_1_2 <= io_B_Valid_40;
    io_B_Valid_40_delay_2_1 <= io_B_Valid_40_delay_1_2;
    io_B_Valid_40_delay_3 <= io_B_Valid_40_delay_2_1;
    io_A_Valid_3_delay_1_40 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_39 <= io_A_Valid_3_delay_1_40;
    io_A_Valid_3_delay_3_38 <= io_A_Valid_3_delay_2_39;
    io_A_Valid_3_delay_4_37 <= io_A_Valid_3_delay_3_38;
    io_A_Valid_3_delay_5_36 <= io_A_Valid_3_delay_4_37;
    io_A_Valid_3_delay_6_35 <= io_A_Valid_3_delay_5_36;
    io_A_Valid_3_delay_7_34 <= io_A_Valid_3_delay_6_35;
    io_A_Valid_3_delay_8_33 <= io_A_Valid_3_delay_7_34;
    io_A_Valid_3_delay_9_32 <= io_A_Valid_3_delay_8_33;
    io_A_Valid_3_delay_10_31 <= io_A_Valid_3_delay_9_32;
    io_A_Valid_3_delay_11_30 <= io_A_Valid_3_delay_10_31;
    io_A_Valid_3_delay_12_29 <= io_A_Valid_3_delay_11_30;
    io_A_Valid_3_delay_13_28 <= io_A_Valid_3_delay_12_29;
    io_A_Valid_3_delay_14_27 <= io_A_Valid_3_delay_13_28;
    io_A_Valid_3_delay_15_26 <= io_A_Valid_3_delay_14_27;
    io_A_Valid_3_delay_16_25 <= io_A_Valid_3_delay_15_26;
    io_A_Valid_3_delay_17_24 <= io_A_Valid_3_delay_16_25;
    io_A_Valid_3_delay_18_23 <= io_A_Valid_3_delay_17_24;
    io_A_Valid_3_delay_19_22 <= io_A_Valid_3_delay_18_23;
    io_A_Valid_3_delay_20_21 <= io_A_Valid_3_delay_19_22;
    io_A_Valid_3_delay_21_20 <= io_A_Valid_3_delay_20_21;
    io_A_Valid_3_delay_22_19 <= io_A_Valid_3_delay_21_20;
    io_A_Valid_3_delay_23_18 <= io_A_Valid_3_delay_22_19;
    io_A_Valid_3_delay_24_17 <= io_A_Valid_3_delay_23_18;
    io_A_Valid_3_delay_25_16 <= io_A_Valid_3_delay_24_17;
    io_A_Valid_3_delay_26_15 <= io_A_Valid_3_delay_25_16;
    io_A_Valid_3_delay_27_14 <= io_A_Valid_3_delay_26_15;
    io_A_Valid_3_delay_28_13 <= io_A_Valid_3_delay_27_14;
    io_A_Valid_3_delay_29_12 <= io_A_Valid_3_delay_28_13;
    io_A_Valid_3_delay_30_11 <= io_A_Valid_3_delay_29_12;
    io_A_Valid_3_delay_31_10 <= io_A_Valid_3_delay_30_11;
    io_A_Valid_3_delay_32_9 <= io_A_Valid_3_delay_31_10;
    io_A_Valid_3_delay_33_8 <= io_A_Valid_3_delay_32_9;
    io_A_Valid_3_delay_34_7 <= io_A_Valid_3_delay_33_8;
    io_A_Valid_3_delay_35_6 <= io_A_Valid_3_delay_34_7;
    io_A_Valid_3_delay_36_5 <= io_A_Valid_3_delay_35_6;
    io_A_Valid_3_delay_37_4 <= io_A_Valid_3_delay_36_5;
    io_A_Valid_3_delay_38_3 <= io_A_Valid_3_delay_37_4;
    io_A_Valid_3_delay_39_2 <= io_A_Valid_3_delay_38_3;
    io_A_Valid_3_delay_40_1 <= io_A_Valid_3_delay_39_2;
    io_A_Valid_3_delay_41 <= io_A_Valid_3_delay_40_1;
    io_B_Valid_41_delay_1_2 <= io_B_Valid_41;
    io_B_Valid_41_delay_2_1 <= io_B_Valid_41_delay_1_2;
    io_B_Valid_41_delay_3 <= io_B_Valid_41_delay_2_1;
    io_A_Valid_3_delay_1_41 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_40 <= io_A_Valid_3_delay_1_41;
    io_A_Valid_3_delay_3_39 <= io_A_Valid_3_delay_2_40;
    io_A_Valid_3_delay_4_38 <= io_A_Valid_3_delay_3_39;
    io_A_Valid_3_delay_5_37 <= io_A_Valid_3_delay_4_38;
    io_A_Valid_3_delay_6_36 <= io_A_Valid_3_delay_5_37;
    io_A_Valid_3_delay_7_35 <= io_A_Valid_3_delay_6_36;
    io_A_Valid_3_delay_8_34 <= io_A_Valid_3_delay_7_35;
    io_A_Valid_3_delay_9_33 <= io_A_Valid_3_delay_8_34;
    io_A_Valid_3_delay_10_32 <= io_A_Valid_3_delay_9_33;
    io_A_Valid_3_delay_11_31 <= io_A_Valid_3_delay_10_32;
    io_A_Valid_3_delay_12_30 <= io_A_Valid_3_delay_11_31;
    io_A_Valid_3_delay_13_29 <= io_A_Valid_3_delay_12_30;
    io_A_Valid_3_delay_14_28 <= io_A_Valid_3_delay_13_29;
    io_A_Valid_3_delay_15_27 <= io_A_Valid_3_delay_14_28;
    io_A_Valid_3_delay_16_26 <= io_A_Valid_3_delay_15_27;
    io_A_Valid_3_delay_17_25 <= io_A_Valid_3_delay_16_26;
    io_A_Valid_3_delay_18_24 <= io_A_Valid_3_delay_17_25;
    io_A_Valid_3_delay_19_23 <= io_A_Valid_3_delay_18_24;
    io_A_Valid_3_delay_20_22 <= io_A_Valid_3_delay_19_23;
    io_A_Valid_3_delay_21_21 <= io_A_Valid_3_delay_20_22;
    io_A_Valid_3_delay_22_20 <= io_A_Valid_3_delay_21_21;
    io_A_Valid_3_delay_23_19 <= io_A_Valid_3_delay_22_20;
    io_A_Valid_3_delay_24_18 <= io_A_Valid_3_delay_23_19;
    io_A_Valid_3_delay_25_17 <= io_A_Valid_3_delay_24_18;
    io_A_Valid_3_delay_26_16 <= io_A_Valid_3_delay_25_17;
    io_A_Valid_3_delay_27_15 <= io_A_Valid_3_delay_26_16;
    io_A_Valid_3_delay_28_14 <= io_A_Valid_3_delay_27_15;
    io_A_Valid_3_delay_29_13 <= io_A_Valid_3_delay_28_14;
    io_A_Valid_3_delay_30_12 <= io_A_Valid_3_delay_29_13;
    io_A_Valid_3_delay_31_11 <= io_A_Valid_3_delay_30_12;
    io_A_Valid_3_delay_32_10 <= io_A_Valid_3_delay_31_11;
    io_A_Valid_3_delay_33_9 <= io_A_Valid_3_delay_32_10;
    io_A_Valid_3_delay_34_8 <= io_A_Valid_3_delay_33_9;
    io_A_Valid_3_delay_35_7 <= io_A_Valid_3_delay_34_8;
    io_A_Valid_3_delay_36_6 <= io_A_Valid_3_delay_35_7;
    io_A_Valid_3_delay_37_5 <= io_A_Valid_3_delay_36_6;
    io_A_Valid_3_delay_38_4 <= io_A_Valid_3_delay_37_5;
    io_A_Valid_3_delay_39_3 <= io_A_Valid_3_delay_38_4;
    io_A_Valid_3_delay_40_2 <= io_A_Valid_3_delay_39_3;
    io_A_Valid_3_delay_41_1 <= io_A_Valid_3_delay_40_2;
    io_A_Valid_3_delay_42 <= io_A_Valid_3_delay_41_1;
    io_B_Valid_42_delay_1_2 <= io_B_Valid_42;
    io_B_Valid_42_delay_2_1 <= io_B_Valid_42_delay_1_2;
    io_B_Valid_42_delay_3 <= io_B_Valid_42_delay_2_1;
    io_A_Valid_3_delay_1_42 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_41 <= io_A_Valid_3_delay_1_42;
    io_A_Valid_3_delay_3_40 <= io_A_Valid_3_delay_2_41;
    io_A_Valid_3_delay_4_39 <= io_A_Valid_3_delay_3_40;
    io_A_Valid_3_delay_5_38 <= io_A_Valid_3_delay_4_39;
    io_A_Valid_3_delay_6_37 <= io_A_Valid_3_delay_5_38;
    io_A_Valid_3_delay_7_36 <= io_A_Valid_3_delay_6_37;
    io_A_Valid_3_delay_8_35 <= io_A_Valid_3_delay_7_36;
    io_A_Valid_3_delay_9_34 <= io_A_Valid_3_delay_8_35;
    io_A_Valid_3_delay_10_33 <= io_A_Valid_3_delay_9_34;
    io_A_Valid_3_delay_11_32 <= io_A_Valid_3_delay_10_33;
    io_A_Valid_3_delay_12_31 <= io_A_Valid_3_delay_11_32;
    io_A_Valid_3_delay_13_30 <= io_A_Valid_3_delay_12_31;
    io_A_Valid_3_delay_14_29 <= io_A_Valid_3_delay_13_30;
    io_A_Valid_3_delay_15_28 <= io_A_Valid_3_delay_14_29;
    io_A_Valid_3_delay_16_27 <= io_A_Valid_3_delay_15_28;
    io_A_Valid_3_delay_17_26 <= io_A_Valid_3_delay_16_27;
    io_A_Valid_3_delay_18_25 <= io_A_Valid_3_delay_17_26;
    io_A_Valid_3_delay_19_24 <= io_A_Valid_3_delay_18_25;
    io_A_Valid_3_delay_20_23 <= io_A_Valid_3_delay_19_24;
    io_A_Valid_3_delay_21_22 <= io_A_Valid_3_delay_20_23;
    io_A_Valid_3_delay_22_21 <= io_A_Valid_3_delay_21_22;
    io_A_Valid_3_delay_23_20 <= io_A_Valid_3_delay_22_21;
    io_A_Valid_3_delay_24_19 <= io_A_Valid_3_delay_23_20;
    io_A_Valid_3_delay_25_18 <= io_A_Valid_3_delay_24_19;
    io_A_Valid_3_delay_26_17 <= io_A_Valid_3_delay_25_18;
    io_A_Valid_3_delay_27_16 <= io_A_Valid_3_delay_26_17;
    io_A_Valid_3_delay_28_15 <= io_A_Valid_3_delay_27_16;
    io_A_Valid_3_delay_29_14 <= io_A_Valid_3_delay_28_15;
    io_A_Valid_3_delay_30_13 <= io_A_Valid_3_delay_29_14;
    io_A_Valid_3_delay_31_12 <= io_A_Valid_3_delay_30_13;
    io_A_Valid_3_delay_32_11 <= io_A_Valid_3_delay_31_12;
    io_A_Valid_3_delay_33_10 <= io_A_Valid_3_delay_32_11;
    io_A_Valid_3_delay_34_9 <= io_A_Valid_3_delay_33_10;
    io_A_Valid_3_delay_35_8 <= io_A_Valid_3_delay_34_9;
    io_A_Valid_3_delay_36_7 <= io_A_Valid_3_delay_35_8;
    io_A_Valid_3_delay_37_6 <= io_A_Valid_3_delay_36_7;
    io_A_Valid_3_delay_38_5 <= io_A_Valid_3_delay_37_6;
    io_A_Valid_3_delay_39_4 <= io_A_Valid_3_delay_38_5;
    io_A_Valid_3_delay_40_3 <= io_A_Valid_3_delay_39_4;
    io_A_Valid_3_delay_41_2 <= io_A_Valid_3_delay_40_3;
    io_A_Valid_3_delay_42_1 <= io_A_Valid_3_delay_41_2;
    io_A_Valid_3_delay_43 <= io_A_Valid_3_delay_42_1;
    io_B_Valid_43_delay_1_2 <= io_B_Valid_43;
    io_B_Valid_43_delay_2_1 <= io_B_Valid_43_delay_1_2;
    io_B_Valid_43_delay_3 <= io_B_Valid_43_delay_2_1;
    io_A_Valid_3_delay_1_43 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_42 <= io_A_Valid_3_delay_1_43;
    io_A_Valid_3_delay_3_41 <= io_A_Valid_3_delay_2_42;
    io_A_Valid_3_delay_4_40 <= io_A_Valid_3_delay_3_41;
    io_A_Valid_3_delay_5_39 <= io_A_Valid_3_delay_4_40;
    io_A_Valid_3_delay_6_38 <= io_A_Valid_3_delay_5_39;
    io_A_Valid_3_delay_7_37 <= io_A_Valid_3_delay_6_38;
    io_A_Valid_3_delay_8_36 <= io_A_Valid_3_delay_7_37;
    io_A_Valid_3_delay_9_35 <= io_A_Valid_3_delay_8_36;
    io_A_Valid_3_delay_10_34 <= io_A_Valid_3_delay_9_35;
    io_A_Valid_3_delay_11_33 <= io_A_Valid_3_delay_10_34;
    io_A_Valid_3_delay_12_32 <= io_A_Valid_3_delay_11_33;
    io_A_Valid_3_delay_13_31 <= io_A_Valid_3_delay_12_32;
    io_A_Valid_3_delay_14_30 <= io_A_Valid_3_delay_13_31;
    io_A_Valid_3_delay_15_29 <= io_A_Valid_3_delay_14_30;
    io_A_Valid_3_delay_16_28 <= io_A_Valid_3_delay_15_29;
    io_A_Valid_3_delay_17_27 <= io_A_Valid_3_delay_16_28;
    io_A_Valid_3_delay_18_26 <= io_A_Valid_3_delay_17_27;
    io_A_Valid_3_delay_19_25 <= io_A_Valid_3_delay_18_26;
    io_A_Valid_3_delay_20_24 <= io_A_Valid_3_delay_19_25;
    io_A_Valid_3_delay_21_23 <= io_A_Valid_3_delay_20_24;
    io_A_Valid_3_delay_22_22 <= io_A_Valid_3_delay_21_23;
    io_A_Valid_3_delay_23_21 <= io_A_Valid_3_delay_22_22;
    io_A_Valid_3_delay_24_20 <= io_A_Valid_3_delay_23_21;
    io_A_Valid_3_delay_25_19 <= io_A_Valid_3_delay_24_20;
    io_A_Valid_3_delay_26_18 <= io_A_Valid_3_delay_25_19;
    io_A_Valid_3_delay_27_17 <= io_A_Valid_3_delay_26_18;
    io_A_Valid_3_delay_28_16 <= io_A_Valid_3_delay_27_17;
    io_A_Valid_3_delay_29_15 <= io_A_Valid_3_delay_28_16;
    io_A_Valid_3_delay_30_14 <= io_A_Valid_3_delay_29_15;
    io_A_Valid_3_delay_31_13 <= io_A_Valid_3_delay_30_14;
    io_A_Valid_3_delay_32_12 <= io_A_Valid_3_delay_31_13;
    io_A_Valid_3_delay_33_11 <= io_A_Valid_3_delay_32_12;
    io_A_Valid_3_delay_34_10 <= io_A_Valid_3_delay_33_11;
    io_A_Valid_3_delay_35_9 <= io_A_Valid_3_delay_34_10;
    io_A_Valid_3_delay_36_8 <= io_A_Valid_3_delay_35_9;
    io_A_Valid_3_delay_37_7 <= io_A_Valid_3_delay_36_8;
    io_A_Valid_3_delay_38_6 <= io_A_Valid_3_delay_37_7;
    io_A_Valid_3_delay_39_5 <= io_A_Valid_3_delay_38_6;
    io_A_Valid_3_delay_40_4 <= io_A_Valid_3_delay_39_5;
    io_A_Valid_3_delay_41_3 <= io_A_Valid_3_delay_40_4;
    io_A_Valid_3_delay_42_2 <= io_A_Valid_3_delay_41_3;
    io_A_Valid_3_delay_43_1 <= io_A_Valid_3_delay_42_2;
    io_A_Valid_3_delay_44 <= io_A_Valid_3_delay_43_1;
    io_B_Valid_44_delay_1_2 <= io_B_Valid_44;
    io_B_Valid_44_delay_2_1 <= io_B_Valid_44_delay_1_2;
    io_B_Valid_44_delay_3 <= io_B_Valid_44_delay_2_1;
    io_A_Valid_3_delay_1_44 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_43 <= io_A_Valid_3_delay_1_44;
    io_A_Valid_3_delay_3_42 <= io_A_Valid_3_delay_2_43;
    io_A_Valid_3_delay_4_41 <= io_A_Valid_3_delay_3_42;
    io_A_Valid_3_delay_5_40 <= io_A_Valid_3_delay_4_41;
    io_A_Valid_3_delay_6_39 <= io_A_Valid_3_delay_5_40;
    io_A_Valid_3_delay_7_38 <= io_A_Valid_3_delay_6_39;
    io_A_Valid_3_delay_8_37 <= io_A_Valid_3_delay_7_38;
    io_A_Valid_3_delay_9_36 <= io_A_Valid_3_delay_8_37;
    io_A_Valid_3_delay_10_35 <= io_A_Valid_3_delay_9_36;
    io_A_Valid_3_delay_11_34 <= io_A_Valid_3_delay_10_35;
    io_A_Valid_3_delay_12_33 <= io_A_Valid_3_delay_11_34;
    io_A_Valid_3_delay_13_32 <= io_A_Valid_3_delay_12_33;
    io_A_Valid_3_delay_14_31 <= io_A_Valid_3_delay_13_32;
    io_A_Valid_3_delay_15_30 <= io_A_Valid_3_delay_14_31;
    io_A_Valid_3_delay_16_29 <= io_A_Valid_3_delay_15_30;
    io_A_Valid_3_delay_17_28 <= io_A_Valid_3_delay_16_29;
    io_A_Valid_3_delay_18_27 <= io_A_Valid_3_delay_17_28;
    io_A_Valid_3_delay_19_26 <= io_A_Valid_3_delay_18_27;
    io_A_Valid_3_delay_20_25 <= io_A_Valid_3_delay_19_26;
    io_A_Valid_3_delay_21_24 <= io_A_Valid_3_delay_20_25;
    io_A_Valid_3_delay_22_23 <= io_A_Valid_3_delay_21_24;
    io_A_Valid_3_delay_23_22 <= io_A_Valid_3_delay_22_23;
    io_A_Valid_3_delay_24_21 <= io_A_Valid_3_delay_23_22;
    io_A_Valid_3_delay_25_20 <= io_A_Valid_3_delay_24_21;
    io_A_Valid_3_delay_26_19 <= io_A_Valid_3_delay_25_20;
    io_A_Valid_3_delay_27_18 <= io_A_Valid_3_delay_26_19;
    io_A_Valid_3_delay_28_17 <= io_A_Valid_3_delay_27_18;
    io_A_Valid_3_delay_29_16 <= io_A_Valid_3_delay_28_17;
    io_A_Valid_3_delay_30_15 <= io_A_Valid_3_delay_29_16;
    io_A_Valid_3_delay_31_14 <= io_A_Valid_3_delay_30_15;
    io_A_Valid_3_delay_32_13 <= io_A_Valid_3_delay_31_14;
    io_A_Valid_3_delay_33_12 <= io_A_Valid_3_delay_32_13;
    io_A_Valid_3_delay_34_11 <= io_A_Valid_3_delay_33_12;
    io_A_Valid_3_delay_35_10 <= io_A_Valid_3_delay_34_11;
    io_A_Valid_3_delay_36_9 <= io_A_Valid_3_delay_35_10;
    io_A_Valid_3_delay_37_8 <= io_A_Valid_3_delay_36_9;
    io_A_Valid_3_delay_38_7 <= io_A_Valid_3_delay_37_8;
    io_A_Valid_3_delay_39_6 <= io_A_Valid_3_delay_38_7;
    io_A_Valid_3_delay_40_5 <= io_A_Valid_3_delay_39_6;
    io_A_Valid_3_delay_41_4 <= io_A_Valid_3_delay_40_5;
    io_A_Valid_3_delay_42_3 <= io_A_Valid_3_delay_41_4;
    io_A_Valid_3_delay_43_2 <= io_A_Valid_3_delay_42_3;
    io_A_Valid_3_delay_44_1 <= io_A_Valid_3_delay_43_2;
    io_A_Valid_3_delay_45 <= io_A_Valid_3_delay_44_1;
    io_B_Valid_45_delay_1_2 <= io_B_Valid_45;
    io_B_Valid_45_delay_2_1 <= io_B_Valid_45_delay_1_2;
    io_B_Valid_45_delay_3 <= io_B_Valid_45_delay_2_1;
    io_A_Valid_3_delay_1_45 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_44 <= io_A_Valid_3_delay_1_45;
    io_A_Valid_3_delay_3_43 <= io_A_Valid_3_delay_2_44;
    io_A_Valid_3_delay_4_42 <= io_A_Valid_3_delay_3_43;
    io_A_Valid_3_delay_5_41 <= io_A_Valid_3_delay_4_42;
    io_A_Valid_3_delay_6_40 <= io_A_Valid_3_delay_5_41;
    io_A_Valid_3_delay_7_39 <= io_A_Valid_3_delay_6_40;
    io_A_Valid_3_delay_8_38 <= io_A_Valid_3_delay_7_39;
    io_A_Valid_3_delay_9_37 <= io_A_Valid_3_delay_8_38;
    io_A_Valid_3_delay_10_36 <= io_A_Valid_3_delay_9_37;
    io_A_Valid_3_delay_11_35 <= io_A_Valid_3_delay_10_36;
    io_A_Valid_3_delay_12_34 <= io_A_Valid_3_delay_11_35;
    io_A_Valid_3_delay_13_33 <= io_A_Valid_3_delay_12_34;
    io_A_Valid_3_delay_14_32 <= io_A_Valid_3_delay_13_33;
    io_A_Valid_3_delay_15_31 <= io_A_Valid_3_delay_14_32;
    io_A_Valid_3_delay_16_30 <= io_A_Valid_3_delay_15_31;
    io_A_Valid_3_delay_17_29 <= io_A_Valid_3_delay_16_30;
    io_A_Valid_3_delay_18_28 <= io_A_Valid_3_delay_17_29;
    io_A_Valid_3_delay_19_27 <= io_A_Valid_3_delay_18_28;
    io_A_Valid_3_delay_20_26 <= io_A_Valid_3_delay_19_27;
    io_A_Valid_3_delay_21_25 <= io_A_Valid_3_delay_20_26;
    io_A_Valid_3_delay_22_24 <= io_A_Valid_3_delay_21_25;
    io_A_Valid_3_delay_23_23 <= io_A_Valid_3_delay_22_24;
    io_A_Valid_3_delay_24_22 <= io_A_Valid_3_delay_23_23;
    io_A_Valid_3_delay_25_21 <= io_A_Valid_3_delay_24_22;
    io_A_Valid_3_delay_26_20 <= io_A_Valid_3_delay_25_21;
    io_A_Valid_3_delay_27_19 <= io_A_Valid_3_delay_26_20;
    io_A_Valid_3_delay_28_18 <= io_A_Valid_3_delay_27_19;
    io_A_Valid_3_delay_29_17 <= io_A_Valid_3_delay_28_18;
    io_A_Valid_3_delay_30_16 <= io_A_Valid_3_delay_29_17;
    io_A_Valid_3_delay_31_15 <= io_A_Valid_3_delay_30_16;
    io_A_Valid_3_delay_32_14 <= io_A_Valid_3_delay_31_15;
    io_A_Valid_3_delay_33_13 <= io_A_Valid_3_delay_32_14;
    io_A_Valid_3_delay_34_12 <= io_A_Valid_3_delay_33_13;
    io_A_Valid_3_delay_35_11 <= io_A_Valid_3_delay_34_12;
    io_A_Valid_3_delay_36_10 <= io_A_Valid_3_delay_35_11;
    io_A_Valid_3_delay_37_9 <= io_A_Valid_3_delay_36_10;
    io_A_Valid_3_delay_38_8 <= io_A_Valid_3_delay_37_9;
    io_A_Valid_3_delay_39_7 <= io_A_Valid_3_delay_38_8;
    io_A_Valid_3_delay_40_6 <= io_A_Valid_3_delay_39_7;
    io_A_Valid_3_delay_41_5 <= io_A_Valid_3_delay_40_6;
    io_A_Valid_3_delay_42_4 <= io_A_Valid_3_delay_41_5;
    io_A_Valid_3_delay_43_3 <= io_A_Valid_3_delay_42_4;
    io_A_Valid_3_delay_44_2 <= io_A_Valid_3_delay_43_3;
    io_A_Valid_3_delay_45_1 <= io_A_Valid_3_delay_44_2;
    io_A_Valid_3_delay_46 <= io_A_Valid_3_delay_45_1;
    io_B_Valid_46_delay_1_2 <= io_B_Valid_46;
    io_B_Valid_46_delay_2_1 <= io_B_Valid_46_delay_1_2;
    io_B_Valid_46_delay_3 <= io_B_Valid_46_delay_2_1;
    io_A_Valid_3_delay_1_46 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_45 <= io_A_Valid_3_delay_1_46;
    io_A_Valid_3_delay_3_44 <= io_A_Valid_3_delay_2_45;
    io_A_Valid_3_delay_4_43 <= io_A_Valid_3_delay_3_44;
    io_A_Valid_3_delay_5_42 <= io_A_Valid_3_delay_4_43;
    io_A_Valid_3_delay_6_41 <= io_A_Valid_3_delay_5_42;
    io_A_Valid_3_delay_7_40 <= io_A_Valid_3_delay_6_41;
    io_A_Valid_3_delay_8_39 <= io_A_Valid_3_delay_7_40;
    io_A_Valid_3_delay_9_38 <= io_A_Valid_3_delay_8_39;
    io_A_Valid_3_delay_10_37 <= io_A_Valid_3_delay_9_38;
    io_A_Valid_3_delay_11_36 <= io_A_Valid_3_delay_10_37;
    io_A_Valid_3_delay_12_35 <= io_A_Valid_3_delay_11_36;
    io_A_Valid_3_delay_13_34 <= io_A_Valid_3_delay_12_35;
    io_A_Valid_3_delay_14_33 <= io_A_Valid_3_delay_13_34;
    io_A_Valid_3_delay_15_32 <= io_A_Valid_3_delay_14_33;
    io_A_Valid_3_delay_16_31 <= io_A_Valid_3_delay_15_32;
    io_A_Valid_3_delay_17_30 <= io_A_Valid_3_delay_16_31;
    io_A_Valid_3_delay_18_29 <= io_A_Valid_3_delay_17_30;
    io_A_Valid_3_delay_19_28 <= io_A_Valid_3_delay_18_29;
    io_A_Valid_3_delay_20_27 <= io_A_Valid_3_delay_19_28;
    io_A_Valid_3_delay_21_26 <= io_A_Valid_3_delay_20_27;
    io_A_Valid_3_delay_22_25 <= io_A_Valid_3_delay_21_26;
    io_A_Valid_3_delay_23_24 <= io_A_Valid_3_delay_22_25;
    io_A_Valid_3_delay_24_23 <= io_A_Valid_3_delay_23_24;
    io_A_Valid_3_delay_25_22 <= io_A_Valid_3_delay_24_23;
    io_A_Valid_3_delay_26_21 <= io_A_Valid_3_delay_25_22;
    io_A_Valid_3_delay_27_20 <= io_A_Valid_3_delay_26_21;
    io_A_Valid_3_delay_28_19 <= io_A_Valid_3_delay_27_20;
    io_A_Valid_3_delay_29_18 <= io_A_Valid_3_delay_28_19;
    io_A_Valid_3_delay_30_17 <= io_A_Valid_3_delay_29_18;
    io_A_Valid_3_delay_31_16 <= io_A_Valid_3_delay_30_17;
    io_A_Valid_3_delay_32_15 <= io_A_Valid_3_delay_31_16;
    io_A_Valid_3_delay_33_14 <= io_A_Valid_3_delay_32_15;
    io_A_Valid_3_delay_34_13 <= io_A_Valid_3_delay_33_14;
    io_A_Valid_3_delay_35_12 <= io_A_Valid_3_delay_34_13;
    io_A_Valid_3_delay_36_11 <= io_A_Valid_3_delay_35_12;
    io_A_Valid_3_delay_37_10 <= io_A_Valid_3_delay_36_11;
    io_A_Valid_3_delay_38_9 <= io_A_Valid_3_delay_37_10;
    io_A_Valid_3_delay_39_8 <= io_A_Valid_3_delay_38_9;
    io_A_Valid_3_delay_40_7 <= io_A_Valid_3_delay_39_8;
    io_A_Valid_3_delay_41_6 <= io_A_Valid_3_delay_40_7;
    io_A_Valid_3_delay_42_5 <= io_A_Valid_3_delay_41_6;
    io_A_Valid_3_delay_43_4 <= io_A_Valid_3_delay_42_5;
    io_A_Valid_3_delay_44_3 <= io_A_Valid_3_delay_43_4;
    io_A_Valid_3_delay_45_2 <= io_A_Valid_3_delay_44_3;
    io_A_Valid_3_delay_46_1 <= io_A_Valid_3_delay_45_2;
    io_A_Valid_3_delay_47 <= io_A_Valid_3_delay_46_1;
    io_B_Valid_47_delay_1_2 <= io_B_Valid_47;
    io_B_Valid_47_delay_2_1 <= io_B_Valid_47_delay_1_2;
    io_B_Valid_47_delay_3 <= io_B_Valid_47_delay_2_1;
    io_A_Valid_3_delay_1_47 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_46 <= io_A_Valid_3_delay_1_47;
    io_A_Valid_3_delay_3_45 <= io_A_Valid_3_delay_2_46;
    io_A_Valid_3_delay_4_44 <= io_A_Valid_3_delay_3_45;
    io_A_Valid_3_delay_5_43 <= io_A_Valid_3_delay_4_44;
    io_A_Valid_3_delay_6_42 <= io_A_Valid_3_delay_5_43;
    io_A_Valid_3_delay_7_41 <= io_A_Valid_3_delay_6_42;
    io_A_Valid_3_delay_8_40 <= io_A_Valid_3_delay_7_41;
    io_A_Valid_3_delay_9_39 <= io_A_Valid_3_delay_8_40;
    io_A_Valid_3_delay_10_38 <= io_A_Valid_3_delay_9_39;
    io_A_Valid_3_delay_11_37 <= io_A_Valid_3_delay_10_38;
    io_A_Valid_3_delay_12_36 <= io_A_Valid_3_delay_11_37;
    io_A_Valid_3_delay_13_35 <= io_A_Valid_3_delay_12_36;
    io_A_Valid_3_delay_14_34 <= io_A_Valid_3_delay_13_35;
    io_A_Valid_3_delay_15_33 <= io_A_Valid_3_delay_14_34;
    io_A_Valid_3_delay_16_32 <= io_A_Valid_3_delay_15_33;
    io_A_Valid_3_delay_17_31 <= io_A_Valid_3_delay_16_32;
    io_A_Valid_3_delay_18_30 <= io_A_Valid_3_delay_17_31;
    io_A_Valid_3_delay_19_29 <= io_A_Valid_3_delay_18_30;
    io_A_Valid_3_delay_20_28 <= io_A_Valid_3_delay_19_29;
    io_A_Valid_3_delay_21_27 <= io_A_Valid_3_delay_20_28;
    io_A_Valid_3_delay_22_26 <= io_A_Valid_3_delay_21_27;
    io_A_Valid_3_delay_23_25 <= io_A_Valid_3_delay_22_26;
    io_A_Valid_3_delay_24_24 <= io_A_Valid_3_delay_23_25;
    io_A_Valid_3_delay_25_23 <= io_A_Valid_3_delay_24_24;
    io_A_Valid_3_delay_26_22 <= io_A_Valid_3_delay_25_23;
    io_A_Valid_3_delay_27_21 <= io_A_Valid_3_delay_26_22;
    io_A_Valid_3_delay_28_20 <= io_A_Valid_3_delay_27_21;
    io_A_Valid_3_delay_29_19 <= io_A_Valid_3_delay_28_20;
    io_A_Valid_3_delay_30_18 <= io_A_Valid_3_delay_29_19;
    io_A_Valid_3_delay_31_17 <= io_A_Valid_3_delay_30_18;
    io_A_Valid_3_delay_32_16 <= io_A_Valid_3_delay_31_17;
    io_A_Valid_3_delay_33_15 <= io_A_Valid_3_delay_32_16;
    io_A_Valid_3_delay_34_14 <= io_A_Valid_3_delay_33_15;
    io_A_Valid_3_delay_35_13 <= io_A_Valid_3_delay_34_14;
    io_A_Valid_3_delay_36_12 <= io_A_Valid_3_delay_35_13;
    io_A_Valid_3_delay_37_11 <= io_A_Valid_3_delay_36_12;
    io_A_Valid_3_delay_38_10 <= io_A_Valid_3_delay_37_11;
    io_A_Valid_3_delay_39_9 <= io_A_Valid_3_delay_38_10;
    io_A_Valid_3_delay_40_8 <= io_A_Valid_3_delay_39_9;
    io_A_Valid_3_delay_41_7 <= io_A_Valid_3_delay_40_8;
    io_A_Valid_3_delay_42_6 <= io_A_Valid_3_delay_41_7;
    io_A_Valid_3_delay_43_5 <= io_A_Valid_3_delay_42_6;
    io_A_Valid_3_delay_44_4 <= io_A_Valid_3_delay_43_5;
    io_A_Valid_3_delay_45_3 <= io_A_Valid_3_delay_44_4;
    io_A_Valid_3_delay_46_2 <= io_A_Valid_3_delay_45_3;
    io_A_Valid_3_delay_47_1 <= io_A_Valid_3_delay_46_2;
    io_A_Valid_3_delay_48 <= io_A_Valid_3_delay_47_1;
    io_B_Valid_48_delay_1_2 <= io_B_Valid_48;
    io_B_Valid_48_delay_2_1 <= io_B_Valid_48_delay_1_2;
    io_B_Valid_48_delay_3 <= io_B_Valid_48_delay_2_1;
    io_A_Valid_3_delay_1_48 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_47 <= io_A_Valid_3_delay_1_48;
    io_A_Valid_3_delay_3_46 <= io_A_Valid_3_delay_2_47;
    io_A_Valid_3_delay_4_45 <= io_A_Valid_3_delay_3_46;
    io_A_Valid_3_delay_5_44 <= io_A_Valid_3_delay_4_45;
    io_A_Valid_3_delay_6_43 <= io_A_Valid_3_delay_5_44;
    io_A_Valid_3_delay_7_42 <= io_A_Valid_3_delay_6_43;
    io_A_Valid_3_delay_8_41 <= io_A_Valid_3_delay_7_42;
    io_A_Valid_3_delay_9_40 <= io_A_Valid_3_delay_8_41;
    io_A_Valid_3_delay_10_39 <= io_A_Valid_3_delay_9_40;
    io_A_Valid_3_delay_11_38 <= io_A_Valid_3_delay_10_39;
    io_A_Valid_3_delay_12_37 <= io_A_Valid_3_delay_11_38;
    io_A_Valid_3_delay_13_36 <= io_A_Valid_3_delay_12_37;
    io_A_Valid_3_delay_14_35 <= io_A_Valid_3_delay_13_36;
    io_A_Valid_3_delay_15_34 <= io_A_Valid_3_delay_14_35;
    io_A_Valid_3_delay_16_33 <= io_A_Valid_3_delay_15_34;
    io_A_Valid_3_delay_17_32 <= io_A_Valid_3_delay_16_33;
    io_A_Valid_3_delay_18_31 <= io_A_Valid_3_delay_17_32;
    io_A_Valid_3_delay_19_30 <= io_A_Valid_3_delay_18_31;
    io_A_Valid_3_delay_20_29 <= io_A_Valid_3_delay_19_30;
    io_A_Valid_3_delay_21_28 <= io_A_Valid_3_delay_20_29;
    io_A_Valid_3_delay_22_27 <= io_A_Valid_3_delay_21_28;
    io_A_Valid_3_delay_23_26 <= io_A_Valid_3_delay_22_27;
    io_A_Valid_3_delay_24_25 <= io_A_Valid_3_delay_23_26;
    io_A_Valid_3_delay_25_24 <= io_A_Valid_3_delay_24_25;
    io_A_Valid_3_delay_26_23 <= io_A_Valid_3_delay_25_24;
    io_A_Valid_3_delay_27_22 <= io_A_Valid_3_delay_26_23;
    io_A_Valid_3_delay_28_21 <= io_A_Valid_3_delay_27_22;
    io_A_Valid_3_delay_29_20 <= io_A_Valid_3_delay_28_21;
    io_A_Valid_3_delay_30_19 <= io_A_Valid_3_delay_29_20;
    io_A_Valid_3_delay_31_18 <= io_A_Valid_3_delay_30_19;
    io_A_Valid_3_delay_32_17 <= io_A_Valid_3_delay_31_18;
    io_A_Valid_3_delay_33_16 <= io_A_Valid_3_delay_32_17;
    io_A_Valid_3_delay_34_15 <= io_A_Valid_3_delay_33_16;
    io_A_Valid_3_delay_35_14 <= io_A_Valid_3_delay_34_15;
    io_A_Valid_3_delay_36_13 <= io_A_Valid_3_delay_35_14;
    io_A_Valid_3_delay_37_12 <= io_A_Valid_3_delay_36_13;
    io_A_Valid_3_delay_38_11 <= io_A_Valid_3_delay_37_12;
    io_A_Valid_3_delay_39_10 <= io_A_Valid_3_delay_38_11;
    io_A_Valid_3_delay_40_9 <= io_A_Valid_3_delay_39_10;
    io_A_Valid_3_delay_41_8 <= io_A_Valid_3_delay_40_9;
    io_A_Valid_3_delay_42_7 <= io_A_Valid_3_delay_41_8;
    io_A_Valid_3_delay_43_6 <= io_A_Valid_3_delay_42_7;
    io_A_Valid_3_delay_44_5 <= io_A_Valid_3_delay_43_6;
    io_A_Valid_3_delay_45_4 <= io_A_Valid_3_delay_44_5;
    io_A_Valid_3_delay_46_3 <= io_A_Valid_3_delay_45_4;
    io_A_Valid_3_delay_47_2 <= io_A_Valid_3_delay_46_3;
    io_A_Valid_3_delay_48_1 <= io_A_Valid_3_delay_47_2;
    io_A_Valid_3_delay_49 <= io_A_Valid_3_delay_48_1;
    io_B_Valid_49_delay_1_2 <= io_B_Valid_49;
    io_B_Valid_49_delay_2_1 <= io_B_Valid_49_delay_1_2;
    io_B_Valid_49_delay_3 <= io_B_Valid_49_delay_2_1;
    io_A_Valid_3_delay_1_49 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_48 <= io_A_Valid_3_delay_1_49;
    io_A_Valid_3_delay_3_47 <= io_A_Valid_3_delay_2_48;
    io_A_Valid_3_delay_4_46 <= io_A_Valid_3_delay_3_47;
    io_A_Valid_3_delay_5_45 <= io_A_Valid_3_delay_4_46;
    io_A_Valid_3_delay_6_44 <= io_A_Valid_3_delay_5_45;
    io_A_Valid_3_delay_7_43 <= io_A_Valid_3_delay_6_44;
    io_A_Valid_3_delay_8_42 <= io_A_Valid_3_delay_7_43;
    io_A_Valid_3_delay_9_41 <= io_A_Valid_3_delay_8_42;
    io_A_Valid_3_delay_10_40 <= io_A_Valid_3_delay_9_41;
    io_A_Valid_3_delay_11_39 <= io_A_Valid_3_delay_10_40;
    io_A_Valid_3_delay_12_38 <= io_A_Valid_3_delay_11_39;
    io_A_Valid_3_delay_13_37 <= io_A_Valid_3_delay_12_38;
    io_A_Valid_3_delay_14_36 <= io_A_Valid_3_delay_13_37;
    io_A_Valid_3_delay_15_35 <= io_A_Valid_3_delay_14_36;
    io_A_Valid_3_delay_16_34 <= io_A_Valid_3_delay_15_35;
    io_A_Valid_3_delay_17_33 <= io_A_Valid_3_delay_16_34;
    io_A_Valid_3_delay_18_32 <= io_A_Valid_3_delay_17_33;
    io_A_Valid_3_delay_19_31 <= io_A_Valid_3_delay_18_32;
    io_A_Valid_3_delay_20_30 <= io_A_Valid_3_delay_19_31;
    io_A_Valid_3_delay_21_29 <= io_A_Valid_3_delay_20_30;
    io_A_Valid_3_delay_22_28 <= io_A_Valid_3_delay_21_29;
    io_A_Valid_3_delay_23_27 <= io_A_Valid_3_delay_22_28;
    io_A_Valid_3_delay_24_26 <= io_A_Valid_3_delay_23_27;
    io_A_Valid_3_delay_25_25 <= io_A_Valid_3_delay_24_26;
    io_A_Valid_3_delay_26_24 <= io_A_Valid_3_delay_25_25;
    io_A_Valid_3_delay_27_23 <= io_A_Valid_3_delay_26_24;
    io_A_Valid_3_delay_28_22 <= io_A_Valid_3_delay_27_23;
    io_A_Valid_3_delay_29_21 <= io_A_Valid_3_delay_28_22;
    io_A_Valid_3_delay_30_20 <= io_A_Valid_3_delay_29_21;
    io_A_Valid_3_delay_31_19 <= io_A_Valid_3_delay_30_20;
    io_A_Valid_3_delay_32_18 <= io_A_Valid_3_delay_31_19;
    io_A_Valid_3_delay_33_17 <= io_A_Valid_3_delay_32_18;
    io_A_Valid_3_delay_34_16 <= io_A_Valid_3_delay_33_17;
    io_A_Valid_3_delay_35_15 <= io_A_Valid_3_delay_34_16;
    io_A_Valid_3_delay_36_14 <= io_A_Valid_3_delay_35_15;
    io_A_Valid_3_delay_37_13 <= io_A_Valid_3_delay_36_14;
    io_A_Valid_3_delay_38_12 <= io_A_Valid_3_delay_37_13;
    io_A_Valid_3_delay_39_11 <= io_A_Valid_3_delay_38_12;
    io_A_Valid_3_delay_40_10 <= io_A_Valid_3_delay_39_11;
    io_A_Valid_3_delay_41_9 <= io_A_Valid_3_delay_40_10;
    io_A_Valid_3_delay_42_8 <= io_A_Valid_3_delay_41_9;
    io_A_Valid_3_delay_43_7 <= io_A_Valid_3_delay_42_8;
    io_A_Valid_3_delay_44_6 <= io_A_Valid_3_delay_43_7;
    io_A_Valid_3_delay_45_5 <= io_A_Valid_3_delay_44_6;
    io_A_Valid_3_delay_46_4 <= io_A_Valid_3_delay_45_5;
    io_A_Valid_3_delay_47_3 <= io_A_Valid_3_delay_46_4;
    io_A_Valid_3_delay_48_2 <= io_A_Valid_3_delay_47_3;
    io_A_Valid_3_delay_49_1 <= io_A_Valid_3_delay_48_2;
    io_A_Valid_3_delay_50 <= io_A_Valid_3_delay_49_1;
    io_B_Valid_50_delay_1_2 <= io_B_Valid_50;
    io_B_Valid_50_delay_2_1 <= io_B_Valid_50_delay_1_2;
    io_B_Valid_50_delay_3 <= io_B_Valid_50_delay_2_1;
    io_A_Valid_3_delay_1_50 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_49 <= io_A_Valid_3_delay_1_50;
    io_A_Valid_3_delay_3_48 <= io_A_Valid_3_delay_2_49;
    io_A_Valid_3_delay_4_47 <= io_A_Valid_3_delay_3_48;
    io_A_Valid_3_delay_5_46 <= io_A_Valid_3_delay_4_47;
    io_A_Valid_3_delay_6_45 <= io_A_Valid_3_delay_5_46;
    io_A_Valid_3_delay_7_44 <= io_A_Valid_3_delay_6_45;
    io_A_Valid_3_delay_8_43 <= io_A_Valid_3_delay_7_44;
    io_A_Valid_3_delay_9_42 <= io_A_Valid_3_delay_8_43;
    io_A_Valid_3_delay_10_41 <= io_A_Valid_3_delay_9_42;
    io_A_Valid_3_delay_11_40 <= io_A_Valid_3_delay_10_41;
    io_A_Valid_3_delay_12_39 <= io_A_Valid_3_delay_11_40;
    io_A_Valid_3_delay_13_38 <= io_A_Valid_3_delay_12_39;
    io_A_Valid_3_delay_14_37 <= io_A_Valid_3_delay_13_38;
    io_A_Valid_3_delay_15_36 <= io_A_Valid_3_delay_14_37;
    io_A_Valid_3_delay_16_35 <= io_A_Valid_3_delay_15_36;
    io_A_Valid_3_delay_17_34 <= io_A_Valid_3_delay_16_35;
    io_A_Valid_3_delay_18_33 <= io_A_Valid_3_delay_17_34;
    io_A_Valid_3_delay_19_32 <= io_A_Valid_3_delay_18_33;
    io_A_Valid_3_delay_20_31 <= io_A_Valid_3_delay_19_32;
    io_A_Valid_3_delay_21_30 <= io_A_Valid_3_delay_20_31;
    io_A_Valid_3_delay_22_29 <= io_A_Valid_3_delay_21_30;
    io_A_Valid_3_delay_23_28 <= io_A_Valid_3_delay_22_29;
    io_A_Valid_3_delay_24_27 <= io_A_Valid_3_delay_23_28;
    io_A_Valid_3_delay_25_26 <= io_A_Valid_3_delay_24_27;
    io_A_Valid_3_delay_26_25 <= io_A_Valid_3_delay_25_26;
    io_A_Valid_3_delay_27_24 <= io_A_Valid_3_delay_26_25;
    io_A_Valid_3_delay_28_23 <= io_A_Valid_3_delay_27_24;
    io_A_Valid_3_delay_29_22 <= io_A_Valid_3_delay_28_23;
    io_A_Valid_3_delay_30_21 <= io_A_Valid_3_delay_29_22;
    io_A_Valid_3_delay_31_20 <= io_A_Valid_3_delay_30_21;
    io_A_Valid_3_delay_32_19 <= io_A_Valid_3_delay_31_20;
    io_A_Valid_3_delay_33_18 <= io_A_Valid_3_delay_32_19;
    io_A_Valid_3_delay_34_17 <= io_A_Valid_3_delay_33_18;
    io_A_Valid_3_delay_35_16 <= io_A_Valid_3_delay_34_17;
    io_A_Valid_3_delay_36_15 <= io_A_Valid_3_delay_35_16;
    io_A_Valid_3_delay_37_14 <= io_A_Valid_3_delay_36_15;
    io_A_Valid_3_delay_38_13 <= io_A_Valid_3_delay_37_14;
    io_A_Valid_3_delay_39_12 <= io_A_Valid_3_delay_38_13;
    io_A_Valid_3_delay_40_11 <= io_A_Valid_3_delay_39_12;
    io_A_Valid_3_delay_41_10 <= io_A_Valid_3_delay_40_11;
    io_A_Valid_3_delay_42_9 <= io_A_Valid_3_delay_41_10;
    io_A_Valid_3_delay_43_8 <= io_A_Valid_3_delay_42_9;
    io_A_Valid_3_delay_44_7 <= io_A_Valid_3_delay_43_8;
    io_A_Valid_3_delay_45_6 <= io_A_Valid_3_delay_44_7;
    io_A_Valid_3_delay_46_5 <= io_A_Valid_3_delay_45_6;
    io_A_Valid_3_delay_47_4 <= io_A_Valid_3_delay_46_5;
    io_A_Valid_3_delay_48_3 <= io_A_Valid_3_delay_47_4;
    io_A_Valid_3_delay_49_2 <= io_A_Valid_3_delay_48_3;
    io_A_Valid_3_delay_50_1 <= io_A_Valid_3_delay_49_2;
    io_A_Valid_3_delay_51 <= io_A_Valid_3_delay_50_1;
    io_B_Valid_51_delay_1_2 <= io_B_Valid_51;
    io_B_Valid_51_delay_2_1 <= io_B_Valid_51_delay_1_2;
    io_B_Valid_51_delay_3 <= io_B_Valid_51_delay_2_1;
    io_A_Valid_3_delay_1_51 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_50 <= io_A_Valid_3_delay_1_51;
    io_A_Valid_3_delay_3_49 <= io_A_Valid_3_delay_2_50;
    io_A_Valid_3_delay_4_48 <= io_A_Valid_3_delay_3_49;
    io_A_Valid_3_delay_5_47 <= io_A_Valid_3_delay_4_48;
    io_A_Valid_3_delay_6_46 <= io_A_Valid_3_delay_5_47;
    io_A_Valid_3_delay_7_45 <= io_A_Valid_3_delay_6_46;
    io_A_Valid_3_delay_8_44 <= io_A_Valid_3_delay_7_45;
    io_A_Valid_3_delay_9_43 <= io_A_Valid_3_delay_8_44;
    io_A_Valid_3_delay_10_42 <= io_A_Valid_3_delay_9_43;
    io_A_Valid_3_delay_11_41 <= io_A_Valid_3_delay_10_42;
    io_A_Valid_3_delay_12_40 <= io_A_Valid_3_delay_11_41;
    io_A_Valid_3_delay_13_39 <= io_A_Valid_3_delay_12_40;
    io_A_Valid_3_delay_14_38 <= io_A_Valid_3_delay_13_39;
    io_A_Valid_3_delay_15_37 <= io_A_Valid_3_delay_14_38;
    io_A_Valid_3_delay_16_36 <= io_A_Valid_3_delay_15_37;
    io_A_Valid_3_delay_17_35 <= io_A_Valid_3_delay_16_36;
    io_A_Valid_3_delay_18_34 <= io_A_Valid_3_delay_17_35;
    io_A_Valid_3_delay_19_33 <= io_A_Valid_3_delay_18_34;
    io_A_Valid_3_delay_20_32 <= io_A_Valid_3_delay_19_33;
    io_A_Valid_3_delay_21_31 <= io_A_Valid_3_delay_20_32;
    io_A_Valid_3_delay_22_30 <= io_A_Valid_3_delay_21_31;
    io_A_Valid_3_delay_23_29 <= io_A_Valid_3_delay_22_30;
    io_A_Valid_3_delay_24_28 <= io_A_Valid_3_delay_23_29;
    io_A_Valid_3_delay_25_27 <= io_A_Valid_3_delay_24_28;
    io_A_Valid_3_delay_26_26 <= io_A_Valid_3_delay_25_27;
    io_A_Valid_3_delay_27_25 <= io_A_Valid_3_delay_26_26;
    io_A_Valid_3_delay_28_24 <= io_A_Valid_3_delay_27_25;
    io_A_Valid_3_delay_29_23 <= io_A_Valid_3_delay_28_24;
    io_A_Valid_3_delay_30_22 <= io_A_Valid_3_delay_29_23;
    io_A_Valid_3_delay_31_21 <= io_A_Valid_3_delay_30_22;
    io_A_Valid_3_delay_32_20 <= io_A_Valid_3_delay_31_21;
    io_A_Valid_3_delay_33_19 <= io_A_Valid_3_delay_32_20;
    io_A_Valid_3_delay_34_18 <= io_A_Valid_3_delay_33_19;
    io_A_Valid_3_delay_35_17 <= io_A_Valid_3_delay_34_18;
    io_A_Valid_3_delay_36_16 <= io_A_Valid_3_delay_35_17;
    io_A_Valid_3_delay_37_15 <= io_A_Valid_3_delay_36_16;
    io_A_Valid_3_delay_38_14 <= io_A_Valid_3_delay_37_15;
    io_A_Valid_3_delay_39_13 <= io_A_Valid_3_delay_38_14;
    io_A_Valid_3_delay_40_12 <= io_A_Valid_3_delay_39_13;
    io_A_Valid_3_delay_41_11 <= io_A_Valid_3_delay_40_12;
    io_A_Valid_3_delay_42_10 <= io_A_Valid_3_delay_41_11;
    io_A_Valid_3_delay_43_9 <= io_A_Valid_3_delay_42_10;
    io_A_Valid_3_delay_44_8 <= io_A_Valid_3_delay_43_9;
    io_A_Valid_3_delay_45_7 <= io_A_Valid_3_delay_44_8;
    io_A_Valid_3_delay_46_6 <= io_A_Valid_3_delay_45_7;
    io_A_Valid_3_delay_47_5 <= io_A_Valid_3_delay_46_6;
    io_A_Valid_3_delay_48_4 <= io_A_Valid_3_delay_47_5;
    io_A_Valid_3_delay_49_3 <= io_A_Valid_3_delay_48_4;
    io_A_Valid_3_delay_50_2 <= io_A_Valid_3_delay_49_3;
    io_A_Valid_3_delay_51_1 <= io_A_Valid_3_delay_50_2;
    io_A_Valid_3_delay_52 <= io_A_Valid_3_delay_51_1;
    io_B_Valid_52_delay_1_2 <= io_B_Valid_52;
    io_B_Valid_52_delay_2_1 <= io_B_Valid_52_delay_1_2;
    io_B_Valid_52_delay_3 <= io_B_Valid_52_delay_2_1;
    io_A_Valid_3_delay_1_52 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_51 <= io_A_Valid_3_delay_1_52;
    io_A_Valid_3_delay_3_50 <= io_A_Valid_3_delay_2_51;
    io_A_Valid_3_delay_4_49 <= io_A_Valid_3_delay_3_50;
    io_A_Valid_3_delay_5_48 <= io_A_Valid_3_delay_4_49;
    io_A_Valid_3_delay_6_47 <= io_A_Valid_3_delay_5_48;
    io_A_Valid_3_delay_7_46 <= io_A_Valid_3_delay_6_47;
    io_A_Valid_3_delay_8_45 <= io_A_Valid_3_delay_7_46;
    io_A_Valid_3_delay_9_44 <= io_A_Valid_3_delay_8_45;
    io_A_Valid_3_delay_10_43 <= io_A_Valid_3_delay_9_44;
    io_A_Valid_3_delay_11_42 <= io_A_Valid_3_delay_10_43;
    io_A_Valid_3_delay_12_41 <= io_A_Valid_3_delay_11_42;
    io_A_Valid_3_delay_13_40 <= io_A_Valid_3_delay_12_41;
    io_A_Valid_3_delay_14_39 <= io_A_Valid_3_delay_13_40;
    io_A_Valid_3_delay_15_38 <= io_A_Valid_3_delay_14_39;
    io_A_Valid_3_delay_16_37 <= io_A_Valid_3_delay_15_38;
    io_A_Valid_3_delay_17_36 <= io_A_Valid_3_delay_16_37;
    io_A_Valid_3_delay_18_35 <= io_A_Valid_3_delay_17_36;
    io_A_Valid_3_delay_19_34 <= io_A_Valid_3_delay_18_35;
    io_A_Valid_3_delay_20_33 <= io_A_Valid_3_delay_19_34;
    io_A_Valid_3_delay_21_32 <= io_A_Valid_3_delay_20_33;
    io_A_Valid_3_delay_22_31 <= io_A_Valid_3_delay_21_32;
    io_A_Valid_3_delay_23_30 <= io_A_Valid_3_delay_22_31;
    io_A_Valid_3_delay_24_29 <= io_A_Valid_3_delay_23_30;
    io_A_Valid_3_delay_25_28 <= io_A_Valid_3_delay_24_29;
    io_A_Valid_3_delay_26_27 <= io_A_Valid_3_delay_25_28;
    io_A_Valid_3_delay_27_26 <= io_A_Valid_3_delay_26_27;
    io_A_Valid_3_delay_28_25 <= io_A_Valid_3_delay_27_26;
    io_A_Valid_3_delay_29_24 <= io_A_Valid_3_delay_28_25;
    io_A_Valid_3_delay_30_23 <= io_A_Valid_3_delay_29_24;
    io_A_Valid_3_delay_31_22 <= io_A_Valid_3_delay_30_23;
    io_A_Valid_3_delay_32_21 <= io_A_Valid_3_delay_31_22;
    io_A_Valid_3_delay_33_20 <= io_A_Valid_3_delay_32_21;
    io_A_Valid_3_delay_34_19 <= io_A_Valid_3_delay_33_20;
    io_A_Valid_3_delay_35_18 <= io_A_Valid_3_delay_34_19;
    io_A_Valid_3_delay_36_17 <= io_A_Valid_3_delay_35_18;
    io_A_Valid_3_delay_37_16 <= io_A_Valid_3_delay_36_17;
    io_A_Valid_3_delay_38_15 <= io_A_Valid_3_delay_37_16;
    io_A_Valid_3_delay_39_14 <= io_A_Valid_3_delay_38_15;
    io_A_Valid_3_delay_40_13 <= io_A_Valid_3_delay_39_14;
    io_A_Valid_3_delay_41_12 <= io_A_Valid_3_delay_40_13;
    io_A_Valid_3_delay_42_11 <= io_A_Valid_3_delay_41_12;
    io_A_Valid_3_delay_43_10 <= io_A_Valid_3_delay_42_11;
    io_A_Valid_3_delay_44_9 <= io_A_Valid_3_delay_43_10;
    io_A_Valid_3_delay_45_8 <= io_A_Valid_3_delay_44_9;
    io_A_Valid_3_delay_46_7 <= io_A_Valid_3_delay_45_8;
    io_A_Valid_3_delay_47_6 <= io_A_Valid_3_delay_46_7;
    io_A_Valid_3_delay_48_5 <= io_A_Valid_3_delay_47_6;
    io_A_Valid_3_delay_49_4 <= io_A_Valid_3_delay_48_5;
    io_A_Valid_3_delay_50_3 <= io_A_Valid_3_delay_49_4;
    io_A_Valid_3_delay_51_2 <= io_A_Valid_3_delay_50_3;
    io_A_Valid_3_delay_52_1 <= io_A_Valid_3_delay_51_2;
    io_A_Valid_3_delay_53 <= io_A_Valid_3_delay_52_1;
    io_B_Valid_53_delay_1_2 <= io_B_Valid_53;
    io_B_Valid_53_delay_2_1 <= io_B_Valid_53_delay_1_2;
    io_B_Valid_53_delay_3 <= io_B_Valid_53_delay_2_1;
    io_A_Valid_3_delay_1_53 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_52 <= io_A_Valid_3_delay_1_53;
    io_A_Valid_3_delay_3_51 <= io_A_Valid_3_delay_2_52;
    io_A_Valid_3_delay_4_50 <= io_A_Valid_3_delay_3_51;
    io_A_Valid_3_delay_5_49 <= io_A_Valid_3_delay_4_50;
    io_A_Valid_3_delay_6_48 <= io_A_Valid_3_delay_5_49;
    io_A_Valid_3_delay_7_47 <= io_A_Valid_3_delay_6_48;
    io_A_Valid_3_delay_8_46 <= io_A_Valid_3_delay_7_47;
    io_A_Valid_3_delay_9_45 <= io_A_Valid_3_delay_8_46;
    io_A_Valid_3_delay_10_44 <= io_A_Valid_3_delay_9_45;
    io_A_Valid_3_delay_11_43 <= io_A_Valid_3_delay_10_44;
    io_A_Valid_3_delay_12_42 <= io_A_Valid_3_delay_11_43;
    io_A_Valid_3_delay_13_41 <= io_A_Valid_3_delay_12_42;
    io_A_Valid_3_delay_14_40 <= io_A_Valid_3_delay_13_41;
    io_A_Valid_3_delay_15_39 <= io_A_Valid_3_delay_14_40;
    io_A_Valid_3_delay_16_38 <= io_A_Valid_3_delay_15_39;
    io_A_Valid_3_delay_17_37 <= io_A_Valid_3_delay_16_38;
    io_A_Valid_3_delay_18_36 <= io_A_Valid_3_delay_17_37;
    io_A_Valid_3_delay_19_35 <= io_A_Valid_3_delay_18_36;
    io_A_Valid_3_delay_20_34 <= io_A_Valid_3_delay_19_35;
    io_A_Valid_3_delay_21_33 <= io_A_Valid_3_delay_20_34;
    io_A_Valid_3_delay_22_32 <= io_A_Valid_3_delay_21_33;
    io_A_Valid_3_delay_23_31 <= io_A_Valid_3_delay_22_32;
    io_A_Valid_3_delay_24_30 <= io_A_Valid_3_delay_23_31;
    io_A_Valid_3_delay_25_29 <= io_A_Valid_3_delay_24_30;
    io_A_Valid_3_delay_26_28 <= io_A_Valid_3_delay_25_29;
    io_A_Valid_3_delay_27_27 <= io_A_Valid_3_delay_26_28;
    io_A_Valid_3_delay_28_26 <= io_A_Valid_3_delay_27_27;
    io_A_Valid_3_delay_29_25 <= io_A_Valid_3_delay_28_26;
    io_A_Valid_3_delay_30_24 <= io_A_Valid_3_delay_29_25;
    io_A_Valid_3_delay_31_23 <= io_A_Valid_3_delay_30_24;
    io_A_Valid_3_delay_32_22 <= io_A_Valid_3_delay_31_23;
    io_A_Valid_3_delay_33_21 <= io_A_Valid_3_delay_32_22;
    io_A_Valid_3_delay_34_20 <= io_A_Valid_3_delay_33_21;
    io_A_Valid_3_delay_35_19 <= io_A_Valid_3_delay_34_20;
    io_A_Valid_3_delay_36_18 <= io_A_Valid_3_delay_35_19;
    io_A_Valid_3_delay_37_17 <= io_A_Valid_3_delay_36_18;
    io_A_Valid_3_delay_38_16 <= io_A_Valid_3_delay_37_17;
    io_A_Valid_3_delay_39_15 <= io_A_Valid_3_delay_38_16;
    io_A_Valid_3_delay_40_14 <= io_A_Valid_3_delay_39_15;
    io_A_Valid_3_delay_41_13 <= io_A_Valid_3_delay_40_14;
    io_A_Valid_3_delay_42_12 <= io_A_Valid_3_delay_41_13;
    io_A_Valid_3_delay_43_11 <= io_A_Valid_3_delay_42_12;
    io_A_Valid_3_delay_44_10 <= io_A_Valid_3_delay_43_11;
    io_A_Valid_3_delay_45_9 <= io_A_Valid_3_delay_44_10;
    io_A_Valid_3_delay_46_8 <= io_A_Valid_3_delay_45_9;
    io_A_Valid_3_delay_47_7 <= io_A_Valid_3_delay_46_8;
    io_A_Valid_3_delay_48_6 <= io_A_Valid_3_delay_47_7;
    io_A_Valid_3_delay_49_5 <= io_A_Valid_3_delay_48_6;
    io_A_Valid_3_delay_50_4 <= io_A_Valid_3_delay_49_5;
    io_A_Valid_3_delay_51_3 <= io_A_Valid_3_delay_50_4;
    io_A_Valid_3_delay_52_2 <= io_A_Valid_3_delay_51_3;
    io_A_Valid_3_delay_53_1 <= io_A_Valid_3_delay_52_2;
    io_A_Valid_3_delay_54 <= io_A_Valid_3_delay_53_1;
    io_B_Valid_54_delay_1_2 <= io_B_Valid_54;
    io_B_Valid_54_delay_2_1 <= io_B_Valid_54_delay_1_2;
    io_B_Valid_54_delay_3 <= io_B_Valid_54_delay_2_1;
    io_A_Valid_3_delay_1_54 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_53 <= io_A_Valid_3_delay_1_54;
    io_A_Valid_3_delay_3_52 <= io_A_Valid_3_delay_2_53;
    io_A_Valid_3_delay_4_51 <= io_A_Valid_3_delay_3_52;
    io_A_Valid_3_delay_5_50 <= io_A_Valid_3_delay_4_51;
    io_A_Valid_3_delay_6_49 <= io_A_Valid_3_delay_5_50;
    io_A_Valid_3_delay_7_48 <= io_A_Valid_3_delay_6_49;
    io_A_Valid_3_delay_8_47 <= io_A_Valid_3_delay_7_48;
    io_A_Valid_3_delay_9_46 <= io_A_Valid_3_delay_8_47;
    io_A_Valid_3_delay_10_45 <= io_A_Valid_3_delay_9_46;
    io_A_Valid_3_delay_11_44 <= io_A_Valid_3_delay_10_45;
    io_A_Valid_3_delay_12_43 <= io_A_Valid_3_delay_11_44;
    io_A_Valid_3_delay_13_42 <= io_A_Valid_3_delay_12_43;
    io_A_Valid_3_delay_14_41 <= io_A_Valid_3_delay_13_42;
    io_A_Valid_3_delay_15_40 <= io_A_Valid_3_delay_14_41;
    io_A_Valid_3_delay_16_39 <= io_A_Valid_3_delay_15_40;
    io_A_Valid_3_delay_17_38 <= io_A_Valid_3_delay_16_39;
    io_A_Valid_3_delay_18_37 <= io_A_Valid_3_delay_17_38;
    io_A_Valid_3_delay_19_36 <= io_A_Valid_3_delay_18_37;
    io_A_Valid_3_delay_20_35 <= io_A_Valid_3_delay_19_36;
    io_A_Valid_3_delay_21_34 <= io_A_Valid_3_delay_20_35;
    io_A_Valid_3_delay_22_33 <= io_A_Valid_3_delay_21_34;
    io_A_Valid_3_delay_23_32 <= io_A_Valid_3_delay_22_33;
    io_A_Valid_3_delay_24_31 <= io_A_Valid_3_delay_23_32;
    io_A_Valid_3_delay_25_30 <= io_A_Valid_3_delay_24_31;
    io_A_Valid_3_delay_26_29 <= io_A_Valid_3_delay_25_30;
    io_A_Valid_3_delay_27_28 <= io_A_Valid_3_delay_26_29;
    io_A_Valid_3_delay_28_27 <= io_A_Valid_3_delay_27_28;
    io_A_Valid_3_delay_29_26 <= io_A_Valid_3_delay_28_27;
    io_A_Valid_3_delay_30_25 <= io_A_Valid_3_delay_29_26;
    io_A_Valid_3_delay_31_24 <= io_A_Valid_3_delay_30_25;
    io_A_Valid_3_delay_32_23 <= io_A_Valid_3_delay_31_24;
    io_A_Valid_3_delay_33_22 <= io_A_Valid_3_delay_32_23;
    io_A_Valid_3_delay_34_21 <= io_A_Valid_3_delay_33_22;
    io_A_Valid_3_delay_35_20 <= io_A_Valid_3_delay_34_21;
    io_A_Valid_3_delay_36_19 <= io_A_Valid_3_delay_35_20;
    io_A_Valid_3_delay_37_18 <= io_A_Valid_3_delay_36_19;
    io_A_Valid_3_delay_38_17 <= io_A_Valid_3_delay_37_18;
    io_A_Valid_3_delay_39_16 <= io_A_Valid_3_delay_38_17;
    io_A_Valid_3_delay_40_15 <= io_A_Valid_3_delay_39_16;
    io_A_Valid_3_delay_41_14 <= io_A_Valid_3_delay_40_15;
    io_A_Valid_3_delay_42_13 <= io_A_Valid_3_delay_41_14;
    io_A_Valid_3_delay_43_12 <= io_A_Valid_3_delay_42_13;
    io_A_Valid_3_delay_44_11 <= io_A_Valid_3_delay_43_12;
    io_A_Valid_3_delay_45_10 <= io_A_Valid_3_delay_44_11;
    io_A_Valid_3_delay_46_9 <= io_A_Valid_3_delay_45_10;
    io_A_Valid_3_delay_47_8 <= io_A_Valid_3_delay_46_9;
    io_A_Valid_3_delay_48_7 <= io_A_Valid_3_delay_47_8;
    io_A_Valid_3_delay_49_6 <= io_A_Valid_3_delay_48_7;
    io_A_Valid_3_delay_50_5 <= io_A_Valid_3_delay_49_6;
    io_A_Valid_3_delay_51_4 <= io_A_Valid_3_delay_50_5;
    io_A_Valid_3_delay_52_3 <= io_A_Valid_3_delay_51_4;
    io_A_Valid_3_delay_53_2 <= io_A_Valid_3_delay_52_3;
    io_A_Valid_3_delay_54_1 <= io_A_Valid_3_delay_53_2;
    io_A_Valid_3_delay_55 <= io_A_Valid_3_delay_54_1;
    io_B_Valid_55_delay_1_2 <= io_B_Valid_55;
    io_B_Valid_55_delay_2_1 <= io_B_Valid_55_delay_1_2;
    io_B_Valid_55_delay_3 <= io_B_Valid_55_delay_2_1;
    io_A_Valid_3_delay_1_55 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_54 <= io_A_Valid_3_delay_1_55;
    io_A_Valid_3_delay_3_53 <= io_A_Valid_3_delay_2_54;
    io_A_Valid_3_delay_4_52 <= io_A_Valid_3_delay_3_53;
    io_A_Valid_3_delay_5_51 <= io_A_Valid_3_delay_4_52;
    io_A_Valid_3_delay_6_50 <= io_A_Valid_3_delay_5_51;
    io_A_Valid_3_delay_7_49 <= io_A_Valid_3_delay_6_50;
    io_A_Valid_3_delay_8_48 <= io_A_Valid_3_delay_7_49;
    io_A_Valid_3_delay_9_47 <= io_A_Valid_3_delay_8_48;
    io_A_Valid_3_delay_10_46 <= io_A_Valid_3_delay_9_47;
    io_A_Valid_3_delay_11_45 <= io_A_Valid_3_delay_10_46;
    io_A_Valid_3_delay_12_44 <= io_A_Valid_3_delay_11_45;
    io_A_Valid_3_delay_13_43 <= io_A_Valid_3_delay_12_44;
    io_A_Valid_3_delay_14_42 <= io_A_Valid_3_delay_13_43;
    io_A_Valid_3_delay_15_41 <= io_A_Valid_3_delay_14_42;
    io_A_Valid_3_delay_16_40 <= io_A_Valid_3_delay_15_41;
    io_A_Valid_3_delay_17_39 <= io_A_Valid_3_delay_16_40;
    io_A_Valid_3_delay_18_38 <= io_A_Valid_3_delay_17_39;
    io_A_Valid_3_delay_19_37 <= io_A_Valid_3_delay_18_38;
    io_A_Valid_3_delay_20_36 <= io_A_Valid_3_delay_19_37;
    io_A_Valid_3_delay_21_35 <= io_A_Valid_3_delay_20_36;
    io_A_Valid_3_delay_22_34 <= io_A_Valid_3_delay_21_35;
    io_A_Valid_3_delay_23_33 <= io_A_Valid_3_delay_22_34;
    io_A_Valid_3_delay_24_32 <= io_A_Valid_3_delay_23_33;
    io_A_Valid_3_delay_25_31 <= io_A_Valid_3_delay_24_32;
    io_A_Valid_3_delay_26_30 <= io_A_Valid_3_delay_25_31;
    io_A_Valid_3_delay_27_29 <= io_A_Valid_3_delay_26_30;
    io_A_Valid_3_delay_28_28 <= io_A_Valid_3_delay_27_29;
    io_A_Valid_3_delay_29_27 <= io_A_Valid_3_delay_28_28;
    io_A_Valid_3_delay_30_26 <= io_A_Valid_3_delay_29_27;
    io_A_Valid_3_delay_31_25 <= io_A_Valid_3_delay_30_26;
    io_A_Valid_3_delay_32_24 <= io_A_Valid_3_delay_31_25;
    io_A_Valid_3_delay_33_23 <= io_A_Valid_3_delay_32_24;
    io_A_Valid_3_delay_34_22 <= io_A_Valid_3_delay_33_23;
    io_A_Valid_3_delay_35_21 <= io_A_Valid_3_delay_34_22;
    io_A_Valid_3_delay_36_20 <= io_A_Valid_3_delay_35_21;
    io_A_Valid_3_delay_37_19 <= io_A_Valid_3_delay_36_20;
    io_A_Valid_3_delay_38_18 <= io_A_Valid_3_delay_37_19;
    io_A_Valid_3_delay_39_17 <= io_A_Valid_3_delay_38_18;
    io_A_Valid_3_delay_40_16 <= io_A_Valid_3_delay_39_17;
    io_A_Valid_3_delay_41_15 <= io_A_Valid_3_delay_40_16;
    io_A_Valid_3_delay_42_14 <= io_A_Valid_3_delay_41_15;
    io_A_Valid_3_delay_43_13 <= io_A_Valid_3_delay_42_14;
    io_A_Valid_3_delay_44_12 <= io_A_Valid_3_delay_43_13;
    io_A_Valid_3_delay_45_11 <= io_A_Valid_3_delay_44_12;
    io_A_Valid_3_delay_46_10 <= io_A_Valid_3_delay_45_11;
    io_A_Valid_3_delay_47_9 <= io_A_Valid_3_delay_46_10;
    io_A_Valid_3_delay_48_8 <= io_A_Valid_3_delay_47_9;
    io_A_Valid_3_delay_49_7 <= io_A_Valid_3_delay_48_8;
    io_A_Valid_3_delay_50_6 <= io_A_Valid_3_delay_49_7;
    io_A_Valid_3_delay_51_5 <= io_A_Valid_3_delay_50_6;
    io_A_Valid_3_delay_52_4 <= io_A_Valid_3_delay_51_5;
    io_A_Valid_3_delay_53_3 <= io_A_Valid_3_delay_52_4;
    io_A_Valid_3_delay_54_2 <= io_A_Valid_3_delay_53_3;
    io_A_Valid_3_delay_55_1 <= io_A_Valid_3_delay_54_2;
    io_A_Valid_3_delay_56 <= io_A_Valid_3_delay_55_1;
    io_B_Valid_56_delay_1_2 <= io_B_Valid_56;
    io_B_Valid_56_delay_2_1 <= io_B_Valid_56_delay_1_2;
    io_B_Valid_56_delay_3 <= io_B_Valid_56_delay_2_1;
    io_A_Valid_3_delay_1_56 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_55 <= io_A_Valid_3_delay_1_56;
    io_A_Valid_3_delay_3_54 <= io_A_Valid_3_delay_2_55;
    io_A_Valid_3_delay_4_53 <= io_A_Valid_3_delay_3_54;
    io_A_Valid_3_delay_5_52 <= io_A_Valid_3_delay_4_53;
    io_A_Valid_3_delay_6_51 <= io_A_Valid_3_delay_5_52;
    io_A_Valid_3_delay_7_50 <= io_A_Valid_3_delay_6_51;
    io_A_Valid_3_delay_8_49 <= io_A_Valid_3_delay_7_50;
    io_A_Valid_3_delay_9_48 <= io_A_Valid_3_delay_8_49;
    io_A_Valid_3_delay_10_47 <= io_A_Valid_3_delay_9_48;
    io_A_Valid_3_delay_11_46 <= io_A_Valid_3_delay_10_47;
    io_A_Valid_3_delay_12_45 <= io_A_Valid_3_delay_11_46;
    io_A_Valid_3_delay_13_44 <= io_A_Valid_3_delay_12_45;
    io_A_Valid_3_delay_14_43 <= io_A_Valid_3_delay_13_44;
    io_A_Valid_3_delay_15_42 <= io_A_Valid_3_delay_14_43;
    io_A_Valid_3_delay_16_41 <= io_A_Valid_3_delay_15_42;
    io_A_Valid_3_delay_17_40 <= io_A_Valid_3_delay_16_41;
    io_A_Valid_3_delay_18_39 <= io_A_Valid_3_delay_17_40;
    io_A_Valid_3_delay_19_38 <= io_A_Valid_3_delay_18_39;
    io_A_Valid_3_delay_20_37 <= io_A_Valid_3_delay_19_38;
    io_A_Valid_3_delay_21_36 <= io_A_Valid_3_delay_20_37;
    io_A_Valid_3_delay_22_35 <= io_A_Valid_3_delay_21_36;
    io_A_Valid_3_delay_23_34 <= io_A_Valid_3_delay_22_35;
    io_A_Valid_3_delay_24_33 <= io_A_Valid_3_delay_23_34;
    io_A_Valid_3_delay_25_32 <= io_A_Valid_3_delay_24_33;
    io_A_Valid_3_delay_26_31 <= io_A_Valid_3_delay_25_32;
    io_A_Valid_3_delay_27_30 <= io_A_Valid_3_delay_26_31;
    io_A_Valid_3_delay_28_29 <= io_A_Valid_3_delay_27_30;
    io_A_Valid_3_delay_29_28 <= io_A_Valid_3_delay_28_29;
    io_A_Valid_3_delay_30_27 <= io_A_Valid_3_delay_29_28;
    io_A_Valid_3_delay_31_26 <= io_A_Valid_3_delay_30_27;
    io_A_Valid_3_delay_32_25 <= io_A_Valid_3_delay_31_26;
    io_A_Valid_3_delay_33_24 <= io_A_Valid_3_delay_32_25;
    io_A_Valid_3_delay_34_23 <= io_A_Valid_3_delay_33_24;
    io_A_Valid_3_delay_35_22 <= io_A_Valid_3_delay_34_23;
    io_A_Valid_3_delay_36_21 <= io_A_Valid_3_delay_35_22;
    io_A_Valid_3_delay_37_20 <= io_A_Valid_3_delay_36_21;
    io_A_Valid_3_delay_38_19 <= io_A_Valid_3_delay_37_20;
    io_A_Valid_3_delay_39_18 <= io_A_Valid_3_delay_38_19;
    io_A_Valid_3_delay_40_17 <= io_A_Valid_3_delay_39_18;
    io_A_Valid_3_delay_41_16 <= io_A_Valid_3_delay_40_17;
    io_A_Valid_3_delay_42_15 <= io_A_Valid_3_delay_41_16;
    io_A_Valid_3_delay_43_14 <= io_A_Valid_3_delay_42_15;
    io_A_Valid_3_delay_44_13 <= io_A_Valid_3_delay_43_14;
    io_A_Valid_3_delay_45_12 <= io_A_Valid_3_delay_44_13;
    io_A_Valid_3_delay_46_11 <= io_A_Valid_3_delay_45_12;
    io_A_Valid_3_delay_47_10 <= io_A_Valid_3_delay_46_11;
    io_A_Valid_3_delay_48_9 <= io_A_Valid_3_delay_47_10;
    io_A_Valid_3_delay_49_8 <= io_A_Valid_3_delay_48_9;
    io_A_Valid_3_delay_50_7 <= io_A_Valid_3_delay_49_8;
    io_A_Valid_3_delay_51_6 <= io_A_Valid_3_delay_50_7;
    io_A_Valid_3_delay_52_5 <= io_A_Valid_3_delay_51_6;
    io_A_Valid_3_delay_53_4 <= io_A_Valid_3_delay_52_5;
    io_A_Valid_3_delay_54_3 <= io_A_Valid_3_delay_53_4;
    io_A_Valid_3_delay_55_2 <= io_A_Valid_3_delay_54_3;
    io_A_Valid_3_delay_56_1 <= io_A_Valid_3_delay_55_2;
    io_A_Valid_3_delay_57 <= io_A_Valid_3_delay_56_1;
    io_B_Valid_57_delay_1_2 <= io_B_Valid_57;
    io_B_Valid_57_delay_2_1 <= io_B_Valid_57_delay_1_2;
    io_B_Valid_57_delay_3 <= io_B_Valid_57_delay_2_1;
    io_A_Valid_3_delay_1_57 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_56 <= io_A_Valid_3_delay_1_57;
    io_A_Valid_3_delay_3_55 <= io_A_Valid_3_delay_2_56;
    io_A_Valid_3_delay_4_54 <= io_A_Valid_3_delay_3_55;
    io_A_Valid_3_delay_5_53 <= io_A_Valid_3_delay_4_54;
    io_A_Valid_3_delay_6_52 <= io_A_Valid_3_delay_5_53;
    io_A_Valid_3_delay_7_51 <= io_A_Valid_3_delay_6_52;
    io_A_Valid_3_delay_8_50 <= io_A_Valid_3_delay_7_51;
    io_A_Valid_3_delay_9_49 <= io_A_Valid_3_delay_8_50;
    io_A_Valid_3_delay_10_48 <= io_A_Valid_3_delay_9_49;
    io_A_Valid_3_delay_11_47 <= io_A_Valid_3_delay_10_48;
    io_A_Valid_3_delay_12_46 <= io_A_Valid_3_delay_11_47;
    io_A_Valid_3_delay_13_45 <= io_A_Valid_3_delay_12_46;
    io_A_Valid_3_delay_14_44 <= io_A_Valid_3_delay_13_45;
    io_A_Valid_3_delay_15_43 <= io_A_Valid_3_delay_14_44;
    io_A_Valid_3_delay_16_42 <= io_A_Valid_3_delay_15_43;
    io_A_Valid_3_delay_17_41 <= io_A_Valid_3_delay_16_42;
    io_A_Valid_3_delay_18_40 <= io_A_Valid_3_delay_17_41;
    io_A_Valid_3_delay_19_39 <= io_A_Valid_3_delay_18_40;
    io_A_Valid_3_delay_20_38 <= io_A_Valid_3_delay_19_39;
    io_A_Valid_3_delay_21_37 <= io_A_Valid_3_delay_20_38;
    io_A_Valid_3_delay_22_36 <= io_A_Valid_3_delay_21_37;
    io_A_Valid_3_delay_23_35 <= io_A_Valid_3_delay_22_36;
    io_A_Valid_3_delay_24_34 <= io_A_Valid_3_delay_23_35;
    io_A_Valid_3_delay_25_33 <= io_A_Valid_3_delay_24_34;
    io_A_Valid_3_delay_26_32 <= io_A_Valid_3_delay_25_33;
    io_A_Valid_3_delay_27_31 <= io_A_Valid_3_delay_26_32;
    io_A_Valid_3_delay_28_30 <= io_A_Valid_3_delay_27_31;
    io_A_Valid_3_delay_29_29 <= io_A_Valid_3_delay_28_30;
    io_A_Valid_3_delay_30_28 <= io_A_Valid_3_delay_29_29;
    io_A_Valid_3_delay_31_27 <= io_A_Valid_3_delay_30_28;
    io_A_Valid_3_delay_32_26 <= io_A_Valid_3_delay_31_27;
    io_A_Valid_3_delay_33_25 <= io_A_Valid_3_delay_32_26;
    io_A_Valid_3_delay_34_24 <= io_A_Valid_3_delay_33_25;
    io_A_Valid_3_delay_35_23 <= io_A_Valid_3_delay_34_24;
    io_A_Valid_3_delay_36_22 <= io_A_Valid_3_delay_35_23;
    io_A_Valid_3_delay_37_21 <= io_A_Valid_3_delay_36_22;
    io_A_Valid_3_delay_38_20 <= io_A_Valid_3_delay_37_21;
    io_A_Valid_3_delay_39_19 <= io_A_Valid_3_delay_38_20;
    io_A_Valid_3_delay_40_18 <= io_A_Valid_3_delay_39_19;
    io_A_Valid_3_delay_41_17 <= io_A_Valid_3_delay_40_18;
    io_A_Valid_3_delay_42_16 <= io_A_Valid_3_delay_41_17;
    io_A_Valid_3_delay_43_15 <= io_A_Valid_3_delay_42_16;
    io_A_Valid_3_delay_44_14 <= io_A_Valid_3_delay_43_15;
    io_A_Valid_3_delay_45_13 <= io_A_Valid_3_delay_44_14;
    io_A_Valid_3_delay_46_12 <= io_A_Valid_3_delay_45_13;
    io_A_Valid_3_delay_47_11 <= io_A_Valid_3_delay_46_12;
    io_A_Valid_3_delay_48_10 <= io_A_Valid_3_delay_47_11;
    io_A_Valid_3_delay_49_9 <= io_A_Valid_3_delay_48_10;
    io_A_Valid_3_delay_50_8 <= io_A_Valid_3_delay_49_9;
    io_A_Valid_3_delay_51_7 <= io_A_Valid_3_delay_50_8;
    io_A_Valid_3_delay_52_6 <= io_A_Valid_3_delay_51_7;
    io_A_Valid_3_delay_53_5 <= io_A_Valid_3_delay_52_6;
    io_A_Valid_3_delay_54_4 <= io_A_Valid_3_delay_53_5;
    io_A_Valid_3_delay_55_3 <= io_A_Valid_3_delay_54_4;
    io_A_Valid_3_delay_56_2 <= io_A_Valid_3_delay_55_3;
    io_A_Valid_3_delay_57_1 <= io_A_Valid_3_delay_56_2;
    io_A_Valid_3_delay_58 <= io_A_Valid_3_delay_57_1;
    io_B_Valid_58_delay_1_2 <= io_B_Valid_58;
    io_B_Valid_58_delay_2_1 <= io_B_Valid_58_delay_1_2;
    io_B_Valid_58_delay_3 <= io_B_Valid_58_delay_2_1;
    io_A_Valid_3_delay_1_58 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_57 <= io_A_Valid_3_delay_1_58;
    io_A_Valid_3_delay_3_56 <= io_A_Valid_3_delay_2_57;
    io_A_Valid_3_delay_4_55 <= io_A_Valid_3_delay_3_56;
    io_A_Valid_3_delay_5_54 <= io_A_Valid_3_delay_4_55;
    io_A_Valid_3_delay_6_53 <= io_A_Valid_3_delay_5_54;
    io_A_Valid_3_delay_7_52 <= io_A_Valid_3_delay_6_53;
    io_A_Valid_3_delay_8_51 <= io_A_Valid_3_delay_7_52;
    io_A_Valid_3_delay_9_50 <= io_A_Valid_3_delay_8_51;
    io_A_Valid_3_delay_10_49 <= io_A_Valid_3_delay_9_50;
    io_A_Valid_3_delay_11_48 <= io_A_Valid_3_delay_10_49;
    io_A_Valid_3_delay_12_47 <= io_A_Valid_3_delay_11_48;
    io_A_Valid_3_delay_13_46 <= io_A_Valid_3_delay_12_47;
    io_A_Valid_3_delay_14_45 <= io_A_Valid_3_delay_13_46;
    io_A_Valid_3_delay_15_44 <= io_A_Valid_3_delay_14_45;
    io_A_Valid_3_delay_16_43 <= io_A_Valid_3_delay_15_44;
    io_A_Valid_3_delay_17_42 <= io_A_Valid_3_delay_16_43;
    io_A_Valid_3_delay_18_41 <= io_A_Valid_3_delay_17_42;
    io_A_Valid_3_delay_19_40 <= io_A_Valid_3_delay_18_41;
    io_A_Valid_3_delay_20_39 <= io_A_Valid_3_delay_19_40;
    io_A_Valid_3_delay_21_38 <= io_A_Valid_3_delay_20_39;
    io_A_Valid_3_delay_22_37 <= io_A_Valid_3_delay_21_38;
    io_A_Valid_3_delay_23_36 <= io_A_Valid_3_delay_22_37;
    io_A_Valid_3_delay_24_35 <= io_A_Valid_3_delay_23_36;
    io_A_Valid_3_delay_25_34 <= io_A_Valid_3_delay_24_35;
    io_A_Valid_3_delay_26_33 <= io_A_Valid_3_delay_25_34;
    io_A_Valid_3_delay_27_32 <= io_A_Valid_3_delay_26_33;
    io_A_Valid_3_delay_28_31 <= io_A_Valid_3_delay_27_32;
    io_A_Valid_3_delay_29_30 <= io_A_Valid_3_delay_28_31;
    io_A_Valid_3_delay_30_29 <= io_A_Valid_3_delay_29_30;
    io_A_Valid_3_delay_31_28 <= io_A_Valid_3_delay_30_29;
    io_A_Valid_3_delay_32_27 <= io_A_Valid_3_delay_31_28;
    io_A_Valid_3_delay_33_26 <= io_A_Valid_3_delay_32_27;
    io_A_Valid_3_delay_34_25 <= io_A_Valid_3_delay_33_26;
    io_A_Valid_3_delay_35_24 <= io_A_Valid_3_delay_34_25;
    io_A_Valid_3_delay_36_23 <= io_A_Valid_3_delay_35_24;
    io_A_Valid_3_delay_37_22 <= io_A_Valid_3_delay_36_23;
    io_A_Valid_3_delay_38_21 <= io_A_Valid_3_delay_37_22;
    io_A_Valid_3_delay_39_20 <= io_A_Valid_3_delay_38_21;
    io_A_Valid_3_delay_40_19 <= io_A_Valid_3_delay_39_20;
    io_A_Valid_3_delay_41_18 <= io_A_Valid_3_delay_40_19;
    io_A_Valid_3_delay_42_17 <= io_A_Valid_3_delay_41_18;
    io_A_Valid_3_delay_43_16 <= io_A_Valid_3_delay_42_17;
    io_A_Valid_3_delay_44_15 <= io_A_Valid_3_delay_43_16;
    io_A_Valid_3_delay_45_14 <= io_A_Valid_3_delay_44_15;
    io_A_Valid_3_delay_46_13 <= io_A_Valid_3_delay_45_14;
    io_A_Valid_3_delay_47_12 <= io_A_Valid_3_delay_46_13;
    io_A_Valid_3_delay_48_11 <= io_A_Valid_3_delay_47_12;
    io_A_Valid_3_delay_49_10 <= io_A_Valid_3_delay_48_11;
    io_A_Valid_3_delay_50_9 <= io_A_Valid_3_delay_49_10;
    io_A_Valid_3_delay_51_8 <= io_A_Valid_3_delay_50_9;
    io_A_Valid_3_delay_52_7 <= io_A_Valid_3_delay_51_8;
    io_A_Valid_3_delay_53_6 <= io_A_Valid_3_delay_52_7;
    io_A_Valid_3_delay_54_5 <= io_A_Valid_3_delay_53_6;
    io_A_Valid_3_delay_55_4 <= io_A_Valid_3_delay_54_5;
    io_A_Valid_3_delay_56_3 <= io_A_Valid_3_delay_55_4;
    io_A_Valid_3_delay_57_2 <= io_A_Valid_3_delay_56_3;
    io_A_Valid_3_delay_58_1 <= io_A_Valid_3_delay_57_2;
    io_A_Valid_3_delay_59 <= io_A_Valid_3_delay_58_1;
    io_B_Valid_59_delay_1_2 <= io_B_Valid_59;
    io_B_Valid_59_delay_2_1 <= io_B_Valid_59_delay_1_2;
    io_B_Valid_59_delay_3 <= io_B_Valid_59_delay_2_1;
    io_A_Valid_3_delay_1_59 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_58 <= io_A_Valid_3_delay_1_59;
    io_A_Valid_3_delay_3_57 <= io_A_Valid_3_delay_2_58;
    io_A_Valid_3_delay_4_56 <= io_A_Valid_3_delay_3_57;
    io_A_Valid_3_delay_5_55 <= io_A_Valid_3_delay_4_56;
    io_A_Valid_3_delay_6_54 <= io_A_Valid_3_delay_5_55;
    io_A_Valid_3_delay_7_53 <= io_A_Valid_3_delay_6_54;
    io_A_Valid_3_delay_8_52 <= io_A_Valid_3_delay_7_53;
    io_A_Valid_3_delay_9_51 <= io_A_Valid_3_delay_8_52;
    io_A_Valid_3_delay_10_50 <= io_A_Valid_3_delay_9_51;
    io_A_Valid_3_delay_11_49 <= io_A_Valid_3_delay_10_50;
    io_A_Valid_3_delay_12_48 <= io_A_Valid_3_delay_11_49;
    io_A_Valid_3_delay_13_47 <= io_A_Valid_3_delay_12_48;
    io_A_Valid_3_delay_14_46 <= io_A_Valid_3_delay_13_47;
    io_A_Valid_3_delay_15_45 <= io_A_Valid_3_delay_14_46;
    io_A_Valid_3_delay_16_44 <= io_A_Valid_3_delay_15_45;
    io_A_Valid_3_delay_17_43 <= io_A_Valid_3_delay_16_44;
    io_A_Valid_3_delay_18_42 <= io_A_Valid_3_delay_17_43;
    io_A_Valid_3_delay_19_41 <= io_A_Valid_3_delay_18_42;
    io_A_Valid_3_delay_20_40 <= io_A_Valid_3_delay_19_41;
    io_A_Valid_3_delay_21_39 <= io_A_Valid_3_delay_20_40;
    io_A_Valid_3_delay_22_38 <= io_A_Valid_3_delay_21_39;
    io_A_Valid_3_delay_23_37 <= io_A_Valid_3_delay_22_38;
    io_A_Valid_3_delay_24_36 <= io_A_Valid_3_delay_23_37;
    io_A_Valid_3_delay_25_35 <= io_A_Valid_3_delay_24_36;
    io_A_Valid_3_delay_26_34 <= io_A_Valid_3_delay_25_35;
    io_A_Valid_3_delay_27_33 <= io_A_Valid_3_delay_26_34;
    io_A_Valid_3_delay_28_32 <= io_A_Valid_3_delay_27_33;
    io_A_Valid_3_delay_29_31 <= io_A_Valid_3_delay_28_32;
    io_A_Valid_3_delay_30_30 <= io_A_Valid_3_delay_29_31;
    io_A_Valid_3_delay_31_29 <= io_A_Valid_3_delay_30_30;
    io_A_Valid_3_delay_32_28 <= io_A_Valid_3_delay_31_29;
    io_A_Valid_3_delay_33_27 <= io_A_Valid_3_delay_32_28;
    io_A_Valid_3_delay_34_26 <= io_A_Valid_3_delay_33_27;
    io_A_Valid_3_delay_35_25 <= io_A_Valid_3_delay_34_26;
    io_A_Valid_3_delay_36_24 <= io_A_Valid_3_delay_35_25;
    io_A_Valid_3_delay_37_23 <= io_A_Valid_3_delay_36_24;
    io_A_Valid_3_delay_38_22 <= io_A_Valid_3_delay_37_23;
    io_A_Valid_3_delay_39_21 <= io_A_Valid_3_delay_38_22;
    io_A_Valid_3_delay_40_20 <= io_A_Valid_3_delay_39_21;
    io_A_Valid_3_delay_41_19 <= io_A_Valid_3_delay_40_20;
    io_A_Valid_3_delay_42_18 <= io_A_Valid_3_delay_41_19;
    io_A_Valid_3_delay_43_17 <= io_A_Valid_3_delay_42_18;
    io_A_Valid_3_delay_44_16 <= io_A_Valid_3_delay_43_17;
    io_A_Valid_3_delay_45_15 <= io_A_Valid_3_delay_44_16;
    io_A_Valid_3_delay_46_14 <= io_A_Valid_3_delay_45_15;
    io_A_Valid_3_delay_47_13 <= io_A_Valid_3_delay_46_14;
    io_A_Valid_3_delay_48_12 <= io_A_Valid_3_delay_47_13;
    io_A_Valid_3_delay_49_11 <= io_A_Valid_3_delay_48_12;
    io_A_Valid_3_delay_50_10 <= io_A_Valid_3_delay_49_11;
    io_A_Valid_3_delay_51_9 <= io_A_Valid_3_delay_50_10;
    io_A_Valid_3_delay_52_8 <= io_A_Valid_3_delay_51_9;
    io_A_Valid_3_delay_53_7 <= io_A_Valid_3_delay_52_8;
    io_A_Valid_3_delay_54_6 <= io_A_Valid_3_delay_53_7;
    io_A_Valid_3_delay_55_5 <= io_A_Valid_3_delay_54_6;
    io_A_Valid_3_delay_56_4 <= io_A_Valid_3_delay_55_5;
    io_A_Valid_3_delay_57_3 <= io_A_Valid_3_delay_56_4;
    io_A_Valid_3_delay_58_2 <= io_A_Valid_3_delay_57_3;
    io_A_Valid_3_delay_59_1 <= io_A_Valid_3_delay_58_2;
    io_A_Valid_3_delay_60 <= io_A_Valid_3_delay_59_1;
    io_B_Valid_60_delay_1_2 <= io_B_Valid_60;
    io_B_Valid_60_delay_2_1 <= io_B_Valid_60_delay_1_2;
    io_B_Valid_60_delay_3 <= io_B_Valid_60_delay_2_1;
    io_A_Valid_3_delay_1_60 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_59 <= io_A_Valid_3_delay_1_60;
    io_A_Valid_3_delay_3_58 <= io_A_Valid_3_delay_2_59;
    io_A_Valid_3_delay_4_57 <= io_A_Valid_3_delay_3_58;
    io_A_Valid_3_delay_5_56 <= io_A_Valid_3_delay_4_57;
    io_A_Valid_3_delay_6_55 <= io_A_Valid_3_delay_5_56;
    io_A_Valid_3_delay_7_54 <= io_A_Valid_3_delay_6_55;
    io_A_Valid_3_delay_8_53 <= io_A_Valid_3_delay_7_54;
    io_A_Valid_3_delay_9_52 <= io_A_Valid_3_delay_8_53;
    io_A_Valid_3_delay_10_51 <= io_A_Valid_3_delay_9_52;
    io_A_Valid_3_delay_11_50 <= io_A_Valid_3_delay_10_51;
    io_A_Valid_3_delay_12_49 <= io_A_Valid_3_delay_11_50;
    io_A_Valid_3_delay_13_48 <= io_A_Valid_3_delay_12_49;
    io_A_Valid_3_delay_14_47 <= io_A_Valid_3_delay_13_48;
    io_A_Valid_3_delay_15_46 <= io_A_Valid_3_delay_14_47;
    io_A_Valid_3_delay_16_45 <= io_A_Valid_3_delay_15_46;
    io_A_Valid_3_delay_17_44 <= io_A_Valid_3_delay_16_45;
    io_A_Valid_3_delay_18_43 <= io_A_Valid_3_delay_17_44;
    io_A_Valid_3_delay_19_42 <= io_A_Valid_3_delay_18_43;
    io_A_Valid_3_delay_20_41 <= io_A_Valid_3_delay_19_42;
    io_A_Valid_3_delay_21_40 <= io_A_Valid_3_delay_20_41;
    io_A_Valid_3_delay_22_39 <= io_A_Valid_3_delay_21_40;
    io_A_Valid_3_delay_23_38 <= io_A_Valid_3_delay_22_39;
    io_A_Valid_3_delay_24_37 <= io_A_Valid_3_delay_23_38;
    io_A_Valid_3_delay_25_36 <= io_A_Valid_3_delay_24_37;
    io_A_Valid_3_delay_26_35 <= io_A_Valid_3_delay_25_36;
    io_A_Valid_3_delay_27_34 <= io_A_Valid_3_delay_26_35;
    io_A_Valid_3_delay_28_33 <= io_A_Valid_3_delay_27_34;
    io_A_Valid_3_delay_29_32 <= io_A_Valid_3_delay_28_33;
    io_A_Valid_3_delay_30_31 <= io_A_Valid_3_delay_29_32;
    io_A_Valid_3_delay_31_30 <= io_A_Valid_3_delay_30_31;
    io_A_Valid_3_delay_32_29 <= io_A_Valid_3_delay_31_30;
    io_A_Valid_3_delay_33_28 <= io_A_Valid_3_delay_32_29;
    io_A_Valid_3_delay_34_27 <= io_A_Valid_3_delay_33_28;
    io_A_Valid_3_delay_35_26 <= io_A_Valid_3_delay_34_27;
    io_A_Valid_3_delay_36_25 <= io_A_Valid_3_delay_35_26;
    io_A_Valid_3_delay_37_24 <= io_A_Valid_3_delay_36_25;
    io_A_Valid_3_delay_38_23 <= io_A_Valid_3_delay_37_24;
    io_A_Valid_3_delay_39_22 <= io_A_Valid_3_delay_38_23;
    io_A_Valid_3_delay_40_21 <= io_A_Valid_3_delay_39_22;
    io_A_Valid_3_delay_41_20 <= io_A_Valid_3_delay_40_21;
    io_A_Valid_3_delay_42_19 <= io_A_Valid_3_delay_41_20;
    io_A_Valid_3_delay_43_18 <= io_A_Valid_3_delay_42_19;
    io_A_Valid_3_delay_44_17 <= io_A_Valid_3_delay_43_18;
    io_A_Valid_3_delay_45_16 <= io_A_Valid_3_delay_44_17;
    io_A_Valid_3_delay_46_15 <= io_A_Valid_3_delay_45_16;
    io_A_Valid_3_delay_47_14 <= io_A_Valid_3_delay_46_15;
    io_A_Valid_3_delay_48_13 <= io_A_Valid_3_delay_47_14;
    io_A_Valid_3_delay_49_12 <= io_A_Valid_3_delay_48_13;
    io_A_Valid_3_delay_50_11 <= io_A_Valid_3_delay_49_12;
    io_A_Valid_3_delay_51_10 <= io_A_Valid_3_delay_50_11;
    io_A_Valid_3_delay_52_9 <= io_A_Valid_3_delay_51_10;
    io_A_Valid_3_delay_53_8 <= io_A_Valid_3_delay_52_9;
    io_A_Valid_3_delay_54_7 <= io_A_Valid_3_delay_53_8;
    io_A_Valid_3_delay_55_6 <= io_A_Valid_3_delay_54_7;
    io_A_Valid_3_delay_56_5 <= io_A_Valid_3_delay_55_6;
    io_A_Valid_3_delay_57_4 <= io_A_Valid_3_delay_56_5;
    io_A_Valid_3_delay_58_3 <= io_A_Valid_3_delay_57_4;
    io_A_Valid_3_delay_59_2 <= io_A_Valid_3_delay_58_3;
    io_A_Valid_3_delay_60_1 <= io_A_Valid_3_delay_59_2;
    io_A_Valid_3_delay_61 <= io_A_Valid_3_delay_60_1;
    io_B_Valid_61_delay_1_2 <= io_B_Valid_61;
    io_B_Valid_61_delay_2_1 <= io_B_Valid_61_delay_1_2;
    io_B_Valid_61_delay_3 <= io_B_Valid_61_delay_2_1;
    io_A_Valid_3_delay_1_61 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_60 <= io_A_Valid_3_delay_1_61;
    io_A_Valid_3_delay_3_59 <= io_A_Valid_3_delay_2_60;
    io_A_Valid_3_delay_4_58 <= io_A_Valid_3_delay_3_59;
    io_A_Valid_3_delay_5_57 <= io_A_Valid_3_delay_4_58;
    io_A_Valid_3_delay_6_56 <= io_A_Valid_3_delay_5_57;
    io_A_Valid_3_delay_7_55 <= io_A_Valid_3_delay_6_56;
    io_A_Valid_3_delay_8_54 <= io_A_Valid_3_delay_7_55;
    io_A_Valid_3_delay_9_53 <= io_A_Valid_3_delay_8_54;
    io_A_Valid_3_delay_10_52 <= io_A_Valid_3_delay_9_53;
    io_A_Valid_3_delay_11_51 <= io_A_Valid_3_delay_10_52;
    io_A_Valid_3_delay_12_50 <= io_A_Valid_3_delay_11_51;
    io_A_Valid_3_delay_13_49 <= io_A_Valid_3_delay_12_50;
    io_A_Valid_3_delay_14_48 <= io_A_Valid_3_delay_13_49;
    io_A_Valid_3_delay_15_47 <= io_A_Valid_3_delay_14_48;
    io_A_Valid_3_delay_16_46 <= io_A_Valid_3_delay_15_47;
    io_A_Valid_3_delay_17_45 <= io_A_Valid_3_delay_16_46;
    io_A_Valid_3_delay_18_44 <= io_A_Valid_3_delay_17_45;
    io_A_Valid_3_delay_19_43 <= io_A_Valid_3_delay_18_44;
    io_A_Valid_3_delay_20_42 <= io_A_Valid_3_delay_19_43;
    io_A_Valid_3_delay_21_41 <= io_A_Valid_3_delay_20_42;
    io_A_Valid_3_delay_22_40 <= io_A_Valid_3_delay_21_41;
    io_A_Valid_3_delay_23_39 <= io_A_Valid_3_delay_22_40;
    io_A_Valid_3_delay_24_38 <= io_A_Valid_3_delay_23_39;
    io_A_Valid_3_delay_25_37 <= io_A_Valid_3_delay_24_38;
    io_A_Valid_3_delay_26_36 <= io_A_Valid_3_delay_25_37;
    io_A_Valid_3_delay_27_35 <= io_A_Valid_3_delay_26_36;
    io_A_Valid_3_delay_28_34 <= io_A_Valid_3_delay_27_35;
    io_A_Valid_3_delay_29_33 <= io_A_Valid_3_delay_28_34;
    io_A_Valid_3_delay_30_32 <= io_A_Valid_3_delay_29_33;
    io_A_Valid_3_delay_31_31 <= io_A_Valid_3_delay_30_32;
    io_A_Valid_3_delay_32_30 <= io_A_Valid_3_delay_31_31;
    io_A_Valid_3_delay_33_29 <= io_A_Valid_3_delay_32_30;
    io_A_Valid_3_delay_34_28 <= io_A_Valid_3_delay_33_29;
    io_A_Valid_3_delay_35_27 <= io_A_Valid_3_delay_34_28;
    io_A_Valid_3_delay_36_26 <= io_A_Valid_3_delay_35_27;
    io_A_Valid_3_delay_37_25 <= io_A_Valid_3_delay_36_26;
    io_A_Valid_3_delay_38_24 <= io_A_Valid_3_delay_37_25;
    io_A_Valid_3_delay_39_23 <= io_A_Valid_3_delay_38_24;
    io_A_Valid_3_delay_40_22 <= io_A_Valid_3_delay_39_23;
    io_A_Valid_3_delay_41_21 <= io_A_Valid_3_delay_40_22;
    io_A_Valid_3_delay_42_20 <= io_A_Valid_3_delay_41_21;
    io_A_Valid_3_delay_43_19 <= io_A_Valid_3_delay_42_20;
    io_A_Valid_3_delay_44_18 <= io_A_Valid_3_delay_43_19;
    io_A_Valid_3_delay_45_17 <= io_A_Valid_3_delay_44_18;
    io_A_Valid_3_delay_46_16 <= io_A_Valid_3_delay_45_17;
    io_A_Valid_3_delay_47_15 <= io_A_Valid_3_delay_46_16;
    io_A_Valid_3_delay_48_14 <= io_A_Valid_3_delay_47_15;
    io_A_Valid_3_delay_49_13 <= io_A_Valid_3_delay_48_14;
    io_A_Valid_3_delay_50_12 <= io_A_Valid_3_delay_49_13;
    io_A_Valid_3_delay_51_11 <= io_A_Valid_3_delay_50_12;
    io_A_Valid_3_delay_52_10 <= io_A_Valid_3_delay_51_11;
    io_A_Valid_3_delay_53_9 <= io_A_Valid_3_delay_52_10;
    io_A_Valid_3_delay_54_8 <= io_A_Valid_3_delay_53_9;
    io_A_Valid_3_delay_55_7 <= io_A_Valid_3_delay_54_8;
    io_A_Valid_3_delay_56_6 <= io_A_Valid_3_delay_55_7;
    io_A_Valid_3_delay_57_5 <= io_A_Valid_3_delay_56_6;
    io_A_Valid_3_delay_58_4 <= io_A_Valid_3_delay_57_5;
    io_A_Valid_3_delay_59_3 <= io_A_Valid_3_delay_58_4;
    io_A_Valid_3_delay_60_2 <= io_A_Valid_3_delay_59_3;
    io_A_Valid_3_delay_61_1 <= io_A_Valid_3_delay_60_2;
    io_A_Valid_3_delay_62 <= io_A_Valid_3_delay_61_1;
    io_B_Valid_62_delay_1_2 <= io_B_Valid_62;
    io_B_Valid_62_delay_2_1 <= io_B_Valid_62_delay_1_2;
    io_B_Valid_62_delay_3 <= io_B_Valid_62_delay_2_1;
    io_A_Valid_3_delay_1_62 <= io_A_Valid_3;
    io_A_Valid_3_delay_2_61 <= io_A_Valid_3_delay_1_62;
    io_A_Valid_3_delay_3_60 <= io_A_Valid_3_delay_2_61;
    io_A_Valid_3_delay_4_59 <= io_A_Valid_3_delay_3_60;
    io_A_Valid_3_delay_5_58 <= io_A_Valid_3_delay_4_59;
    io_A_Valid_3_delay_6_57 <= io_A_Valid_3_delay_5_58;
    io_A_Valid_3_delay_7_56 <= io_A_Valid_3_delay_6_57;
    io_A_Valid_3_delay_8_55 <= io_A_Valid_3_delay_7_56;
    io_A_Valid_3_delay_9_54 <= io_A_Valid_3_delay_8_55;
    io_A_Valid_3_delay_10_53 <= io_A_Valid_3_delay_9_54;
    io_A_Valid_3_delay_11_52 <= io_A_Valid_3_delay_10_53;
    io_A_Valid_3_delay_12_51 <= io_A_Valid_3_delay_11_52;
    io_A_Valid_3_delay_13_50 <= io_A_Valid_3_delay_12_51;
    io_A_Valid_3_delay_14_49 <= io_A_Valid_3_delay_13_50;
    io_A_Valid_3_delay_15_48 <= io_A_Valid_3_delay_14_49;
    io_A_Valid_3_delay_16_47 <= io_A_Valid_3_delay_15_48;
    io_A_Valid_3_delay_17_46 <= io_A_Valid_3_delay_16_47;
    io_A_Valid_3_delay_18_45 <= io_A_Valid_3_delay_17_46;
    io_A_Valid_3_delay_19_44 <= io_A_Valid_3_delay_18_45;
    io_A_Valid_3_delay_20_43 <= io_A_Valid_3_delay_19_44;
    io_A_Valid_3_delay_21_42 <= io_A_Valid_3_delay_20_43;
    io_A_Valid_3_delay_22_41 <= io_A_Valid_3_delay_21_42;
    io_A_Valid_3_delay_23_40 <= io_A_Valid_3_delay_22_41;
    io_A_Valid_3_delay_24_39 <= io_A_Valid_3_delay_23_40;
    io_A_Valid_3_delay_25_38 <= io_A_Valid_3_delay_24_39;
    io_A_Valid_3_delay_26_37 <= io_A_Valid_3_delay_25_38;
    io_A_Valid_3_delay_27_36 <= io_A_Valid_3_delay_26_37;
    io_A_Valid_3_delay_28_35 <= io_A_Valid_3_delay_27_36;
    io_A_Valid_3_delay_29_34 <= io_A_Valid_3_delay_28_35;
    io_A_Valid_3_delay_30_33 <= io_A_Valid_3_delay_29_34;
    io_A_Valid_3_delay_31_32 <= io_A_Valid_3_delay_30_33;
    io_A_Valid_3_delay_32_31 <= io_A_Valid_3_delay_31_32;
    io_A_Valid_3_delay_33_30 <= io_A_Valid_3_delay_32_31;
    io_A_Valid_3_delay_34_29 <= io_A_Valid_3_delay_33_30;
    io_A_Valid_3_delay_35_28 <= io_A_Valid_3_delay_34_29;
    io_A_Valid_3_delay_36_27 <= io_A_Valid_3_delay_35_28;
    io_A_Valid_3_delay_37_26 <= io_A_Valid_3_delay_36_27;
    io_A_Valid_3_delay_38_25 <= io_A_Valid_3_delay_37_26;
    io_A_Valid_3_delay_39_24 <= io_A_Valid_3_delay_38_25;
    io_A_Valid_3_delay_40_23 <= io_A_Valid_3_delay_39_24;
    io_A_Valid_3_delay_41_22 <= io_A_Valid_3_delay_40_23;
    io_A_Valid_3_delay_42_21 <= io_A_Valid_3_delay_41_22;
    io_A_Valid_3_delay_43_20 <= io_A_Valid_3_delay_42_21;
    io_A_Valid_3_delay_44_19 <= io_A_Valid_3_delay_43_20;
    io_A_Valid_3_delay_45_18 <= io_A_Valid_3_delay_44_19;
    io_A_Valid_3_delay_46_17 <= io_A_Valid_3_delay_45_18;
    io_A_Valid_3_delay_47_16 <= io_A_Valid_3_delay_46_17;
    io_A_Valid_3_delay_48_15 <= io_A_Valid_3_delay_47_16;
    io_A_Valid_3_delay_49_14 <= io_A_Valid_3_delay_48_15;
    io_A_Valid_3_delay_50_13 <= io_A_Valid_3_delay_49_14;
    io_A_Valid_3_delay_51_12 <= io_A_Valid_3_delay_50_13;
    io_A_Valid_3_delay_52_11 <= io_A_Valid_3_delay_51_12;
    io_A_Valid_3_delay_53_10 <= io_A_Valid_3_delay_52_11;
    io_A_Valid_3_delay_54_9 <= io_A_Valid_3_delay_53_10;
    io_A_Valid_3_delay_55_8 <= io_A_Valid_3_delay_54_9;
    io_A_Valid_3_delay_56_7 <= io_A_Valid_3_delay_55_8;
    io_A_Valid_3_delay_57_6 <= io_A_Valid_3_delay_56_7;
    io_A_Valid_3_delay_58_5 <= io_A_Valid_3_delay_57_6;
    io_A_Valid_3_delay_59_4 <= io_A_Valid_3_delay_58_5;
    io_A_Valid_3_delay_60_3 <= io_A_Valid_3_delay_59_4;
    io_A_Valid_3_delay_61_2 <= io_A_Valid_3_delay_60_3;
    io_A_Valid_3_delay_62_1 <= io_A_Valid_3_delay_61_2;
    io_A_Valid_3_delay_63 <= io_A_Valid_3_delay_62_1;
    io_B_Valid_63_delay_1_2 <= io_B_Valid_63;
    io_B_Valid_63_delay_2_1 <= io_B_Valid_63_delay_1_2;
    io_B_Valid_63_delay_3 <= io_B_Valid_63_delay_2_1;
    io_B_Valid_0_delay_1_3 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_2 <= io_B_Valid_0_delay_1_3;
    io_B_Valid_0_delay_3_1 <= io_B_Valid_0_delay_2_2;
    io_B_Valid_0_delay_4 <= io_B_Valid_0_delay_3_1;
    io_A_Valid_4_delay_1 <= io_A_Valid_4;
    io_B_Valid_1_delay_1_3 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_2 <= io_B_Valid_1_delay_1_3;
    io_B_Valid_1_delay_3_1 <= io_B_Valid_1_delay_2_2;
    io_B_Valid_1_delay_4 <= io_B_Valid_1_delay_3_1;
    io_A_Valid_4_delay_1_1 <= io_A_Valid_4;
    io_A_Valid_4_delay_2 <= io_A_Valid_4_delay_1_1;
    io_B_Valid_2_delay_1_3 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_2 <= io_B_Valid_2_delay_1_3;
    io_B_Valid_2_delay_3_1 <= io_B_Valid_2_delay_2_2;
    io_B_Valid_2_delay_4 <= io_B_Valid_2_delay_3_1;
    io_A_Valid_4_delay_1_2 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_1 <= io_A_Valid_4_delay_1_2;
    io_A_Valid_4_delay_3 <= io_A_Valid_4_delay_2_1;
    io_B_Valid_3_delay_1_3 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_2 <= io_B_Valid_3_delay_1_3;
    io_B_Valid_3_delay_3_1 <= io_B_Valid_3_delay_2_2;
    io_B_Valid_3_delay_4 <= io_B_Valid_3_delay_3_1;
    io_A_Valid_4_delay_1_3 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_2 <= io_A_Valid_4_delay_1_3;
    io_A_Valid_4_delay_3_1 <= io_A_Valid_4_delay_2_2;
    io_A_Valid_4_delay_4 <= io_A_Valid_4_delay_3_1;
    io_B_Valid_4_delay_1_3 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_2 <= io_B_Valid_4_delay_1_3;
    io_B_Valid_4_delay_3_1 <= io_B_Valid_4_delay_2_2;
    io_B_Valid_4_delay_4 <= io_B_Valid_4_delay_3_1;
    io_A_Valid_4_delay_1_4 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_3 <= io_A_Valid_4_delay_1_4;
    io_A_Valid_4_delay_3_2 <= io_A_Valid_4_delay_2_3;
    io_A_Valid_4_delay_4_1 <= io_A_Valid_4_delay_3_2;
    io_A_Valid_4_delay_5 <= io_A_Valid_4_delay_4_1;
    io_B_Valid_5_delay_1_3 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_2 <= io_B_Valid_5_delay_1_3;
    io_B_Valid_5_delay_3_1 <= io_B_Valid_5_delay_2_2;
    io_B_Valid_5_delay_4 <= io_B_Valid_5_delay_3_1;
    io_A_Valid_4_delay_1_5 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_4 <= io_A_Valid_4_delay_1_5;
    io_A_Valid_4_delay_3_3 <= io_A_Valid_4_delay_2_4;
    io_A_Valid_4_delay_4_2 <= io_A_Valid_4_delay_3_3;
    io_A_Valid_4_delay_5_1 <= io_A_Valid_4_delay_4_2;
    io_A_Valid_4_delay_6 <= io_A_Valid_4_delay_5_1;
    io_B_Valid_6_delay_1_3 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_2 <= io_B_Valid_6_delay_1_3;
    io_B_Valid_6_delay_3_1 <= io_B_Valid_6_delay_2_2;
    io_B_Valid_6_delay_4 <= io_B_Valid_6_delay_3_1;
    io_A_Valid_4_delay_1_6 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_5 <= io_A_Valid_4_delay_1_6;
    io_A_Valid_4_delay_3_4 <= io_A_Valid_4_delay_2_5;
    io_A_Valid_4_delay_4_3 <= io_A_Valid_4_delay_3_4;
    io_A_Valid_4_delay_5_2 <= io_A_Valid_4_delay_4_3;
    io_A_Valid_4_delay_6_1 <= io_A_Valid_4_delay_5_2;
    io_A_Valid_4_delay_7 <= io_A_Valid_4_delay_6_1;
    io_B_Valid_7_delay_1_3 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_2 <= io_B_Valid_7_delay_1_3;
    io_B_Valid_7_delay_3_1 <= io_B_Valid_7_delay_2_2;
    io_B_Valid_7_delay_4 <= io_B_Valid_7_delay_3_1;
    io_A_Valid_4_delay_1_7 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_6 <= io_A_Valid_4_delay_1_7;
    io_A_Valid_4_delay_3_5 <= io_A_Valid_4_delay_2_6;
    io_A_Valid_4_delay_4_4 <= io_A_Valid_4_delay_3_5;
    io_A_Valid_4_delay_5_3 <= io_A_Valid_4_delay_4_4;
    io_A_Valid_4_delay_6_2 <= io_A_Valid_4_delay_5_3;
    io_A_Valid_4_delay_7_1 <= io_A_Valid_4_delay_6_2;
    io_A_Valid_4_delay_8 <= io_A_Valid_4_delay_7_1;
    io_B_Valid_8_delay_1_3 <= io_B_Valid_8;
    io_B_Valid_8_delay_2_2 <= io_B_Valid_8_delay_1_3;
    io_B_Valid_8_delay_3_1 <= io_B_Valid_8_delay_2_2;
    io_B_Valid_8_delay_4 <= io_B_Valid_8_delay_3_1;
    io_A_Valid_4_delay_1_8 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_7 <= io_A_Valid_4_delay_1_8;
    io_A_Valid_4_delay_3_6 <= io_A_Valid_4_delay_2_7;
    io_A_Valid_4_delay_4_5 <= io_A_Valid_4_delay_3_6;
    io_A_Valid_4_delay_5_4 <= io_A_Valid_4_delay_4_5;
    io_A_Valid_4_delay_6_3 <= io_A_Valid_4_delay_5_4;
    io_A_Valid_4_delay_7_2 <= io_A_Valid_4_delay_6_3;
    io_A_Valid_4_delay_8_1 <= io_A_Valid_4_delay_7_2;
    io_A_Valid_4_delay_9 <= io_A_Valid_4_delay_8_1;
    io_B_Valid_9_delay_1_3 <= io_B_Valid_9;
    io_B_Valid_9_delay_2_2 <= io_B_Valid_9_delay_1_3;
    io_B_Valid_9_delay_3_1 <= io_B_Valid_9_delay_2_2;
    io_B_Valid_9_delay_4 <= io_B_Valid_9_delay_3_1;
    io_A_Valid_4_delay_1_9 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_8 <= io_A_Valid_4_delay_1_9;
    io_A_Valid_4_delay_3_7 <= io_A_Valid_4_delay_2_8;
    io_A_Valid_4_delay_4_6 <= io_A_Valid_4_delay_3_7;
    io_A_Valid_4_delay_5_5 <= io_A_Valid_4_delay_4_6;
    io_A_Valid_4_delay_6_4 <= io_A_Valid_4_delay_5_5;
    io_A_Valid_4_delay_7_3 <= io_A_Valid_4_delay_6_4;
    io_A_Valid_4_delay_8_2 <= io_A_Valid_4_delay_7_3;
    io_A_Valid_4_delay_9_1 <= io_A_Valid_4_delay_8_2;
    io_A_Valid_4_delay_10 <= io_A_Valid_4_delay_9_1;
    io_B_Valid_10_delay_1_3 <= io_B_Valid_10;
    io_B_Valid_10_delay_2_2 <= io_B_Valid_10_delay_1_3;
    io_B_Valid_10_delay_3_1 <= io_B_Valid_10_delay_2_2;
    io_B_Valid_10_delay_4 <= io_B_Valid_10_delay_3_1;
    io_A_Valid_4_delay_1_10 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_9 <= io_A_Valid_4_delay_1_10;
    io_A_Valid_4_delay_3_8 <= io_A_Valid_4_delay_2_9;
    io_A_Valid_4_delay_4_7 <= io_A_Valid_4_delay_3_8;
    io_A_Valid_4_delay_5_6 <= io_A_Valid_4_delay_4_7;
    io_A_Valid_4_delay_6_5 <= io_A_Valid_4_delay_5_6;
    io_A_Valid_4_delay_7_4 <= io_A_Valid_4_delay_6_5;
    io_A_Valid_4_delay_8_3 <= io_A_Valid_4_delay_7_4;
    io_A_Valid_4_delay_9_2 <= io_A_Valid_4_delay_8_3;
    io_A_Valid_4_delay_10_1 <= io_A_Valid_4_delay_9_2;
    io_A_Valid_4_delay_11 <= io_A_Valid_4_delay_10_1;
    io_B_Valid_11_delay_1_3 <= io_B_Valid_11;
    io_B_Valid_11_delay_2_2 <= io_B_Valid_11_delay_1_3;
    io_B_Valid_11_delay_3_1 <= io_B_Valid_11_delay_2_2;
    io_B_Valid_11_delay_4 <= io_B_Valid_11_delay_3_1;
    io_A_Valid_4_delay_1_11 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_10 <= io_A_Valid_4_delay_1_11;
    io_A_Valid_4_delay_3_9 <= io_A_Valid_4_delay_2_10;
    io_A_Valid_4_delay_4_8 <= io_A_Valid_4_delay_3_9;
    io_A_Valid_4_delay_5_7 <= io_A_Valid_4_delay_4_8;
    io_A_Valid_4_delay_6_6 <= io_A_Valid_4_delay_5_7;
    io_A_Valid_4_delay_7_5 <= io_A_Valid_4_delay_6_6;
    io_A_Valid_4_delay_8_4 <= io_A_Valid_4_delay_7_5;
    io_A_Valid_4_delay_9_3 <= io_A_Valid_4_delay_8_4;
    io_A_Valid_4_delay_10_2 <= io_A_Valid_4_delay_9_3;
    io_A_Valid_4_delay_11_1 <= io_A_Valid_4_delay_10_2;
    io_A_Valid_4_delay_12 <= io_A_Valid_4_delay_11_1;
    io_B_Valid_12_delay_1_3 <= io_B_Valid_12;
    io_B_Valid_12_delay_2_2 <= io_B_Valid_12_delay_1_3;
    io_B_Valid_12_delay_3_1 <= io_B_Valid_12_delay_2_2;
    io_B_Valid_12_delay_4 <= io_B_Valid_12_delay_3_1;
    io_A_Valid_4_delay_1_12 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_11 <= io_A_Valid_4_delay_1_12;
    io_A_Valid_4_delay_3_10 <= io_A_Valid_4_delay_2_11;
    io_A_Valid_4_delay_4_9 <= io_A_Valid_4_delay_3_10;
    io_A_Valid_4_delay_5_8 <= io_A_Valid_4_delay_4_9;
    io_A_Valid_4_delay_6_7 <= io_A_Valid_4_delay_5_8;
    io_A_Valid_4_delay_7_6 <= io_A_Valid_4_delay_6_7;
    io_A_Valid_4_delay_8_5 <= io_A_Valid_4_delay_7_6;
    io_A_Valid_4_delay_9_4 <= io_A_Valid_4_delay_8_5;
    io_A_Valid_4_delay_10_3 <= io_A_Valid_4_delay_9_4;
    io_A_Valid_4_delay_11_2 <= io_A_Valid_4_delay_10_3;
    io_A_Valid_4_delay_12_1 <= io_A_Valid_4_delay_11_2;
    io_A_Valid_4_delay_13 <= io_A_Valid_4_delay_12_1;
    io_B_Valid_13_delay_1_3 <= io_B_Valid_13;
    io_B_Valid_13_delay_2_2 <= io_B_Valid_13_delay_1_3;
    io_B_Valid_13_delay_3_1 <= io_B_Valid_13_delay_2_2;
    io_B_Valid_13_delay_4 <= io_B_Valid_13_delay_3_1;
    io_A_Valid_4_delay_1_13 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_12 <= io_A_Valid_4_delay_1_13;
    io_A_Valid_4_delay_3_11 <= io_A_Valid_4_delay_2_12;
    io_A_Valid_4_delay_4_10 <= io_A_Valid_4_delay_3_11;
    io_A_Valid_4_delay_5_9 <= io_A_Valid_4_delay_4_10;
    io_A_Valid_4_delay_6_8 <= io_A_Valid_4_delay_5_9;
    io_A_Valid_4_delay_7_7 <= io_A_Valid_4_delay_6_8;
    io_A_Valid_4_delay_8_6 <= io_A_Valid_4_delay_7_7;
    io_A_Valid_4_delay_9_5 <= io_A_Valid_4_delay_8_6;
    io_A_Valid_4_delay_10_4 <= io_A_Valid_4_delay_9_5;
    io_A_Valid_4_delay_11_3 <= io_A_Valid_4_delay_10_4;
    io_A_Valid_4_delay_12_2 <= io_A_Valid_4_delay_11_3;
    io_A_Valid_4_delay_13_1 <= io_A_Valid_4_delay_12_2;
    io_A_Valid_4_delay_14 <= io_A_Valid_4_delay_13_1;
    io_B_Valid_14_delay_1_3 <= io_B_Valid_14;
    io_B_Valid_14_delay_2_2 <= io_B_Valid_14_delay_1_3;
    io_B_Valid_14_delay_3_1 <= io_B_Valid_14_delay_2_2;
    io_B_Valid_14_delay_4 <= io_B_Valid_14_delay_3_1;
    io_A_Valid_4_delay_1_14 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_13 <= io_A_Valid_4_delay_1_14;
    io_A_Valid_4_delay_3_12 <= io_A_Valid_4_delay_2_13;
    io_A_Valid_4_delay_4_11 <= io_A_Valid_4_delay_3_12;
    io_A_Valid_4_delay_5_10 <= io_A_Valid_4_delay_4_11;
    io_A_Valid_4_delay_6_9 <= io_A_Valid_4_delay_5_10;
    io_A_Valid_4_delay_7_8 <= io_A_Valid_4_delay_6_9;
    io_A_Valid_4_delay_8_7 <= io_A_Valid_4_delay_7_8;
    io_A_Valid_4_delay_9_6 <= io_A_Valid_4_delay_8_7;
    io_A_Valid_4_delay_10_5 <= io_A_Valid_4_delay_9_6;
    io_A_Valid_4_delay_11_4 <= io_A_Valid_4_delay_10_5;
    io_A_Valid_4_delay_12_3 <= io_A_Valid_4_delay_11_4;
    io_A_Valid_4_delay_13_2 <= io_A_Valid_4_delay_12_3;
    io_A_Valid_4_delay_14_1 <= io_A_Valid_4_delay_13_2;
    io_A_Valid_4_delay_15 <= io_A_Valid_4_delay_14_1;
    io_B_Valid_15_delay_1_3 <= io_B_Valid_15;
    io_B_Valid_15_delay_2_2 <= io_B_Valid_15_delay_1_3;
    io_B_Valid_15_delay_3_1 <= io_B_Valid_15_delay_2_2;
    io_B_Valid_15_delay_4 <= io_B_Valid_15_delay_3_1;
    io_A_Valid_4_delay_1_15 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_14 <= io_A_Valid_4_delay_1_15;
    io_A_Valid_4_delay_3_13 <= io_A_Valid_4_delay_2_14;
    io_A_Valid_4_delay_4_12 <= io_A_Valid_4_delay_3_13;
    io_A_Valid_4_delay_5_11 <= io_A_Valid_4_delay_4_12;
    io_A_Valid_4_delay_6_10 <= io_A_Valid_4_delay_5_11;
    io_A_Valid_4_delay_7_9 <= io_A_Valid_4_delay_6_10;
    io_A_Valid_4_delay_8_8 <= io_A_Valid_4_delay_7_9;
    io_A_Valid_4_delay_9_7 <= io_A_Valid_4_delay_8_8;
    io_A_Valid_4_delay_10_6 <= io_A_Valid_4_delay_9_7;
    io_A_Valid_4_delay_11_5 <= io_A_Valid_4_delay_10_6;
    io_A_Valid_4_delay_12_4 <= io_A_Valid_4_delay_11_5;
    io_A_Valid_4_delay_13_3 <= io_A_Valid_4_delay_12_4;
    io_A_Valid_4_delay_14_2 <= io_A_Valid_4_delay_13_3;
    io_A_Valid_4_delay_15_1 <= io_A_Valid_4_delay_14_2;
    io_A_Valid_4_delay_16 <= io_A_Valid_4_delay_15_1;
    io_B_Valid_16_delay_1_3 <= io_B_Valid_16;
    io_B_Valid_16_delay_2_2 <= io_B_Valid_16_delay_1_3;
    io_B_Valid_16_delay_3_1 <= io_B_Valid_16_delay_2_2;
    io_B_Valid_16_delay_4 <= io_B_Valid_16_delay_3_1;
    io_A_Valid_4_delay_1_16 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_15 <= io_A_Valid_4_delay_1_16;
    io_A_Valid_4_delay_3_14 <= io_A_Valid_4_delay_2_15;
    io_A_Valid_4_delay_4_13 <= io_A_Valid_4_delay_3_14;
    io_A_Valid_4_delay_5_12 <= io_A_Valid_4_delay_4_13;
    io_A_Valid_4_delay_6_11 <= io_A_Valid_4_delay_5_12;
    io_A_Valid_4_delay_7_10 <= io_A_Valid_4_delay_6_11;
    io_A_Valid_4_delay_8_9 <= io_A_Valid_4_delay_7_10;
    io_A_Valid_4_delay_9_8 <= io_A_Valid_4_delay_8_9;
    io_A_Valid_4_delay_10_7 <= io_A_Valid_4_delay_9_8;
    io_A_Valid_4_delay_11_6 <= io_A_Valid_4_delay_10_7;
    io_A_Valid_4_delay_12_5 <= io_A_Valid_4_delay_11_6;
    io_A_Valid_4_delay_13_4 <= io_A_Valid_4_delay_12_5;
    io_A_Valid_4_delay_14_3 <= io_A_Valid_4_delay_13_4;
    io_A_Valid_4_delay_15_2 <= io_A_Valid_4_delay_14_3;
    io_A_Valid_4_delay_16_1 <= io_A_Valid_4_delay_15_2;
    io_A_Valid_4_delay_17 <= io_A_Valid_4_delay_16_1;
    io_B_Valid_17_delay_1_3 <= io_B_Valid_17;
    io_B_Valid_17_delay_2_2 <= io_B_Valid_17_delay_1_3;
    io_B_Valid_17_delay_3_1 <= io_B_Valid_17_delay_2_2;
    io_B_Valid_17_delay_4 <= io_B_Valid_17_delay_3_1;
    io_A_Valid_4_delay_1_17 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_16 <= io_A_Valid_4_delay_1_17;
    io_A_Valid_4_delay_3_15 <= io_A_Valid_4_delay_2_16;
    io_A_Valid_4_delay_4_14 <= io_A_Valid_4_delay_3_15;
    io_A_Valid_4_delay_5_13 <= io_A_Valid_4_delay_4_14;
    io_A_Valid_4_delay_6_12 <= io_A_Valid_4_delay_5_13;
    io_A_Valid_4_delay_7_11 <= io_A_Valid_4_delay_6_12;
    io_A_Valid_4_delay_8_10 <= io_A_Valid_4_delay_7_11;
    io_A_Valid_4_delay_9_9 <= io_A_Valid_4_delay_8_10;
    io_A_Valid_4_delay_10_8 <= io_A_Valid_4_delay_9_9;
    io_A_Valid_4_delay_11_7 <= io_A_Valid_4_delay_10_8;
    io_A_Valid_4_delay_12_6 <= io_A_Valid_4_delay_11_7;
    io_A_Valid_4_delay_13_5 <= io_A_Valid_4_delay_12_6;
    io_A_Valid_4_delay_14_4 <= io_A_Valid_4_delay_13_5;
    io_A_Valid_4_delay_15_3 <= io_A_Valid_4_delay_14_4;
    io_A_Valid_4_delay_16_2 <= io_A_Valid_4_delay_15_3;
    io_A_Valid_4_delay_17_1 <= io_A_Valid_4_delay_16_2;
    io_A_Valid_4_delay_18 <= io_A_Valid_4_delay_17_1;
    io_B_Valid_18_delay_1_3 <= io_B_Valid_18;
    io_B_Valid_18_delay_2_2 <= io_B_Valid_18_delay_1_3;
    io_B_Valid_18_delay_3_1 <= io_B_Valid_18_delay_2_2;
    io_B_Valid_18_delay_4 <= io_B_Valid_18_delay_3_1;
    io_A_Valid_4_delay_1_18 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_17 <= io_A_Valid_4_delay_1_18;
    io_A_Valid_4_delay_3_16 <= io_A_Valid_4_delay_2_17;
    io_A_Valid_4_delay_4_15 <= io_A_Valid_4_delay_3_16;
    io_A_Valid_4_delay_5_14 <= io_A_Valid_4_delay_4_15;
    io_A_Valid_4_delay_6_13 <= io_A_Valid_4_delay_5_14;
    io_A_Valid_4_delay_7_12 <= io_A_Valid_4_delay_6_13;
    io_A_Valid_4_delay_8_11 <= io_A_Valid_4_delay_7_12;
    io_A_Valid_4_delay_9_10 <= io_A_Valid_4_delay_8_11;
    io_A_Valid_4_delay_10_9 <= io_A_Valid_4_delay_9_10;
    io_A_Valid_4_delay_11_8 <= io_A_Valid_4_delay_10_9;
    io_A_Valid_4_delay_12_7 <= io_A_Valid_4_delay_11_8;
    io_A_Valid_4_delay_13_6 <= io_A_Valid_4_delay_12_7;
    io_A_Valid_4_delay_14_5 <= io_A_Valid_4_delay_13_6;
    io_A_Valid_4_delay_15_4 <= io_A_Valid_4_delay_14_5;
    io_A_Valid_4_delay_16_3 <= io_A_Valid_4_delay_15_4;
    io_A_Valid_4_delay_17_2 <= io_A_Valid_4_delay_16_3;
    io_A_Valid_4_delay_18_1 <= io_A_Valid_4_delay_17_2;
    io_A_Valid_4_delay_19 <= io_A_Valid_4_delay_18_1;
    io_B_Valid_19_delay_1_3 <= io_B_Valid_19;
    io_B_Valid_19_delay_2_2 <= io_B_Valid_19_delay_1_3;
    io_B_Valid_19_delay_3_1 <= io_B_Valid_19_delay_2_2;
    io_B_Valid_19_delay_4 <= io_B_Valid_19_delay_3_1;
    io_A_Valid_4_delay_1_19 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_18 <= io_A_Valid_4_delay_1_19;
    io_A_Valid_4_delay_3_17 <= io_A_Valid_4_delay_2_18;
    io_A_Valid_4_delay_4_16 <= io_A_Valid_4_delay_3_17;
    io_A_Valid_4_delay_5_15 <= io_A_Valid_4_delay_4_16;
    io_A_Valid_4_delay_6_14 <= io_A_Valid_4_delay_5_15;
    io_A_Valid_4_delay_7_13 <= io_A_Valid_4_delay_6_14;
    io_A_Valid_4_delay_8_12 <= io_A_Valid_4_delay_7_13;
    io_A_Valid_4_delay_9_11 <= io_A_Valid_4_delay_8_12;
    io_A_Valid_4_delay_10_10 <= io_A_Valid_4_delay_9_11;
    io_A_Valid_4_delay_11_9 <= io_A_Valid_4_delay_10_10;
    io_A_Valid_4_delay_12_8 <= io_A_Valid_4_delay_11_9;
    io_A_Valid_4_delay_13_7 <= io_A_Valid_4_delay_12_8;
    io_A_Valid_4_delay_14_6 <= io_A_Valid_4_delay_13_7;
    io_A_Valid_4_delay_15_5 <= io_A_Valid_4_delay_14_6;
    io_A_Valid_4_delay_16_4 <= io_A_Valid_4_delay_15_5;
    io_A_Valid_4_delay_17_3 <= io_A_Valid_4_delay_16_4;
    io_A_Valid_4_delay_18_2 <= io_A_Valid_4_delay_17_3;
    io_A_Valid_4_delay_19_1 <= io_A_Valid_4_delay_18_2;
    io_A_Valid_4_delay_20 <= io_A_Valid_4_delay_19_1;
    io_B_Valid_20_delay_1_3 <= io_B_Valid_20;
    io_B_Valid_20_delay_2_2 <= io_B_Valid_20_delay_1_3;
    io_B_Valid_20_delay_3_1 <= io_B_Valid_20_delay_2_2;
    io_B_Valid_20_delay_4 <= io_B_Valid_20_delay_3_1;
    io_A_Valid_4_delay_1_20 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_19 <= io_A_Valid_4_delay_1_20;
    io_A_Valid_4_delay_3_18 <= io_A_Valid_4_delay_2_19;
    io_A_Valid_4_delay_4_17 <= io_A_Valid_4_delay_3_18;
    io_A_Valid_4_delay_5_16 <= io_A_Valid_4_delay_4_17;
    io_A_Valid_4_delay_6_15 <= io_A_Valid_4_delay_5_16;
    io_A_Valid_4_delay_7_14 <= io_A_Valid_4_delay_6_15;
    io_A_Valid_4_delay_8_13 <= io_A_Valid_4_delay_7_14;
    io_A_Valid_4_delay_9_12 <= io_A_Valid_4_delay_8_13;
    io_A_Valid_4_delay_10_11 <= io_A_Valid_4_delay_9_12;
    io_A_Valid_4_delay_11_10 <= io_A_Valid_4_delay_10_11;
    io_A_Valid_4_delay_12_9 <= io_A_Valid_4_delay_11_10;
    io_A_Valid_4_delay_13_8 <= io_A_Valid_4_delay_12_9;
    io_A_Valid_4_delay_14_7 <= io_A_Valid_4_delay_13_8;
    io_A_Valid_4_delay_15_6 <= io_A_Valid_4_delay_14_7;
    io_A_Valid_4_delay_16_5 <= io_A_Valid_4_delay_15_6;
    io_A_Valid_4_delay_17_4 <= io_A_Valid_4_delay_16_5;
    io_A_Valid_4_delay_18_3 <= io_A_Valid_4_delay_17_4;
    io_A_Valid_4_delay_19_2 <= io_A_Valid_4_delay_18_3;
    io_A_Valid_4_delay_20_1 <= io_A_Valid_4_delay_19_2;
    io_A_Valid_4_delay_21 <= io_A_Valid_4_delay_20_1;
    io_B_Valid_21_delay_1_3 <= io_B_Valid_21;
    io_B_Valid_21_delay_2_2 <= io_B_Valid_21_delay_1_3;
    io_B_Valid_21_delay_3_1 <= io_B_Valid_21_delay_2_2;
    io_B_Valid_21_delay_4 <= io_B_Valid_21_delay_3_1;
    io_A_Valid_4_delay_1_21 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_20 <= io_A_Valid_4_delay_1_21;
    io_A_Valid_4_delay_3_19 <= io_A_Valid_4_delay_2_20;
    io_A_Valid_4_delay_4_18 <= io_A_Valid_4_delay_3_19;
    io_A_Valid_4_delay_5_17 <= io_A_Valid_4_delay_4_18;
    io_A_Valid_4_delay_6_16 <= io_A_Valid_4_delay_5_17;
    io_A_Valid_4_delay_7_15 <= io_A_Valid_4_delay_6_16;
    io_A_Valid_4_delay_8_14 <= io_A_Valid_4_delay_7_15;
    io_A_Valid_4_delay_9_13 <= io_A_Valid_4_delay_8_14;
    io_A_Valid_4_delay_10_12 <= io_A_Valid_4_delay_9_13;
    io_A_Valid_4_delay_11_11 <= io_A_Valid_4_delay_10_12;
    io_A_Valid_4_delay_12_10 <= io_A_Valid_4_delay_11_11;
    io_A_Valid_4_delay_13_9 <= io_A_Valid_4_delay_12_10;
    io_A_Valid_4_delay_14_8 <= io_A_Valid_4_delay_13_9;
    io_A_Valid_4_delay_15_7 <= io_A_Valid_4_delay_14_8;
    io_A_Valid_4_delay_16_6 <= io_A_Valid_4_delay_15_7;
    io_A_Valid_4_delay_17_5 <= io_A_Valid_4_delay_16_6;
    io_A_Valid_4_delay_18_4 <= io_A_Valid_4_delay_17_5;
    io_A_Valid_4_delay_19_3 <= io_A_Valid_4_delay_18_4;
    io_A_Valid_4_delay_20_2 <= io_A_Valid_4_delay_19_3;
    io_A_Valid_4_delay_21_1 <= io_A_Valid_4_delay_20_2;
    io_A_Valid_4_delay_22 <= io_A_Valid_4_delay_21_1;
    io_B_Valid_22_delay_1_3 <= io_B_Valid_22;
    io_B_Valid_22_delay_2_2 <= io_B_Valid_22_delay_1_3;
    io_B_Valid_22_delay_3_1 <= io_B_Valid_22_delay_2_2;
    io_B_Valid_22_delay_4 <= io_B_Valid_22_delay_3_1;
    io_A_Valid_4_delay_1_22 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_21 <= io_A_Valid_4_delay_1_22;
    io_A_Valid_4_delay_3_20 <= io_A_Valid_4_delay_2_21;
    io_A_Valid_4_delay_4_19 <= io_A_Valid_4_delay_3_20;
    io_A_Valid_4_delay_5_18 <= io_A_Valid_4_delay_4_19;
    io_A_Valid_4_delay_6_17 <= io_A_Valid_4_delay_5_18;
    io_A_Valid_4_delay_7_16 <= io_A_Valid_4_delay_6_17;
    io_A_Valid_4_delay_8_15 <= io_A_Valid_4_delay_7_16;
    io_A_Valid_4_delay_9_14 <= io_A_Valid_4_delay_8_15;
    io_A_Valid_4_delay_10_13 <= io_A_Valid_4_delay_9_14;
    io_A_Valid_4_delay_11_12 <= io_A_Valid_4_delay_10_13;
    io_A_Valid_4_delay_12_11 <= io_A_Valid_4_delay_11_12;
    io_A_Valid_4_delay_13_10 <= io_A_Valid_4_delay_12_11;
    io_A_Valid_4_delay_14_9 <= io_A_Valid_4_delay_13_10;
    io_A_Valid_4_delay_15_8 <= io_A_Valid_4_delay_14_9;
    io_A_Valid_4_delay_16_7 <= io_A_Valid_4_delay_15_8;
    io_A_Valid_4_delay_17_6 <= io_A_Valid_4_delay_16_7;
    io_A_Valid_4_delay_18_5 <= io_A_Valid_4_delay_17_6;
    io_A_Valid_4_delay_19_4 <= io_A_Valid_4_delay_18_5;
    io_A_Valid_4_delay_20_3 <= io_A_Valid_4_delay_19_4;
    io_A_Valid_4_delay_21_2 <= io_A_Valid_4_delay_20_3;
    io_A_Valid_4_delay_22_1 <= io_A_Valid_4_delay_21_2;
    io_A_Valid_4_delay_23 <= io_A_Valid_4_delay_22_1;
    io_B_Valid_23_delay_1_3 <= io_B_Valid_23;
    io_B_Valid_23_delay_2_2 <= io_B_Valid_23_delay_1_3;
    io_B_Valid_23_delay_3_1 <= io_B_Valid_23_delay_2_2;
    io_B_Valid_23_delay_4 <= io_B_Valid_23_delay_3_1;
    io_A_Valid_4_delay_1_23 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_22 <= io_A_Valid_4_delay_1_23;
    io_A_Valid_4_delay_3_21 <= io_A_Valid_4_delay_2_22;
    io_A_Valid_4_delay_4_20 <= io_A_Valid_4_delay_3_21;
    io_A_Valid_4_delay_5_19 <= io_A_Valid_4_delay_4_20;
    io_A_Valid_4_delay_6_18 <= io_A_Valid_4_delay_5_19;
    io_A_Valid_4_delay_7_17 <= io_A_Valid_4_delay_6_18;
    io_A_Valid_4_delay_8_16 <= io_A_Valid_4_delay_7_17;
    io_A_Valid_4_delay_9_15 <= io_A_Valid_4_delay_8_16;
    io_A_Valid_4_delay_10_14 <= io_A_Valid_4_delay_9_15;
    io_A_Valid_4_delay_11_13 <= io_A_Valid_4_delay_10_14;
    io_A_Valid_4_delay_12_12 <= io_A_Valid_4_delay_11_13;
    io_A_Valid_4_delay_13_11 <= io_A_Valid_4_delay_12_12;
    io_A_Valid_4_delay_14_10 <= io_A_Valid_4_delay_13_11;
    io_A_Valid_4_delay_15_9 <= io_A_Valid_4_delay_14_10;
    io_A_Valid_4_delay_16_8 <= io_A_Valid_4_delay_15_9;
    io_A_Valid_4_delay_17_7 <= io_A_Valid_4_delay_16_8;
    io_A_Valid_4_delay_18_6 <= io_A_Valid_4_delay_17_7;
    io_A_Valid_4_delay_19_5 <= io_A_Valid_4_delay_18_6;
    io_A_Valid_4_delay_20_4 <= io_A_Valid_4_delay_19_5;
    io_A_Valid_4_delay_21_3 <= io_A_Valid_4_delay_20_4;
    io_A_Valid_4_delay_22_2 <= io_A_Valid_4_delay_21_3;
    io_A_Valid_4_delay_23_1 <= io_A_Valid_4_delay_22_2;
    io_A_Valid_4_delay_24 <= io_A_Valid_4_delay_23_1;
    io_B_Valid_24_delay_1_3 <= io_B_Valid_24;
    io_B_Valid_24_delay_2_2 <= io_B_Valid_24_delay_1_3;
    io_B_Valid_24_delay_3_1 <= io_B_Valid_24_delay_2_2;
    io_B_Valid_24_delay_4 <= io_B_Valid_24_delay_3_1;
    io_A_Valid_4_delay_1_24 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_23 <= io_A_Valid_4_delay_1_24;
    io_A_Valid_4_delay_3_22 <= io_A_Valid_4_delay_2_23;
    io_A_Valid_4_delay_4_21 <= io_A_Valid_4_delay_3_22;
    io_A_Valid_4_delay_5_20 <= io_A_Valid_4_delay_4_21;
    io_A_Valid_4_delay_6_19 <= io_A_Valid_4_delay_5_20;
    io_A_Valid_4_delay_7_18 <= io_A_Valid_4_delay_6_19;
    io_A_Valid_4_delay_8_17 <= io_A_Valid_4_delay_7_18;
    io_A_Valid_4_delay_9_16 <= io_A_Valid_4_delay_8_17;
    io_A_Valid_4_delay_10_15 <= io_A_Valid_4_delay_9_16;
    io_A_Valid_4_delay_11_14 <= io_A_Valid_4_delay_10_15;
    io_A_Valid_4_delay_12_13 <= io_A_Valid_4_delay_11_14;
    io_A_Valid_4_delay_13_12 <= io_A_Valid_4_delay_12_13;
    io_A_Valid_4_delay_14_11 <= io_A_Valid_4_delay_13_12;
    io_A_Valid_4_delay_15_10 <= io_A_Valid_4_delay_14_11;
    io_A_Valid_4_delay_16_9 <= io_A_Valid_4_delay_15_10;
    io_A_Valid_4_delay_17_8 <= io_A_Valid_4_delay_16_9;
    io_A_Valid_4_delay_18_7 <= io_A_Valid_4_delay_17_8;
    io_A_Valid_4_delay_19_6 <= io_A_Valid_4_delay_18_7;
    io_A_Valid_4_delay_20_5 <= io_A_Valid_4_delay_19_6;
    io_A_Valid_4_delay_21_4 <= io_A_Valid_4_delay_20_5;
    io_A_Valid_4_delay_22_3 <= io_A_Valid_4_delay_21_4;
    io_A_Valid_4_delay_23_2 <= io_A_Valid_4_delay_22_3;
    io_A_Valid_4_delay_24_1 <= io_A_Valid_4_delay_23_2;
    io_A_Valid_4_delay_25 <= io_A_Valid_4_delay_24_1;
    io_B_Valid_25_delay_1_3 <= io_B_Valid_25;
    io_B_Valid_25_delay_2_2 <= io_B_Valid_25_delay_1_3;
    io_B_Valid_25_delay_3_1 <= io_B_Valid_25_delay_2_2;
    io_B_Valid_25_delay_4 <= io_B_Valid_25_delay_3_1;
    io_A_Valid_4_delay_1_25 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_24 <= io_A_Valid_4_delay_1_25;
    io_A_Valid_4_delay_3_23 <= io_A_Valid_4_delay_2_24;
    io_A_Valid_4_delay_4_22 <= io_A_Valid_4_delay_3_23;
    io_A_Valid_4_delay_5_21 <= io_A_Valid_4_delay_4_22;
    io_A_Valid_4_delay_6_20 <= io_A_Valid_4_delay_5_21;
    io_A_Valid_4_delay_7_19 <= io_A_Valid_4_delay_6_20;
    io_A_Valid_4_delay_8_18 <= io_A_Valid_4_delay_7_19;
    io_A_Valid_4_delay_9_17 <= io_A_Valid_4_delay_8_18;
    io_A_Valid_4_delay_10_16 <= io_A_Valid_4_delay_9_17;
    io_A_Valid_4_delay_11_15 <= io_A_Valid_4_delay_10_16;
    io_A_Valid_4_delay_12_14 <= io_A_Valid_4_delay_11_15;
    io_A_Valid_4_delay_13_13 <= io_A_Valid_4_delay_12_14;
    io_A_Valid_4_delay_14_12 <= io_A_Valid_4_delay_13_13;
    io_A_Valid_4_delay_15_11 <= io_A_Valid_4_delay_14_12;
    io_A_Valid_4_delay_16_10 <= io_A_Valid_4_delay_15_11;
    io_A_Valid_4_delay_17_9 <= io_A_Valid_4_delay_16_10;
    io_A_Valid_4_delay_18_8 <= io_A_Valid_4_delay_17_9;
    io_A_Valid_4_delay_19_7 <= io_A_Valid_4_delay_18_8;
    io_A_Valid_4_delay_20_6 <= io_A_Valid_4_delay_19_7;
    io_A_Valid_4_delay_21_5 <= io_A_Valid_4_delay_20_6;
    io_A_Valid_4_delay_22_4 <= io_A_Valid_4_delay_21_5;
    io_A_Valid_4_delay_23_3 <= io_A_Valid_4_delay_22_4;
    io_A_Valid_4_delay_24_2 <= io_A_Valid_4_delay_23_3;
    io_A_Valid_4_delay_25_1 <= io_A_Valid_4_delay_24_2;
    io_A_Valid_4_delay_26 <= io_A_Valid_4_delay_25_1;
    io_B_Valid_26_delay_1_3 <= io_B_Valid_26;
    io_B_Valid_26_delay_2_2 <= io_B_Valid_26_delay_1_3;
    io_B_Valid_26_delay_3_1 <= io_B_Valid_26_delay_2_2;
    io_B_Valid_26_delay_4 <= io_B_Valid_26_delay_3_1;
    io_A_Valid_4_delay_1_26 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_25 <= io_A_Valid_4_delay_1_26;
    io_A_Valid_4_delay_3_24 <= io_A_Valid_4_delay_2_25;
    io_A_Valid_4_delay_4_23 <= io_A_Valid_4_delay_3_24;
    io_A_Valid_4_delay_5_22 <= io_A_Valid_4_delay_4_23;
    io_A_Valid_4_delay_6_21 <= io_A_Valid_4_delay_5_22;
    io_A_Valid_4_delay_7_20 <= io_A_Valid_4_delay_6_21;
    io_A_Valid_4_delay_8_19 <= io_A_Valid_4_delay_7_20;
    io_A_Valid_4_delay_9_18 <= io_A_Valid_4_delay_8_19;
    io_A_Valid_4_delay_10_17 <= io_A_Valid_4_delay_9_18;
    io_A_Valid_4_delay_11_16 <= io_A_Valid_4_delay_10_17;
    io_A_Valid_4_delay_12_15 <= io_A_Valid_4_delay_11_16;
    io_A_Valid_4_delay_13_14 <= io_A_Valid_4_delay_12_15;
    io_A_Valid_4_delay_14_13 <= io_A_Valid_4_delay_13_14;
    io_A_Valid_4_delay_15_12 <= io_A_Valid_4_delay_14_13;
    io_A_Valid_4_delay_16_11 <= io_A_Valid_4_delay_15_12;
    io_A_Valid_4_delay_17_10 <= io_A_Valid_4_delay_16_11;
    io_A_Valid_4_delay_18_9 <= io_A_Valid_4_delay_17_10;
    io_A_Valid_4_delay_19_8 <= io_A_Valid_4_delay_18_9;
    io_A_Valid_4_delay_20_7 <= io_A_Valid_4_delay_19_8;
    io_A_Valid_4_delay_21_6 <= io_A_Valid_4_delay_20_7;
    io_A_Valid_4_delay_22_5 <= io_A_Valid_4_delay_21_6;
    io_A_Valid_4_delay_23_4 <= io_A_Valid_4_delay_22_5;
    io_A_Valid_4_delay_24_3 <= io_A_Valid_4_delay_23_4;
    io_A_Valid_4_delay_25_2 <= io_A_Valid_4_delay_24_3;
    io_A_Valid_4_delay_26_1 <= io_A_Valid_4_delay_25_2;
    io_A_Valid_4_delay_27 <= io_A_Valid_4_delay_26_1;
    io_B_Valid_27_delay_1_3 <= io_B_Valid_27;
    io_B_Valid_27_delay_2_2 <= io_B_Valid_27_delay_1_3;
    io_B_Valid_27_delay_3_1 <= io_B_Valid_27_delay_2_2;
    io_B_Valid_27_delay_4 <= io_B_Valid_27_delay_3_1;
    io_A_Valid_4_delay_1_27 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_26 <= io_A_Valid_4_delay_1_27;
    io_A_Valid_4_delay_3_25 <= io_A_Valid_4_delay_2_26;
    io_A_Valid_4_delay_4_24 <= io_A_Valid_4_delay_3_25;
    io_A_Valid_4_delay_5_23 <= io_A_Valid_4_delay_4_24;
    io_A_Valid_4_delay_6_22 <= io_A_Valid_4_delay_5_23;
    io_A_Valid_4_delay_7_21 <= io_A_Valid_4_delay_6_22;
    io_A_Valid_4_delay_8_20 <= io_A_Valid_4_delay_7_21;
    io_A_Valid_4_delay_9_19 <= io_A_Valid_4_delay_8_20;
    io_A_Valid_4_delay_10_18 <= io_A_Valid_4_delay_9_19;
    io_A_Valid_4_delay_11_17 <= io_A_Valid_4_delay_10_18;
    io_A_Valid_4_delay_12_16 <= io_A_Valid_4_delay_11_17;
    io_A_Valid_4_delay_13_15 <= io_A_Valid_4_delay_12_16;
    io_A_Valid_4_delay_14_14 <= io_A_Valid_4_delay_13_15;
    io_A_Valid_4_delay_15_13 <= io_A_Valid_4_delay_14_14;
    io_A_Valid_4_delay_16_12 <= io_A_Valid_4_delay_15_13;
    io_A_Valid_4_delay_17_11 <= io_A_Valid_4_delay_16_12;
    io_A_Valid_4_delay_18_10 <= io_A_Valid_4_delay_17_11;
    io_A_Valid_4_delay_19_9 <= io_A_Valid_4_delay_18_10;
    io_A_Valid_4_delay_20_8 <= io_A_Valid_4_delay_19_9;
    io_A_Valid_4_delay_21_7 <= io_A_Valid_4_delay_20_8;
    io_A_Valid_4_delay_22_6 <= io_A_Valid_4_delay_21_7;
    io_A_Valid_4_delay_23_5 <= io_A_Valid_4_delay_22_6;
    io_A_Valid_4_delay_24_4 <= io_A_Valid_4_delay_23_5;
    io_A_Valid_4_delay_25_3 <= io_A_Valid_4_delay_24_4;
    io_A_Valid_4_delay_26_2 <= io_A_Valid_4_delay_25_3;
    io_A_Valid_4_delay_27_1 <= io_A_Valid_4_delay_26_2;
    io_A_Valid_4_delay_28 <= io_A_Valid_4_delay_27_1;
    io_B_Valid_28_delay_1_3 <= io_B_Valid_28;
    io_B_Valid_28_delay_2_2 <= io_B_Valid_28_delay_1_3;
    io_B_Valid_28_delay_3_1 <= io_B_Valid_28_delay_2_2;
    io_B_Valid_28_delay_4 <= io_B_Valid_28_delay_3_1;
    io_A_Valid_4_delay_1_28 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_27 <= io_A_Valid_4_delay_1_28;
    io_A_Valid_4_delay_3_26 <= io_A_Valid_4_delay_2_27;
    io_A_Valid_4_delay_4_25 <= io_A_Valid_4_delay_3_26;
    io_A_Valid_4_delay_5_24 <= io_A_Valid_4_delay_4_25;
    io_A_Valid_4_delay_6_23 <= io_A_Valid_4_delay_5_24;
    io_A_Valid_4_delay_7_22 <= io_A_Valid_4_delay_6_23;
    io_A_Valid_4_delay_8_21 <= io_A_Valid_4_delay_7_22;
    io_A_Valid_4_delay_9_20 <= io_A_Valid_4_delay_8_21;
    io_A_Valid_4_delay_10_19 <= io_A_Valid_4_delay_9_20;
    io_A_Valid_4_delay_11_18 <= io_A_Valid_4_delay_10_19;
    io_A_Valid_4_delay_12_17 <= io_A_Valid_4_delay_11_18;
    io_A_Valid_4_delay_13_16 <= io_A_Valid_4_delay_12_17;
    io_A_Valid_4_delay_14_15 <= io_A_Valid_4_delay_13_16;
    io_A_Valid_4_delay_15_14 <= io_A_Valid_4_delay_14_15;
    io_A_Valid_4_delay_16_13 <= io_A_Valid_4_delay_15_14;
    io_A_Valid_4_delay_17_12 <= io_A_Valid_4_delay_16_13;
    io_A_Valid_4_delay_18_11 <= io_A_Valid_4_delay_17_12;
    io_A_Valid_4_delay_19_10 <= io_A_Valid_4_delay_18_11;
    io_A_Valid_4_delay_20_9 <= io_A_Valid_4_delay_19_10;
    io_A_Valid_4_delay_21_8 <= io_A_Valid_4_delay_20_9;
    io_A_Valid_4_delay_22_7 <= io_A_Valid_4_delay_21_8;
    io_A_Valid_4_delay_23_6 <= io_A_Valid_4_delay_22_7;
    io_A_Valid_4_delay_24_5 <= io_A_Valid_4_delay_23_6;
    io_A_Valid_4_delay_25_4 <= io_A_Valid_4_delay_24_5;
    io_A_Valid_4_delay_26_3 <= io_A_Valid_4_delay_25_4;
    io_A_Valid_4_delay_27_2 <= io_A_Valid_4_delay_26_3;
    io_A_Valid_4_delay_28_1 <= io_A_Valid_4_delay_27_2;
    io_A_Valid_4_delay_29 <= io_A_Valid_4_delay_28_1;
    io_B_Valid_29_delay_1_3 <= io_B_Valid_29;
    io_B_Valid_29_delay_2_2 <= io_B_Valid_29_delay_1_3;
    io_B_Valid_29_delay_3_1 <= io_B_Valid_29_delay_2_2;
    io_B_Valid_29_delay_4 <= io_B_Valid_29_delay_3_1;
    io_A_Valid_4_delay_1_29 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_28 <= io_A_Valid_4_delay_1_29;
    io_A_Valid_4_delay_3_27 <= io_A_Valid_4_delay_2_28;
    io_A_Valid_4_delay_4_26 <= io_A_Valid_4_delay_3_27;
    io_A_Valid_4_delay_5_25 <= io_A_Valid_4_delay_4_26;
    io_A_Valid_4_delay_6_24 <= io_A_Valid_4_delay_5_25;
    io_A_Valid_4_delay_7_23 <= io_A_Valid_4_delay_6_24;
    io_A_Valid_4_delay_8_22 <= io_A_Valid_4_delay_7_23;
    io_A_Valid_4_delay_9_21 <= io_A_Valid_4_delay_8_22;
    io_A_Valid_4_delay_10_20 <= io_A_Valid_4_delay_9_21;
    io_A_Valid_4_delay_11_19 <= io_A_Valid_4_delay_10_20;
    io_A_Valid_4_delay_12_18 <= io_A_Valid_4_delay_11_19;
    io_A_Valid_4_delay_13_17 <= io_A_Valid_4_delay_12_18;
    io_A_Valid_4_delay_14_16 <= io_A_Valid_4_delay_13_17;
    io_A_Valid_4_delay_15_15 <= io_A_Valid_4_delay_14_16;
    io_A_Valid_4_delay_16_14 <= io_A_Valid_4_delay_15_15;
    io_A_Valid_4_delay_17_13 <= io_A_Valid_4_delay_16_14;
    io_A_Valid_4_delay_18_12 <= io_A_Valid_4_delay_17_13;
    io_A_Valid_4_delay_19_11 <= io_A_Valid_4_delay_18_12;
    io_A_Valid_4_delay_20_10 <= io_A_Valid_4_delay_19_11;
    io_A_Valid_4_delay_21_9 <= io_A_Valid_4_delay_20_10;
    io_A_Valid_4_delay_22_8 <= io_A_Valid_4_delay_21_9;
    io_A_Valid_4_delay_23_7 <= io_A_Valid_4_delay_22_8;
    io_A_Valid_4_delay_24_6 <= io_A_Valid_4_delay_23_7;
    io_A_Valid_4_delay_25_5 <= io_A_Valid_4_delay_24_6;
    io_A_Valid_4_delay_26_4 <= io_A_Valid_4_delay_25_5;
    io_A_Valid_4_delay_27_3 <= io_A_Valid_4_delay_26_4;
    io_A_Valid_4_delay_28_2 <= io_A_Valid_4_delay_27_3;
    io_A_Valid_4_delay_29_1 <= io_A_Valid_4_delay_28_2;
    io_A_Valid_4_delay_30 <= io_A_Valid_4_delay_29_1;
    io_B_Valid_30_delay_1_3 <= io_B_Valid_30;
    io_B_Valid_30_delay_2_2 <= io_B_Valid_30_delay_1_3;
    io_B_Valid_30_delay_3_1 <= io_B_Valid_30_delay_2_2;
    io_B_Valid_30_delay_4 <= io_B_Valid_30_delay_3_1;
    io_A_Valid_4_delay_1_30 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_29 <= io_A_Valid_4_delay_1_30;
    io_A_Valid_4_delay_3_28 <= io_A_Valid_4_delay_2_29;
    io_A_Valid_4_delay_4_27 <= io_A_Valid_4_delay_3_28;
    io_A_Valid_4_delay_5_26 <= io_A_Valid_4_delay_4_27;
    io_A_Valid_4_delay_6_25 <= io_A_Valid_4_delay_5_26;
    io_A_Valid_4_delay_7_24 <= io_A_Valid_4_delay_6_25;
    io_A_Valid_4_delay_8_23 <= io_A_Valid_4_delay_7_24;
    io_A_Valid_4_delay_9_22 <= io_A_Valid_4_delay_8_23;
    io_A_Valid_4_delay_10_21 <= io_A_Valid_4_delay_9_22;
    io_A_Valid_4_delay_11_20 <= io_A_Valid_4_delay_10_21;
    io_A_Valid_4_delay_12_19 <= io_A_Valid_4_delay_11_20;
    io_A_Valid_4_delay_13_18 <= io_A_Valid_4_delay_12_19;
    io_A_Valid_4_delay_14_17 <= io_A_Valid_4_delay_13_18;
    io_A_Valid_4_delay_15_16 <= io_A_Valid_4_delay_14_17;
    io_A_Valid_4_delay_16_15 <= io_A_Valid_4_delay_15_16;
    io_A_Valid_4_delay_17_14 <= io_A_Valid_4_delay_16_15;
    io_A_Valid_4_delay_18_13 <= io_A_Valid_4_delay_17_14;
    io_A_Valid_4_delay_19_12 <= io_A_Valid_4_delay_18_13;
    io_A_Valid_4_delay_20_11 <= io_A_Valid_4_delay_19_12;
    io_A_Valid_4_delay_21_10 <= io_A_Valid_4_delay_20_11;
    io_A_Valid_4_delay_22_9 <= io_A_Valid_4_delay_21_10;
    io_A_Valid_4_delay_23_8 <= io_A_Valid_4_delay_22_9;
    io_A_Valid_4_delay_24_7 <= io_A_Valid_4_delay_23_8;
    io_A_Valid_4_delay_25_6 <= io_A_Valid_4_delay_24_7;
    io_A_Valid_4_delay_26_5 <= io_A_Valid_4_delay_25_6;
    io_A_Valid_4_delay_27_4 <= io_A_Valid_4_delay_26_5;
    io_A_Valid_4_delay_28_3 <= io_A_Valid_4_delay_27_4;
    io_A_Valid_4_delay_29_2 <= io_A_Valid_4_delay_28_3;
    io_A_Valid_4_delay_30_1 <= io_A_Valid_4_delay_29_2;
    io_A_Valid_4_delay_31 <= io_A_Valid_4_delay_30_1;
    io_B_Valid_31_delay_1_3 <= io_B_Valid_31;
    io_B_Valid_31_delay_2_2 <= io_B_Valid_31_delay_1_3;
    io_B_Valid_31_delay_3_1 <= io_B_Valid_31_delay_2_2;
    io_B_Valid_31_delay_4 <= io_B_Valid_31_delay_3_1;
    io_A_Valid_4_delay_1_31 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_30 <= io_A_Valid_4_delay_1_31;
    io_A_Valid_4_delay_3_29 <= io_A_Valid_4_delay_2_30;
    io_A_Valid_4_delay_4_28 <= io_A_Valid_4_delay_3_29;
    io_A_Valid_4_delay_5_27 <= io_A_Valid_4_delay_4_28;
    io_A_Valid_4_delay_6_26 <= io_A_Valid_4_delay_5_27;
    io_A_Valid_4_delay_7_25 <= io_A_Valid_4_delay_6_26;
    io_A_Valid_4_delay_8_24 <= io_A_Valid_4_delay_7_25;
    io_A_Valid_4_delay_9_23 <= io_A_Valid_4_delay_8_24;
    io_A_Valid_4_delay_10_22 <= io_A_Valid_4_delay_9_23;
    io_A_Valid_4_delay_11_21 <= io_A_Valid_4_delay_10_22;
    io_A_Valid_4_delay_12_20 <= io_A_Valid_4_delay_11_21;
    io_A_Valid_4_delay_13_19 <= io_A_Valid_4_delay_12_20;
    io_A_Valid_4_delay_14_18 <= io_A_Valid_4_delay_13_19;
    io_A_Valid_4_delay_15_17 <= io_A_Valid_4_delay_14_18;
    io_A_Valid_4_delay_16_16 <= io_A_Valid_4_delay_15_17;
    io_A_Valid_4_delay_17_15 <= io_A_Valid_4_delay_16_16;
    io_A_Valid_4_delay_18_14 <= io_A_Valid_4_delay_17_15;
    io_A_Valid_4_delay_19_13 <= io_A_Valid_4_delay_18_14;
    io_A_Valid_4_delay_20_12 <= io_A_Valid_4_delay_19_13;
    io_A_Valid_4_delay_21_11 <= io_A_Valid_4_delay_20_12;
    io_A_Valid_4_delay_22_10 <= io_A_Valid_4_delay_21_11;
    io_A_Valid_4_delay_23_9 <= io_A_Valid_4_delay_22_10;
    io_A_Valid_4_delay_24_8 <= io_A_Valid_4_delay_23_9;
    io_A_Valid_4_delay_25_7 <= io_A_Valid_4_delay_24_8;
    io_A_Valid_4_delay_26_6 <= io_A_Valid_4_delay_25_7;
    io_A_Valid_4_delay_27_5 <= io_A_Valid_4_delay_26_6;
    io_A_Valid_4_delay_28_4 <= io_A_Valid_4_delay_27_5;
    io_A_Valid_4_delay_29_3 <= io_A_Valid_4_delay_28_4;
    io_A_Valid_4_delay_30_2 <= io_A_Valid_4_delay_29_3;
    io_A_Valid_4_delay_31_1 <= io_A_Valid_4_delay_30_2;
    io_A_Valid_4_delay_32 <= io_A_Valid_4_delay_31_1;
    io_B_Valid_32_delay_1_3 <= io_B_Valid_32;
    io_B_Valid_32_delay_2_2 <= io_B_Valid_32_delay_1_3;
    io_B_Valid_32_delay_3_1 <= io_B_Valid_32_delay_2_2;
    io_B_Valid_32_delay_4 <= io_B_Valid_32_delay_3_1;
    io_A_Valid_4_delay_1_32 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_31 <= io_A_Valid_4_delay_1_32;
    io_A_Valid_4_delay_3_30 <= io_A_Valid_4_delay_2_31;
    io_A_Valid_4_delay_4_29 <= io_A_Valid_4_delay_3_30;
    io_A_Valid_4_delay_5_28 <= io_A_Valid_4_delay_4_29;
    io_A_Valid_4_delay_6_27 <= io_A_Valid_4_delay_5_28;
    io_A_Valid_4_delay_7_26 <= io_A_Valid_4_delay_6_27;
    io_A_Valid_4_delay_8_25 <= io_A_Valid_4_delay_7_26;
    io_A_Valid_4_delay_9_24 <= io_A_Valid_4_delay_8_25;
    io_A_Valid_4_delay_10_23 <= io_A_Valid_4_delay_9_24;
    io_A_Valid_4_delay_11_22 <= io_A_Valid_4_delay_10_23;
    io_A_Valid_4_delay_12_21 <= io_A_Valid_4_delay_11_22;
    io_A_Valid_4_delay_13_20 <= io_A_Valid_4_delay_12_21;
    io_A_Valid_4_delay_14_19 <= io_A_Valid_4_delay_13_20;
    io_A_Valid_4_delay_15_18 <= io_A_Valid_4_delay_14_19;
    io_A_Valid_4_delay_16_17 <= io_A_Valid_4_delay_15_18;
    io_A_Valid_4_delay_17_16 <= io_A_Valid_4_delay_16_17;
    io_A_Valid_4_delay_18_15 <= io_A_Valid_4_delay_17_16;
    io_A_Valid_4_delay_19_14 <= io_A_Valid_4_delay_18_15;
    io_A_Valid_4_delay_20_13 <= io_A_Valid_4_delay_19_14;
    io_A_Valid_4_delay_21_12 <= io_A_Valid_4_delay_20_13;
    io_A_Valid_4_delay_22_11 <= io_A_Valid_4_delay_21_12;
    io_A_Valid_4_delay_23_10 <= io_A_Valid_4_delay_22_11;
    io_A_Valid_4_delay_24_9 <= io_A_Valid_4_delay_23_10;
    io_A_Valid_4_delay_25_8 <= io_A_Valid_4_delay_24_9;
    io_A_Valid_4_delay_26_7 <= io_A_Valid_4_delay_25_8;
    io_A_Valid_4_delay_27_6 <= io_A_Valid_4_delay_26_7;
    io_A_Valid_4_delay_28_5 <= io_A_Valid_4_delay_27_6;
    io_A_Valid_4_delay_29_4 <= io_A_Valid_4_delay_28_5;
    io_A_Valid_4_delay_30_3 <= io_A_Valid_4_delay_29_4;
    io_A_Valid_4_delay_31_2 <= io_A_Valid_4_delay_30_3;
    io_A_Valid_4_delay_32_1 <= io_A_Valid_4_delay_31_2;
    io_A_Valid_4_delay_33 <= io_A_Valid_4_delay_32_1;
    io_B_Valid_33_delay_1_3 <= io_B_Valid_33;
    io_B_Valid_33_delay_2_2 <= io_B_Valid_33_delay_1_3;
    io_B_Valid_33_delay_3_1 <= io_B_Valid_33_delay_2_2;
    io_B_Valid_33_delay_4 <= io_B_Valid_33_delay_3_1;
    io_A_Valid_4_delay_1_33 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_32 <= io_A_Valid_4_delay_1_33;
    io_A_Valid_4_delay_3_31 <= io_A_Valid_4_delay_2_32;
    io_A_Valid_4_delay_4_30 <= io_A_Valid_4_delay_3_31;
    io_A_Valid_4_delay_5_29 <= io_A_Valid_4_delay_4_30;
    io_A_Valid_4_delay_6_28 <= io_A_Valid_4_delay_5_29;
    io_A_Valid_4_delay_7_27 <= io_A_Valid_4_delay_6_28;
    io_A_Valid_4_delay_8_26 <= io_A_Valid_4_delay_7_27;
    io_A_Valid_4_delay_9_25 <= io_A_Valid_4_delay_8_26;
    io_A_Valid_4_delay_10_24 <= io_A_Valid_4_delay_9_25;
    io_A_Valid_4_delay_11_23 <= io_A_Valid_4_delay_10_24;
    io_A_Valid_4_delay_12_22 <= io_A_Valid_4_delay_11_23;
    io_A_Valid_4_delay_13_21 <= io_A_Valid_4_delay_12_22;
    io_A_Valid_4_delay_14_20 <= io_A_Valid_4_delay_13_21;
    io_A_Valid_4_delay_15_19 <= io_A_Valid_4_delay_14_20;
    io_A_Valid_4_delay_16_18 <= io_A_Valid_4_delay_15_19;
    io_A_Valid_4_delay_17_17 <= io_A_Valid_4_delay_16_18;
    io_A_Valid_4_delay_18_16 <= io_A_Valid_4_delay_17_17;
    io_A_Valid_4_delay_19_15 <= io_A_Valid_4_delay_18_16;
    io_A_Valid_4_delay_20_14 <= io_A_Valid_4_delay_19_15;
    io_A_Valid_4_delay_21_13 <= io_A_Valid_4_delay_20_14;
    io_A_Valid_4_delay_22_12 <= io_A_Valid_4_delay_21_13;
    io_A_Valid_4_delay_23_11 <= io_A_Valid_4_delay_22_12;
    io_A_Valid_4_delay_24_10 <= io_A_Valid_4_delay_23_11;
    io_A_Valid_4_delay_25_9 <= io_A_Valid_4_delay_24_10;
    io_A_Valid_4_delay_26_8 <= io_A_Valid_4_delay_25_9;
    io_A_Valid_4_delay_27_7 <= io_A_Valid_4_delay_26_8;
    io_A_Valid_4_delay_28_6 <= io_A_Valid_4_delay_27_7;
    io_A_Valid_4_delay_29_5 <= io_A_Valid_4_delay_28_6;
    io_A_Valid_4_delay_30_4 <= io_A_Valid_4_delay_29_5;
    io_A_Valid_4_delay_31_3 <= io_A_Valid_4_delay_30_4;
    io_A_Valid_4_delay_32_2 <= io_A_Valid_4_delay_31_3;
    io_A_Valid_4_delay_33_1 <= io_A_Valid_4_delay_32_2;
    io_A_Valid_4_delay_34 <= io_A_Valid_4_delay_33_1;
    io_B_Valid_34_delay_1_3 <= io_B_Valid_34;
    io_B_Valid_34_delay_2_2 <= io_B_Valid_34_delay_1_3;
    io_B_Valid_34_delay_3_1 <= io_B_Valid_34_delay_2_2;
    io_B_Valid_34_delay_4 <= io_B_Valid_34_delay_3_1;
    io_A_Valid_4_delay_1_34 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_33 <= io_A_Valid_4_delay_1_34;
    io_A_Valid_4_delay_3_32 <= io_A_Valid_4_delay_2_33;
    io_A_Valid_4_delay_4_31 <= io_A_Valid_4_delay_3_32;
    io_A_Valid_4_delay_5_30 <= io_A_Valid_4_delay_4_31;
    io_A_Valid_4_delay_6_29 <= io_A_Valid_4_delay_5_30;
    io_A_Valid_4_delay_7_28 <= io_A_Valid_4_delay_6_29;
    io_A_Valid_4_delay_8_27 <= io_A_Valid_4_delay_7_28;
    io_A_Valid_4_delay_9_26 <= io_A_Valid_4_delay_8_27;
    io_A_Valid_4_delay_10_25 <= io_A_Valid_4_delay_9_26;
    io_A_Valid_4_delay_11_24 <= io_A_Valid_4_delay_10_25;
    io_A_Valid_4_delay_12_23 <= io_A_Valid_4_delay_11_24;
    io_A_Valid_4_delay_13_22 <= io_A_Valid_4_delay_12_23;
    io_A_Valid_4_delay_14_21 <= io_A_Valid_4_delay_13_22;
    io_A_Valid_4_delay_15_20 <= io_A_Valid_4_delay_14_21;
    io_A_Valid_4_delay_16_19 <= io_A_Valid_4_delay_15_20;
    io_A_Valid_4_delay_17_18 <= io_A_Valid_4_delay_16_19;
    io_A_Valid_4_delay_18_17 <= io_A_Valid_4_delay_17_18;
    io_A_Valid_4_delay_19_16 <= io_A_Valid_4_delay_18_17;
    io_A_Valid_4_delay_20_15 <= io_A_Valid_4_delay_19_16;
    io_A_Valid_4_delay_21_14 <= io_A_Valid_4_delay_20_15;
    io_A_Valid_4_delay_22_13 <= io_A_Valid_4_delay_21_14;
    io_A_Valid_4_delay_23_12 <= io_A_Valid_4_delay_22_13;
    io_A_Valid_4_delay_24_11 <= io_A_Valid_4_delay_23_12;
    io_A_Valid_4_delay_25_10 <= io_A_Valid_4_delay_24_11;
    io_A_Valid_4_delay_26_9 <= io_A_Valid_4_delay_25_10;
    io_A_Valid_4_delay_27_8 <= io_A_Valid_4_delay_26_9;
    io_A_Valid_4_delay_28_7 <= io_A_Valid_4_delay_27_8;
    io_A_Valid_4_delay_29_6 <= io_A_Valid_4_delay_28_7;
    io_A_Valid_4_delay_30_5 <= io_A_Valid_4_delay_29_6;
    io_A_Valid_4_delay_31_4 <= io_A_Valid_4_delay_30_5;
    io_A_Valid_4_delay_32_3 <= io_A_Valid_4_delay_31_4;
    io_A_Valid_4_delay_33_2 <= io_A_Valid_4_delay_32_3;
    io_A_Valid_4_delay_34_1 <= io_A_Valid_4_delay_33_2;
    io_A_Valid_4_delay_35 <= io_A_Valid_4_delay_34_1;
    io_B_Valid_35_delay_1_3 <= io_B_Valid_35;
    io_B_Valid_35_delay_2_2 <= io_B_Valid_35_delay_1_3;
    io_B_Valid_35_delay_3_1 <= io_B_Valid_35_delay_2_2;
    io_B_Valid_35_delay_4 <= io_B_Valid_35_delay_3_1;
    io_A_Valid_4_delay_1_35 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_34 <= io_A_Valid_4_delay_1_35;
    io_A_Valid_4_delay_3_33 <= io_A_Valid_4_delay_2_34;
    io_A_Valid_4_delay_4_32 <= io_A_Valid_4_delay_3_33;
    io_A_Valid_4_delay_5_31 <= io_A_Valid_4_delay_4_32;
    io_A_Valid_4_delay_6_30 <= io_A_Valid_4_delay_5_31;
    io_A_Valid_4_delay_7_29 <= io_A_Valid_4_delay_6_30;
    io_A_Valid_4_delay_8_28 <= io_A_Valid_4_delay_7_29;
    io_A_Valid_4_delay_9_27 <= io_A_Valid_4_delay_8_28;
    io_A_Valid_4_delay_10_26 <= io_A_Valid_4_delay_9_27;
    io_A_Valid_4_delay_11_25 <= io_A_Valid_4_delay_10_26;
    io_A_Valid_4_delay_12_24 <= io_A_Valid_4_delay_11_25;
    io_A_Valid_4_delay_13_23 <= io_A_Valid_4_delay_12_24;
    io_A_Valid_4_delay_14_22 <= io_A_Valid_4_delay_13_23;
    io_A_Valid_4_delay_15_21 <= io_A_Valid_4_delay_14_22;
    io_A_Valid_4_delay_16_20 <= io_A_Valid_4_delay_15_21;
    io_A_Valid_4_delay_17_19 <= io_A_Valid_4_delay_16_20;
    io_A_Valid_4_delay_18_18 <= io_A_Valid_4_delay_17_19;
    io_A_Valid_4_delay_19_17 <= io_A_Valid_4_delay_18_18;
    io_A_Valid_4_delay_20_16 <= io_A_Valid_4_delay_19_17;
    io_A_Valid_4_delay_21_15 <= io_A_Valid_4_delay_20_16;
    io_A_Valid_4_delay_22_14 <= io_A_Valid_4_delay_21_15;
    io_A_Valid_4_delay_23_13 <= io_A_Valid_4_delay_22_14;
    io_A_Valid_4_delay_24_12 <= io_A_Valid_4_delay_23_13;
    io_A_Valid_4_delay_25_11 <= io_A_Valid_4_delay_24_12;
    io_A_Valid_4_delay_26_10 <= io_A_Valid_4_delay_25_11;
    io_A_Valid_4_delay_27_9 <= io_A_Valid_4_delay_26_10;
    io_A_Valid_4_delay_28_8 <= io_A_Valid_4_delay_27_9;
    io_A_Valid_4_delay_29_7 <= io_A_Valid_4_delay_28_8;
    io_A_Valid_4_delay_30_6 <= io_A_Valid_4_delay_29_7;
    io_A_Valid_4_delay_31_5 <= io_A_Valid_4_delay_30_6;
    io_A_Valid_4_delay_32_4 <= io_A_Valid_4_delay_31_5;
    io_A_Valid_4_delay_33_3 <= io_A_Valid_4_delay_32_4;
    io_A_Valid_4_delay_34_2 <= io_A_Valid_4_delay_33_3;
    io_A_Valid_4_delay_35_1 <= io_A_Valid_4_delay_34_2;
    io_A_Valid_4_delay_36 <= io_A_Valid_4_delay_35_1;
    io_B_Valid_36_delay_1_3 <= io_B_Valid_36;
    io_B_Valid_36_delay_2_2 <= io_B_Valid_36_delay_1_3;
    io_B_Valid_36_delay_3_1 <= io_B_Valid_36_delay_2_2;
    io_B_Valid_36_delay_4 <= io_B_Valid_36_delay_3_1;
    io_A_Valid_4_delay_1_36 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_35 <= io_A_Valid_4_delay_1_36;
    io_A_Valid_4_delay_3_34 <= io_A_Valid_4_delay_2_35;
    io_A_Valid_4_delay_4_33 <= io_A_Valid_4_delay_3_34;
    io_A_Valid_4_delay_5_32 <= io_A_Valid_4_delay_4_33;
    io_A_Valid_4_delay_6_31 <= io_A_Valid_4_delay_5_32;
    io_A_Valid_4_delay_7_30 <= io_A_Valid_4_delay_6_31;
    io_A_Valid_4_delay_8_29 <= io_A_Valid_4_delay_7_30;
    io_A_Valid_4_delay_9_28 <= io_A_Valid_4_delay_8_29;
    io_A_Valid_4_delay_10_27 <= io_A_Valid_4_delay_9_28;
    io_A_Valid_4_delay_11_26 <= io_A_Valid_4_delay_10_27;
    io_A_Valid_4_delay_12_25 <= io_A_Valid_4_delay_11_26;
    io_A_Valid_4_delay_13_24 <= io_A_Valid_4_delay_12_25;
    io_A_Valid_4_delay_14_23 <= io_A_Valid_4_delay_13_24;
    io_A_Valid_4_delay_15_22 <= io_A_Valid_4_delay_14_23;
    io_A_Valid_4_delay_16_21 <= io_A_Valid_4_delay_15_22;
    io_A_Valid_4_delay_17_20 <= io_A_Valid_4_delay_16_21;
    io_A_Valid_4_delay_18_19 <= io_A_Valid_4_delay_17_20;
    io_A_Valid_4_delay_19_18 <= io_A_Valid_4_delay_18_19;
    io_A_Valid_4_delay_20_17 <= io_A_Valid_4_delay_19_18;
    io_A_Valid_4_delay_21_16 <= io_A_Valid_4_delay_20_17;
    io_A_Valid_4_delay_22_15 <= io_A_Valid_4_delay_21_16;
    io_A_Valid_4_delay_23_14 <= io_A_Valid_4_delay_22_15;
    io_A_Valid_4_delay_24_13 <= io_A_Valid_4_delay_23_14;
    io_A_Valid_4_delay_25_12 <= io_A_Valid_4_delay_24_13;
    io_A_Valid_4_delay_26_11 <= io_A_Valid_4_delay_25_12;
    io_A_Valid_4_delay_27_10 <= io_A_Valid_4_delay_26_11;
    io_A_Valid_4_delay_28_9 <= io_A_Valid_4_delay_27_10;
    io_A_Valid_4_delay_29_8 <= io_A_Valid_4_delay_28_9;
    io_A_Valid_4_delay_30_7 <= io_A_Valid_4_delay_29_8;
    io_A_Valid_4_delay_31_6 <= io_A_Valid_4_delay_30_7;
    io_A_Valid_4_delay_32_5 <= io_A_Valid_4_delay_31_6;
    io_A_Valid_4_delay_33_4 <= io_A_Valid_4_delay_32_5;
    io_A_Valid_4_delay_34_3 <= io_A_Valid_4_delay_33_4;
    io_A_Valid_4_delay_35_2 <= io_A_Valid_4_delay_34_3;
    io_A_Valid_4_delay_36_1 <= io_A_Valid_4_delay_35_2;
    io_A_Valid_4_delay_37 <= io_A_Valid_4_delay_36_1;
    io_B_Valid_37_delay_1_3 <= io_B_Valid_37;
    io_B_Valid_37_delay_2_2 <= io_B_Valid_37_delay_1_3;
    io_B_Valid_37_delay_3_1 <= io_B_Valid_37_delay_2_2;
    io_B_Valid_37_delay_4 <= io_B_Valid_37_delay_3_1;
    io_A_Valid_4_delay_1_37 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_36 <= io_A_Valid_4_delay_1_37;
    io_A_Valid_4_delay_3_35 <= io_A_Valid_4_delay_2_36;
    io_A_Valid_4_delay_4_34 <= io_A_Valid_4_delay_3_35;
    io_A_Valid_4_delay_5_33 <= io_A_Valid_4_delay_4_34;
    io_A_Valid_4_delay_6_32 <= io_A_Valid_4_delay_5_33;
    io_A_Valid_4_delay_7_31 <= io_A_Valid_4_delay_6_32;
    io_A_Valid_4_delay_8_30 <= io_A_Valid_4_delay_7_31;
    io_A_Valid_4_delay_9_29 <= io_A_Valid_4_delay_8_30;
    io_A_Valid_4_delay_10_28 <= io_A_Valid_4_delay_9_29;
    io_A_Valid_4_delay_11_27 <= io_A_Valid_4_delay_10_28;
    io_A_Valid_4_delay_12_26 <= io_A_Valid_4_delay_11_27;
    io_A_Valid_4_delay_13_25 <= io_A_Valid_4_delay_12_26;
    io_A_Valid_4_delay_14_24 <= io_A_Valid_4_delay_13_25;
    io_A_Valid_4_delay_15_23 <= io_A_Valid_4_delay_14_24;
    io_A_Valid_4_delay_16_22 <= io_A_Valid_4_delay_15_23;
    io_A_Valid_4_delay_17_21 <= io_A_Valid_4_delay_16_22;
    io_A_Valid_4_delay_18_20 <= io_A_Valid_4_delay_17_21;
    io_A_Valid_4_delay_19_19 <= io_A_Valid_4_delay_18_20;
    io_A_Valid_4_delay_20_18 <= io_A_Valid_4_delay_19_19;
    io_A_Valid_4_delay_21_17 <= io_A_Valid_4_delay_20_18;
    io_A_Valid_4_delay_22_16 <= io_A_Valid_4_delay_21_17;
    io_A_Valid_4_delay_23_15 <= io_A_Valid_4_delay_22_16;
    io_A_Valid_4_delay_24_14 <= io_A_Valid_4_delay_23_15;
    io_A_Valid_4_delay_25_13 <= io_A_Valid_4_delay_24_14;
    io_A_Valid_4_delay_26_12 <= io_A_Valid_4_delay_25_13;
    io_A_Valid_4_delay_27_11 <= io_A_Valid_4_delay_26_12;
    io_A_Valid_4_delay_28_10 <= io_A_Valid_4_delay_27_11;
    io_A_Valid_4_delay_29_9 <= io_A_Valid_4_delay_28_10;
    io_A_Valid_4_delay_30_8 <= io_A_Valid_4_delay_29_9;
    io_A_Valid_4_delay_31_7 <= io_A_Valid_4_delay_30_8;
    io_A_Valid_4_delay_32_6 <= io_A_Valid_4_delay_31_7;
    io_A_Valid_4_delay_33_5 <= io_A_Valid_4_delay_32_6;
    io_A_Valid_4_delay_34_4 <= io_A_Valid_4_delay_33_5;
    io_A_Valid_4_delay_35_3 <= io_A_Valid_4_delay_34_4;
    io_A_Valid_4_delay_36_2 <= io_A_Valid_4_delay_35_3;
    io_A_Valid_4_delay_37_1 <= io_A_Valid_4_delay_36_2;
    io_A_Valid_4_delay_38 <= io_A_Valid_4_delay_37_1;
    io_B_Valid_38_delay_1_3 <= io_B_Valid_38;
    io_B_Valid_38_delay_2_2 <= io_B_Valid_38_delay_1_3;
    io_B_Valid_38_delay_3_1 <= io_B_Valid_38_delay_2_2;
    io_B_Valid_38_delay_4 <= io_B_Valid_38_delay_3_1;
    io_A_Valid_4_delay_1_38 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_37 <= io_A_Valid_4_delay_1_38;
    io_A_Valid_4_delay_3_36 <= io_A_Valid_4_delay_2_37;
    io_A_Valid_4_delay_4_35 <= io_A_Valid_4_delay_3_36;
    io_A_Valid_4_delay_5_34 <= io_A_Valid_4_delay_4_35;
    io_A_Valid_4_delay_6_33 <= io_A_Valid_4_delay_5_34;
    io_A_Valid_4_delay_7_32 <= io_A_Valid_4_delay_6_33;
    io_A_Valid_4_delay_8_31 <= io_A_Valid_4_delay_7_32;
    io_A_Valid_4_delay_9_30 <= io_A_Valid_4_delay_8_31;
    io_A_Valid_4_delay_10_29 <= io_A_Valid_4_delay_9_30;
    io_A_Valid_4_delay_11_28 <= io_A_Valid_4_delay_10_29;
    io_A_Valid_4_delay_12_27 <= io_A_Valid_4_delay_11_28;
    io_A_Valid_4_delay_13_26 <= io_A_Valid_4_delay_12_27;
    io_A_Valid_4_delay_14_25 <= io_A_Valid_4_delay_13_26;
    io_A_Valid_4_delay_15_24 <= io_A_Valid_4_delay_14_25;
    io_A_Valid_4_delay_16_23 <= io_A_Valid_4_delay_15_24;
    io_A_Valid_4_delay_17_22 <= io_A_Valid_4_delay_16_23;
    io_A_Valid_4_delay_18_21 <= io_A_Valid_4_delay_17_22;
    io_A_Valid_4_delay_19_20 <= io_A_Valid_4_delay_18_21;
    io_A_Valid_4_delay_20_19 <= io_A_Valid_4_delay_19_20;
    io_A_Valid_4_delay_21_18 <= io_A_Valid_4_delay_20_19;
    io_A_Valid_4_delay_22_17 <= io_A_Valid_4_delay_21_18;
    io_A_Valid_4_delay_23_16 <= io_A_Valid_4_delay_22_17;
    io_A_Valid_4_delay_24_15 <= io_A_Valid_4_delay_23_16;
    io_A_Valid_4_delay_25_14 <= io_A_Valid_4_delay_24_15;
    io_A_Valid_4_delay_26_13 <= io_A_Valid_4_delay_25_14;
    io_A_Valid_4_delay_27_12 <= io_A_Valid_4_delay_26_13;
    io_A_Valid_4_delay_28_11 <= io_A_Valid_4_delay_27_12;
    io_A_Valid_4_delay_29_10 <= io_A_Valid_4_delay_28_11;
    io_A_Valid_4_delay_30_9 <= io_A_Valid_4_delay_29_10;
    io_A_Valid_4_delay_31_8 <= io_A_Valid_4_delay_30_9;
    io_A_Valid_4_delay_32_7 <= io_A_Valid_4_delay_31_8;
    io_A_Valid_4_delay_33_6 <= io_A_Valid_4_delay_32_7;
    io_A_Valid_4_delay_34_5 <= io_A_Valid_4_delay_33_6;
    io_A_Valid_4_delay_35_4 <= io_A_Valid_4_delay_34_5;
    io_A_Valid_4_delay_36_3 <= io_A_Valid_4_delay_35_4;
    io_A_Valid_4_delay_37_2 <= io_A_Valid_4_delay_36_3;
    io_A_Valid_4_delay_38_1 <= io_A_Valid_4_delay_37_2;
    io_A_Valid_4_delay_39 <= io_A_Valid_4_delay_38_1;
    io_B_Valid_39_delay_1_3 <= io_B_Valid_39;
    io_B_Valid_39_delay_2_2 <= io_B_Valid_39_delay_1_3;
    io_B_Valid_39_delay_3_1 <= io_B_Valid_39_delay_2_2;
    io_B_Valid_39_delay_4 <= io_B_Valid_39_delay_3_1;
    io_A_Valid_4_delay_1_39 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_38 <= io_A_Valid_4_delay_1_39;
    io_A_Valid_4_delay_3_37 <= io_A_Valid_4_delay_2_38;
    io_A_Valid_4_delay_4_36 <= io_A_Valid_4_delay_3_37;
    io_A_Valid_4_delay_5_35 <= io_A_Valid_4_delay_4_36;
    io_A_Valid_4_delay_6_34 <= io_A_Valid_4_delay_5_35;
    io_A_Valid_4_delay_7_33 <= io_A_Valid_4_delay_6_34;
    io_A_Valid_4_delay_8_32 <= io_A_Valid_4_delay_7_33;
    io_A_Valid_4_delay_9_31 <= io_A_Valid_4_delay_8_32;
    io_A_Valid_4_delay_10_30 <= io_A_Valid_4_delay_9_31;
    io_A_Valid_4_delay_11_29 <= io_A_Valid_4_delay_10_30;
    io_A_Valid_4_delay_12_28 <= io_A_Valid_4_delay_11_29;
    io_A_Valid_4_delay_13_27 <= io_A_Valid_4_delay_12_28;
    io_A_Valid_4_delay_14_26 <= io_A_Valid_4_delay_13_27;
    io_A_Valid_4_delay_15_25 <= io_A_Valid_4_delay_14_26;
    io_A_Valid_4_delay_16_24 <= io_A_Valid_4_delay_15_25;
    io_A_Valid_4_delay_17_23 <= io_A_Valid_4_delay_16_24;
    io_A_Valid_4_delay_18_22 <= io_A_Valid_4_delay_17_23;
    io_A_Valid_4_delay_19_21 <= io_A_Valid_4_delay_18_22;
    io_A_Valid_4_delay_20_20 <= io_A_Valid_4_delay_19_21;
    io_A_Valid_4_delay_21_19 <= io_A_Valid_4_delay_20_20;
    io_A_Valid_4_delay_22_18 <= io_A_Valid_4_delay_21_19;
    io_A_Valid_4_delay_23_17 <= io_A_Valid_4_delay_22_18;
    io_A_Valid_4_delay_24_16 <= io_A_Valid_4_delay_23_17;
    io_A_Valid_4_delay_25_15 <= io_A_Valid_4_delay_24_16;
    io_A_Valid_4_delay_26_14 <= io_A_Valid_4_delay_25_15;
    io_A_Valid_4_delay_27_13 <= io_A_Valid_4_delay_26_14;
    io_A_Valid_4_delay_28_12 <= io_A_Valid_4_delay_27_13;
    io_A_Valid_4_delay_29_11 <= io_A_Valid_4_delay_28_12;
    io_A_Valid_4_delay_30_10 <= io_A_Valid_4_delay_29_11;
    io_A_Valid_4_delay_31_9 <= io_A_Valid_4_delay_30_10;
    io_A_Valid_4_delay_32_8 <= io_A_Valid_4_delay_31_9;
    io_A_Valid_4_delay_33_7 <= io_A_Valid_4_delay_32_8;
    io_A_Valid_4_delay_34_6 <= io_A_Valid_4_delay_33_7;
    io_A_Valid_4_delay_35_5 <= io_A_Valid_4_delay_34_6;
    io_A_Valid_4_delay_36_4 <= io_A_Valid_4_delay_35_5;
    io_A_Valid_4_delay_37_3 <= io_A_Valid_4_delay_36_4;
    io_A_Valid_4_delay_38_2 <= io_A_Valid_4_delay_37_3;
    io_A_Valid_4_delay_39_1 <= io_A_Valid_4_delay_38_2;
    io_A_Valid_4_delay_40 <= io_A_Valid_4_delay_39_1;
    io_B_Valid_40_delay_1_3 <= io_B_Valid_40;
    io_B_Valid_40_delay_2_2 <= io_B_Valid_40_delay_1_3;
    io_B_Valid_40_delay_3_1 <= io_B_Valid_40_delay_2_2;
    io_B_Valid_40_delay_4 <= io_B_Valid_40_delay_3_1;
    io_A_Valid_4_delay_1_40 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_39 <= io_A_Valid_4_delay_1_40;
    io_A_Valid_4_delay_3_38 <= io_A_Valid_4_delay_2_39;
    io_A_Valid_4_delay_4_37 <= io_A_Valid_4_delay_3_38;
    io_A_Valid_4_delay_5_36 <= io_A_Valid_4_delay_4_37;
    io_A_Valid_4_delay_6_35 <= io_A_Valid_4_delay_5_36;
    io_A_Valid_4_delay_7_34 <= io_A_Valid_4_delay_6_35;
    io_A_Valid_4_delay_8_33 <= io_A_Valid_4_delay_7_34;
    io_A_Valid_4_delay_9_32 <= io_A_Valid_4_delay_8_33;
    io_A_Valid_4_delay_10_31 <= io_A_Valid_4_delay_9_32;
    io_A_Valid_4_delay_11_30 <= io_A_Valid_4_delay_10_31;
    io_A_Valid_4_delay_12_29 <= io_A_Valid_4_delay_11_30;
    io_A_Valid_4_delay_13_28 <= io_A_Valid_4_delay_12_29;
    io_A_Valid_4_delay_14_27 <= io_A_Valid_4_delay_13_28;
    io_A_Valid_4_delay_15_26 <= io_A_Valid_4_delay_14_27;
    io_A_Valid_4_delay_16_25 <= io_A_Valid_4_delay_15_26;
    io_A_Valid_4_delay_17_24 <= io_A_Valid_4_delay_16_25;
    io_A_Valid_4_delay_18_23 <= io_A_Valid_4_delay_17_24;
    io_A_Valid_4_delay_19_22 <= io_A_Valid_4_delay_18_23;
    io_A_Valid_4_delay_20_21 <= io_A_Valid_4_delay_19_22;
    io_A_Valid_4_delay_21_20 <= io_A_Valid_4_delay_20_21;
    io_A_Valid_4_delay_22_19 <= io_A_Valid_4_delay_21_20;
    io_A_Valid_4_delay_23_18 <= io_A_Valid_4_delay_22_19;
    io_A_Valid_4_delay_24_17 <= io_A_Valid_4_delay_23_18;
    io_A_Valid_4_delay_25_16 <= io_A_Valid_4_delay_24_17;
    io_A_Valid_4_delay_26_15 <= io_A_Valid_4_delay_25_16;
    io_A_Valid_4_delay_27_14 <= io_A_Valid_4_delay_26_15;
    io_A_Valid_4_delay_28_13 <= io_A_Valid_4_delay_27_14;
    io_A_Valid_4_delay_29_12 <= io_A_Valid_4_delay_28_13;
    io_A_Valid_4_delay_30_11 <= io_A_Valid_4_delay_29_12;
    io_A_Valid_4_delay_31_10 <= io_A_Valid_4_delay_30_11;
    io_A_Valid_4_delay_32_9 <= io_A_Valid_4_delay_31_10;
    io_A_Valid_4_delay_33_8 <= io_A_Valid_4_delay_32_9;
    io_A_Valid_4_delay_34_7 <= io_A_Valid_4_delay_33_8;
    io_A_Valid_4_delay_35_6 <= io_A_Valid_4_delay_34_7;
    io_A_Valid_4_delay_36_5 <= io_A_Valid_4_delay_35_6;
    io_A_Valid_4_delay_37_4 <= io_A_Valid_4_delay_36_5;
    io_A_Valid_4_delay_38_3 <= io_A_Valid_4_delay_37_4;
    io_A_Valid_4_delay_39_2 <= io_A_Valid_4_delay_38_3;
    io_A_Valid_4_delay_40_1 <= io_A_Valid_4_delay_39_2;
    io_A_Valid_4_delay_41 <= io_A_Valid_4_delay_40_1;
    io_B_Valid_41_delay_1_3 <= io_B_Valid_41;
    io_B_Valid_41_delay_2_2 <= io_B_Valid_41_delay_1_3;
    io_B_Valid_41_delay_3_1 <= io_B_Valid_41_delay_2_2;
    io_B_Valid_41_delay_4 <= io_B_Valid_41_delay_3_1;
    io_A_Valid_4_delay_1_41 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_40 <= io_A_Valid_4_delay_1_41;
    io_A_Valid_4_delay_3_39 <= io_A_Valid_4_delay_2_40;
    io_A_Valid_4_delay_4_38 <= io_A_Valid_4_delay_3_39;
    io_A_Valid_4_delay_5_37 <= io_A_Valid_4_delay_4_38;
    io_A_Valid_4_delay_6_36 <= io_A_Valid_4_delay_5_37;
    io_A_Valid_4_delay_7_35 <= io_A_Valid_4_delay_6_36;
    io_A_Valid_4_delay_8_34 <= io_A_Valid_4_delay_7_35;
    io_A_Valid_4_delay_9_33 <= io_A_Valid_4_delay_8_34;
    io_A_Valid_4_delay_10_32 <= io_A_Valid_4_delay_9_33;
    io_A_Valid_4_delay_11_31 <= io_A_Valid_4_delay_10_32;
    io_A_Valid_4_delay_12_30 <= io_A_Valid_4_delay_11_31;
    io_A_Valid_4_delay_13_29 <= io_A_Valid_4_delay_12_30;
    io_A_Valid_4_delay_14_28 <= io_A_Valid_4_delay_13_29;
    io_A_Valid_4_delay_15_27 <= io_A_Valid_4_delay_14_28;
    io_A_Valid_4_delay_16_26 <= io_A_Valid_4_delay_15_27;
    io_A_Valid_4_delay_17_25 <= io_A_Valid_4_delay_16_26;
    io_A_Valid_4_delay_18_24 <= io_A_Valid_4_delay_17_25;
    io_A_Valid_4_delay_19_23 <= io_A_Valid_4_delay_18_24;
    io_A_Valid_4_delay_20_22 <= io_A_Valid_4_delay_19_23;
    io_A_Valid_4_delay_21_21 <= io_A_Valid_4_delay_20_22;
    io_A_Valid_4_delay_22_20 <= io_A_Valid_4_delay_21_21;
    io_A_Valid_4_delay_23_19 <= io_A_Valid_4_delay_22_20;
    io_A_Valid_4_delay_24_18 <= io_A_Valid_4_delay_23_19;
    io_A_Valid_4_delay_25_17 <= io_A_Valid_4_delay_24_18;
    io_A_Valid_4_delay_26_16 <= io_A_Valid_4_delay_25_17;
    io_A_Valid_4_delay_27_15 <= io_A_Valid_4_delay_26_16;
    io_A_Valid_4_delay_28_14 <= io_A_Valid_4_delay_27_15;
    io_A_Valid_4_delay_29_13 <= io_A_Valid_4_delay_28_14;
    io_A_Valid_4_delay_30_12 <= io_A_Valid_4_delay_29_13;
    io_A_Valid_4_delay_31_11 <= io_A_Valid_4_delay_30_12;
    io_A_Valid_4_delay_32_10 <= io_A_Valid_4_delay_31_11;
    io_A_Valid_4_delay_33_9 <= io_A_Valid_4_delay_32_10;
    io_A_Valid_4_delay_34_8 <= io_A_Valid_4_delay_33_9;
    io_A_Valid_4_delay_35_7 <= io_A_Valid_4_delay_34_8;
    io_A_Valid_4_delay_36_6 <= io_A_Valid_4_delay_35_7;
    io_A_Valid_4_delay_37_5 <= io_A_Valid_4_delay_36_6;
    io_A_Valid_4_delay_38_4 <= io_A_Valid_4_delay_37_5;
    io_A_Valid_4_delay_39_3 <= io_A_Valid_4_delay_38_4;
    io_A_Valid_4_delay_40_2 <= io_A_Valid_4_delay_39_3;
    io_A_Valid_4_delay_41_1 <= io_A_Valid_4_delay_40_2;
    io_A_Valid_4_delay_42 <= io_A_Valid_4_delay_41_1;
    io_B_Valid_42_delay_1_3 <= io_B_Valid_42;
    io_B_Valid_42_delay_2_2 <= io_B_Valid_42_delay_1_3;
    io_B_Valid_42_delay_3_1 <= io_B_Valid_42_delay_2_2;
    io_B_Valid_42_delay_4 <= io_B_Valid_42_delay_3_1;
    io_A_Valid_4_delay_1_42 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_41 <= io_A_Valid_4_delay_1_42;
    io_A_Valid_4_delay_3_40 <= io_A_Valid_4_delay_2_41;
    io_A_Valid_4_delay_4_39 <= io_A_Valid_4_delay_3_40;
    io_A_Valid_4_delay_5_38 <= io_A_Valid_4_delay_4_39;
    io_A_Valid_4_delay_6_37 <= io_A_Valid_4_delay_5_38;
    io_A_Valid_4_delay_7_36 <= io_A_Valid_4_delay_6_37;
    io_A_Valid_4_delay_8_35 <= io_A_Valid_4_delay_7_36;
    io_A_Valid_4_delay_9_34 <= io_A_Valid_4_delay_8_35;
    io_A_Valid_4_delay_10_33 <= io_A_Valid_4_delay_9_34;
    io_A_Valid_4_delay_11_32 <= io_A_Valid_4_delay_10_33;
    io_A_Valid_4_delay_12_31 <= io_A_Valid_4_delay_11_32;
    io_A_Valid_4_delay_13_30 <= io_A_Valid_4_delay_12_31;
    io_A_Valid_4_delay_14_29 <= io_A_Valid_4_delay_13_30;
    io_A_Valid_4_delay_15_28 <= io_A_Valid_4_delay_14_29;
    io_A_Valid_4_delay_16_27 <= io_A_Valid_4_delay_15_28;
    io_A_Valid_4_delay_17_26 <= io_A_Valid_4_delay_16_27;
    io_A_Valid_4_delay_18_25 <= io_A_Valid_4_delay_17_26;
    io_A_Valid_4_delay_19_24 <= io_A_Valid_4_delay_18_25;
    io_A_Valid_4_delay_20_23 <= io_A_Valid_4_delay_19_24;
    io_A_Valid_4_delay_21_22 <= io_A_Valid_4_delay_20_23;
    io_A_Valid_4_delay_22_21 <= io_A_Valid_4_delay_21_22;
    io_A_Valid_4_delay_23_20 <= io_A_Valid_4_delay_22_21;
    io_A_Valid_4_delay_24_19 <= io_A_Valid_4_delay_23_20;
    io_A_Valid_4_delay_25_18 <= io_A_Valid_4_delay_24_19;
    io_A_Valid_4_delay_26_17 <= io_A_Valid_4_delay_25_18;
    io_A_Valid_4_delay_27_16 <= io_A_Valid_4_delay_26_17;
    io_A_Valid_4_delay_28_15 <= io_A_Valid_4_delay_27_16;
    io_A_Valid_4_delay_29_14 <= io_A_Valid_4_delay_28_15;
    io_A_Valid_4_delay_30_13 <= io_A_Valid_4_delay_29_14;
    io_A_Valid_4_delay_31_12 <= io_A_Valid_4_delay_30_13;
    io_A_Valid_4_delay_32_11 <= io_A_Valid_4_delay_31_12;
    io_A_Valid_4_delay_33_10 <= io_A_Valid_4_delay_32_11;
    io_A_Valid_4_delay_34_9 <= io_A_Valid_4_delay_33_10;
    io_A_Valid_4_delay_35_8 <= io_A_Valid_4_delay_34_9;
    io_A_Valid_4_delay_36_7 <= io_A_Valid_4_delay_35_8;
    io_A_Valid_4_delay_37_6 <= io_A_Valid_4_delay_36_7;
    io_A_Valid_4_delay_38_5 <= io_A_Valid_4_delay_37_6;
    io_A_Valid_4_delay_39_4 <= io_A_Valid_4_delay_38_5;
    io_A_Valid_4_delay_40_3 <= io_A_Valid_4_delay_39_4;
    io_A_Valid_4_delay_41_2 <= io_A_Valid_4_delay_40_3;
    io_A_Valid_4_delay_42_1 <= io_A_Valid_4_delay_41_2;
    io_A_Valid_4_delay_43 <= io_A_Valid_4_delay_42_1;
    io_B_Valid_43_delay_1_3 <= io_B_Valid_43;
    io_B_Valid_43_delay_2_2 <= io_B_Valid_43_delay_1_3;
    io_B_Valid_43_delay_3_1 <= io_B_Valid_43_delay_2_2;
    io_B_Valid_43_delay_4 <= io_B_Valid_43_delay_3_1;
    io_A_Valid_4_delay_1_43 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_42 <= io_A_Valid_4_delay_1_43;
    io_A_Valid_4_delay_3_41 <= io_A_Valid_4_delay_2_42;
    io_A_Valid_4_delay_4_40 <= io_A_Valid_4_delay_3_41;
    io_A_Valid_4_delay_5_39 <= io_A_Valid_4_delay_4_40;
    io_A_Valid_4_delay_6_38 <= io_A_Valid_4_delay_5_39;
    io_A_Valid_4_delay_7_37 <= io_A_Valid_4_delay_6_38;
    io_A_Valid_4_delay_8_36 <= io_A_Valid_4_delay_7_37;
    io_A_Valid_4_delay_9_35 <= io_A_Valid_4_delay_8_36;
    io_A_Valid_4_delay_10_34 <= io_A_Valid_4_delay_9_35;
    io_A_Valid_4_delay_11_33 <= io_A_Valid_4_delay_10_34;
    io_A_Valid_4_delay_12_32 <= io_A_Valid_4_delay_11_33;
    io_A_Valid_4_delay_13_31 <= io_A_Valid_4_delay_12_32;
    io_A_Valid_4_delay_14_30 <= io_A_Valid_4_delay_13_31;
    io_A_Valid_4_delay_15_29 <= io_A_Valid_4_delay_14_30;
    io_A_Valid_4_delay_16_28 <= io_A_Valid_4_delay_15_29;
    io_A_Valid_4_delay_17_27 <= io_A_Valid_4_delay_16_28;
    io_A_Valid_4_delay_18_26 <= io_A_Valid_4_delay_17_27;
    io_A_Valid_4_delay_19_25 <= io_A_Valid_4_delay_18_26;
    io_A_Valid_4_delay_20_24 <= io_A_Valid_4_delay_19_25;
    io_A_Valid_4_delay_21_23 <= io_A_Valid_4_delay_20_24;
    io_A_Valid_4_delay_22_22 <= io_A_Valid_4_delay_21_23;
    io_A_Valid_4_delay_23_21 <= io_A_Valid_4_delay_22_22;
    io_A_Valid_4_delay_24_20 <= io_A_Valid_4_delay_23_21;
    io_A_Valid_4_delay_25_19 <= io_A_Valid_4_delay_24_20;
    io_A_Valid_4_delay_26_18 <= io_A_Valid_4_delay_25_19;
    io_A_Valid_4_delay_27_17 <= io_A_Valid_4_delay_26_18;
    io_A_Valid_4_delay_28_16 <= io_A_Valid_4_delay_27_17;
    io_A_Valid_4_delay_29_15 <= io_A_Valid_4_delay_28_16;
    io_A_Valid_4_delay_30_14 <= io_A_Valid_4_delay_29_15;
    io_A_Valid_4_delay_31_13 <= io_A_Valid_4_delay_30_14;
    io_A_Valid_4_delay_32_12 <= io_A_Valid_4_delay_31_13;
    io_A_Valid_4_delay_33_11 <= io_A_Valid_4_delay_32_12;
    io_A_Valid_4_delay_34_10 <= io_A_Valid_4_delay_33_11;
    io_A_Valid_4_delay_35_9 <= io_A_Valid_4_delay_34_10;
    io_A_Valid_4_delay_36_8 <= io_A_Valid_4_delay_35_9;
    io_A_Valid_4_delay_37_7 <= io_A_Valid_4_delay_36_8;
    io_A_Valid_4_delay_38_6 <= io_A_Valid_4_delay_37_7;
    io_A_Valid_4_delay_39_5 <= io_A_Valid_4_delay_38_6;
    io_A_Valid_4_delay_40_4 <= io_A_Valid_4_delay_39_5;
    io_A_Valid_4_delay_41_3 <= io_A_Valid_4_delay_40_4;
    io_A_Valid_4_delay_42_2 <= io_A_Valid_4_delay_41_3;
    io_A_Valid_4_delay_43_1 <= io_A_Valid_4_delay_42_2;
    io_A_Valid_4_delay_44 <= io_A_Valid_4_delay_43_1;
    io_B_Valid_44_delay_1_3 <= io_B_Valid_44;
    io_B_Valid_44_delay_2_2 <= io_B_Valid_44_delay_1_3;
    io_B_Valid_44_delay_3_1 <= io_B_Valid_44_delay_2_2;
    io_B_Valid_44_delay_4 <= io_B_Valid_44_delay_3_1;
    io_A_Valid_4_delay_1_44 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_43 <= io_A_Valid_4_delay_1_44;
    io_A_Valid_4_delay_3_42 <= io_A_Valid_4_delay_2_43;
    io_A_Valid_4_delay_4_41 <= io_A_Valid_4_delay_3_42;
    io_A_Valid_4_delay_5_40 <= io_A_Valid_4_delay_4_41;
    io_A_Valid_4_delay_6_39 <= io_A_Valid_4_delay_5_40;
    io_A_Valid_4_delay_7_38 <= io_A_Valid_4_delay_6_39;
    io_A_Valid_4_delay_8_37 <= io_A_Valid_4_delay_7_38;
    io_A_Valid_4_delay_9_36 <= io_A_Valid_4_delay_8_37;
    io_A_Valid_4_delay_10_35 <= io_A_Valid_4_delay_9_36;
    io_A_Valid_4_delay_11_34 <= io_A_Valid_4_delay_10_35;
    io_A_Valid_4_delay_12_33 <= io_A_Valid_4_delay_11_34;
    io_A_Valid_4_delay_13_32 <= io_A_Valid_4_delay_12_33;
    io_A_Valid_4_delay_14_31 <= io_A_Valid_4_delay_13_32;
    io_A_Valid_4_delay_15_30 <= io_A_Valid_4_delay_14_31;
    io_A_Valid_4_delay_16_29 <= io_A_Valid_4_delay_15_30;
    io_A_Valid_4_delay_17_28 <= io_A_Valid_4_delay_16_29;
    io_A_Valid_4_delay_18_27 <= io_A_Valid_4_delay_17_28;
    io_A_Valid_4_delay_19_26 <= io_A_Valid_4_delay_18_27;
    io_A_Valid_4_delay_20_25 <= io_A_Valid_4_delay_19_26;
    io_A_Valid_4_delay_21_24 <= io_A_Valid_4_delay_20_25;
    io_A_Valid_4_delay_22_23 <= io_A_Valid_4_delay_21_24;
    io_A_Valid_4_delay_23_22 <= io_A_Valid_4_delay_22_23;
    io_A_Valid_4_delay_24_21 <= io_A_Valid_4_delay_23_22;
    io_A_Valid_4_delay_25_20 <= io_A_Valid_4_delay_24_21;
    io_A_Valid_4_delay_26_19 <= io_A_Valid_4_delay_25_20;
    io_A_Valid_4_delay_27_18 <= io_A_Valid_4_delay_26_19;
    io_A_Valid_4_delay_28_17 <= io_A_Valid_4_delay_27_18;
    io_A_Valid_4_delay_29_16 <= io_A_Valid_4_delay_28_17;
    io_A_Valid_4_delay_30_15 <= io_A_Valid_4_delay_29_16;
    io_A_Valid_4_delay_31_14 <= io_A_Valid_4_delay_30_15;
    io_A_Valid_4_delay_32_13 <= io_A_Valid_4_delay_31_14;
    io_A_Valid_4_delay_33_12 <= io_A_Valid_4_delay_32_13;
    io_A_Valid_4_delay_34_11 <= io_A_Valid_4_delay_33_12;
    io_A_Valid_4_delay_35_10 <= io_A_Valid_4_delay_34_11;
    io_A_Valid_4_delay_36_9 <= io_A_Valid_4_delay_35_10;
    io_A_Valid_4_delay_37_8 <= io_A_Valid_4_delay_36_9;
    io_A_Valid_4_delay_38_7 <= io_A_Valid_4_delay_37_8;
    io_A_Valid_4_delay_39_6 <= io_A_Valid_4_delay_38_7;
    io_A_Valid_4_delay_40_5 <= io_A_Valid_4_delay_39_6;
    io_A_Valid_4_delay_41_4 <= io_A_Valid_4_delay_40_5;
    io_A_Valid_4_delay_42_3 <= io_A_Valid_4_delay_41_4;
    io_A_Valid_4_delay_43_2 <= io_A_Valid_4_delay_42_3;
    io_A_Valid_4_delay_44_1 <= io_A_Valid_4_delay_43_2;
    io_A_Valid_4_delay_45 <= io_A_Valid_4_delay_44_1;
    io_B_Valid_45_delay_1_3 <= io_B_Valid_45;
    io_B_Valid_45_delay_2_2 <= io_B_Valid_45_delay_1_3;
    io_B_Valid_45_delay_3_1 <= io_B_Valid_45_delay_2_2;
    io_B_Valid_45_delay_4 <= io_B_Valid_45_delay_3_1;
    io_A_Valid_4_delay_1_45 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_44 <= io_A_Valid_4_delay_1_45;
    io_A_Valid_4_delay_3_43 <= io_A_Valid_4_delay_2_44;
    io_A_Valid_4_delay_4_42 <= io_A_Valid_4_delay_3_43;
    io_A_Valid_4_delay_5_41 <= io_A_Valid_4_delay_4_42;
    io_A_Valid_4_delay_6_40 <= io_A_Valid_4_delay_5_41;
    io_A_Valid_4_delay_7_39 <= io_A_Valid_4_delay_6_40;
    io_A_Valid_4_delay_8_38 <= io_A_Valid_4_delay_7_39;
    io_A_Valid_4_delay_9_37 <= io_A_Valid_4_delay_8_38;
    io_A_Valid_4_delay_10_36 <= io_A_Valid_4_delay_9_37;
    io_A_Valid_4_delay_11_35 <= io_A_Valid_4_delay_10_36;
    io_A_Valid_4_delay_12_34 <= io_A_Valid_4_delay_11_35;
    io_A_Valid_4_delay_13_33 <= io_A_Valid_4_delay_12_34;
    io_A_Valid_4_delay_14_32 <= io_A_Valid_4_delay_13_33;
    io_A_Valid_4_delay_15_31 <= io_A_Valid_4_delay_14_32;
    io_A_Valid_4_delay_16_30 <= io_A_Valid_4_delay_15_31;
    io_A_Valid_4_delay_17_29 <= io_A_Valid_4_delay_16_30;
    io_A_Valid_4_delay_18_28 <= io_A_Valid_4_delay_17_29;
    io_A_Valid_4_delay_19_27 <= io_A_Valid_4_delay_18_28;
    io_A_Valid_4_delay_20_26 <= io_A_Valid_4_delay_19_27;
    io_A_Valid_4_delay_21_25 <= io_A_Valid_4_delay_20_26;
    io_A_Valid_4_delay_22_24 <= io_A_Valid_4_delay_21_25;
    io_A_Valid_4_delay_23_23 <= io_A_Valid_4_delay_22_24;
    io_A_Valid_4_delay_24_22 <= io_A_Valid_4_delay_23_23;
    io_A_Valid_4_delay_25_21 <= io_A_Valid_4_delay_24_22;
    io_A_Valid_4_delay_26_20 <= io_A_Valid_4_delay_25_21;
    io_A_Valid_4_delay_27_19 <= io_A_Valid_4_delay_26_20;
    io_A_Valid_4_delay_28_18 <= io_A_Valid_4_delay_27_19;
    io_A_Valid_4_delay_29_17 <= io_A_Valid_4_delay_28_18;
    io_A_Valid_4_delay_30_16 <= io_A_Valid_4_delay_29_17;
    io_A_Valid_4_delay_31_15 <= io_A_Valid_4_delay_30_16;
    io_A_Valid_4_delay_32_14 <= io_A_Valid_4_delay_31_15;
    io_A_Valid_4_delay_33_13 <= io_A_Valid_4_delay_32_14;
    io_A_Valid_4_delay_34_12 <= io_A_Valid_4_delay_33_13;
    io_A_Valid_4_delay_35_11 <= io_A_Valid_4_delay_34_12;
    io_A_Valid_4_delay_36_10 <= io_A_Valid_4_delay_35_11;
    io_A_Valid_4_delay_37_9 <= io_A_Valid_4_delay_36_10;
    io_A_Valid_4_delay_38_8 <= io_A_Valid_4_delay_37_9;
    io_A_Valid_4_delay_39_7 <= io_A_Valid_4_delay_38_8;
    io_A_Valid_4_delay_40_6 <= io_A_Valid_4_delay_39_7;
    io_A_Valid_4_delay_41_5 <= io_A_Valid_4_delay_40_6;
    io_A_Valid_4_delay_42_4 <= io_A_Valid_4_delay_41_5;
    io_A_Valid_4_delay_43_3 <= io_A_Valid_4_delay_42_4;
    io_A_Valid_4_delay_44_2 <= io_A_Valid_4_delay_43_3;
    io_A_Valid_4_delay_45_1 <= io_A_Valid_4_delay_44_2;
    io_A_Valid_4_delay_46 <= io_A_Valid_4_delay_45_1;
    io_B_Valid_46_delay_1_3 <= io_B_Valid_46;
    io_B_Valid_46_delay_2_2 <= io_B_Valid_46_delay_1_3;
    io_B_Valid_46_delay_3_1 <= io_B_Valid_46_delay_2_2;
    io_B_Valid_46_delay_4 <= io_B_Valid_46_delay_3_1;
    io_A_Valid_4_delay_1_46 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_45 <= io_A_Valid_4_delay_1_46;
    io_A_Valid_4_delay_3_44 <= io_A_Valid_4_delay_2_45;
    io_A_Valid_4_delay_4_43 <= io_A_Valid_4_delay_3_44;
    io_A_Valid_4_delay_5_42 <= io_A_Valid_4_delay_4_43;
    io_A_Valid_4_delay_6_41 <= io_A_Valid_4_delay_5_42;
    io_A_Valid_4_delay_7_40 <= io_A_Valid_4_delay_6_41;
    io_A_Valid_4_delay_8_39 <= io_A_Valid_4_delay_7_40;
    io_A_Valid_4_delay_9_38 <= io_A_Valid_4_delay_8_39;
    io_A_Valid_4_delay_10_37 <= io_A_Valid_4_delay_9_38;
    io_A_Valid_4_delay_11_36 <= io_A_Valid_4_delay_10_37;
    io_A_Valid_4_delay_12_35 <= io_A_Valid_4_delay_11_36;
    io_A_Valid_4_delay_13_34 <= io_A_Valid_4_delay_12_35;
    io_A_Valid_4_delay_14_33 <= io_A_Valid_4_delay_13_34;
    io_A_Valid_4_delay_15_32 <= io_A_Valid_4_delay_14_33;
    io_A_Valid_4_delay_16_31 <= io_A_Valid_4_delay_15_32;
    io_A_Valid_4_delay_17_30 <= io_A_Valid_4_delay_16_31;
    io_A_Valid_4_delay_18_29 <= io_A_Valid_4_delay_17_30;
    io_A_Valid_4_delay_19_28 <= io_A_Valid_4_delay_18_29;
    io_A_Valid_4_delay_20_27 <= io_A_Valid_4_delay_19_28;
    io_A_Valid_4_delay_21_26 <= io_A_Valid_4_delay_20_27;
    io_A_Valid_4_delay_22_25 <= io_A_Valid_4_delay_21_26;
    io_A_Valid_4_delay_23_24 <= io_A_Valid_4_delay_22_25;
    io_A_Valid_4_delay_24_23 <= io_A_Valid_4_delay_23_24;
    io_A_Valid_4_delay_25_22 <= io_A_Valid_4_delay_24_23;
    io_A_Valid_4_delay_26_21 <= io_A_Valid_4_delay_25_22;
    io_A_Valid_4_delay_27_20 <= io_A_Valid_4_delay_26_21;
    io_A_Valid_4_delay_28_19 <= io_A_Valid_4_delay_27_20;
    io_A_Valid_4_delay_29_18 <= io_A_Valid_4_delay_28_19;
    io_A_Valid_4_delay_30_17 <= io_A_Valid_4_delay_29_18;
    io_A_Valid_4_delay_31_16 <= io_A_Valid_4_delay_30_17;
    io_A_Valid_4_delay_32_15 <= io_A_Valid_4_delay_31_16;
    io_A_Valid_4_delay_33_14 <= io_A_Valid_4_delay_32_15;
    io_A_Valid_4_delay_34_13 <= io_A_Valid_4_delay_33_14;
    io_A_Valid_4_delay_35_12 <= io_A_Valid_4_delay_34_13;
    io_A_Valid_4_delay_36_11 <= io_A_Valid_4_delay_35_12;
    io_A_Valid_4_delay_37_10 <= io_A_Valid_4_delay_36_11;
    io_A_Valid_4_delay_38_9 <= io_A_Valid_4_delay_37_10;
    io_A_Valid_4_delay_39_8 <= io_A_Valid_4_delay_38_9;
    io_A_Valid_4_delay_40_7 <= io_A_Valid_4_delay_39_8;
    io_A_Valid_4_delay_41_6 <= io_A_Valid_4_delay_40_7;
    io_A_Valid_4_delay_42_5 <= io_A_Valid_4_delay_41_6;
    io_A_Valid_4_delay_43_4 <= io_A_Valid_4_delay_42_5;
    io_A_Valid_4_delay_44_3 <= io_A_Valid_4_delay_43_4;
    io_A_Valid_4_delay_45_2 <= io_A_Valid_4_delay_44_3;
    io_A_Valid_4_delay_46_1 <= io_A_Valid_4_delay_45_2;
    io_A_Valid_4_delay_47 <= io_A_Valid_4_delay_46_1;
    io_B_Valid_47_delay_1_3 <= io_B_Valid_47;
    io_B_Valid_47_delay_2_2 <= io_B_Valid_47_delay_1_3;
    io_B_Valid_47_delay_3_1 <= io_B_Valid_47_delay_2_2;
    io_B_Valid_47_delay_4 <= io_B_Valid_47_delay_3_1;
    io_A_Valid_4_delay_1_47 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_46 <= io_A_Valid_4_delay_1_47;
    io_A_Valid_4_delay_3_45 <= io_A_Valid_4_delay_2_46;
    io_A_Valid_4_delay_4_44 <= io_A_Valid_4_delay_3_45;
    io_A_Valid_4_delay_5_43 <= io_A_Valid_4_delay_4_44;
    io_A_Valid_4_delay_6_42 <= io_A_Valid_4_delay_5_43;
    io_A_Valid_4_delay_7_41 <= io_A_Valid_4_delay_6_42;
    io_A_Valid_4_delay_8_40 <= io_A_Valid_4_delay_7_41;
    io_A_Valid_4_delay_9_39 <= io_A_Valid_4_delay_8_40;
    io_A_Valid_4_delay_10_38 <= io_A_Valid_4_delay_9_39;
    io_A_Valid_4_delay_11_37 <= io_A_Valid_4_delay_10_38;
    io_A_Valid_4_delay_12_36 <= io_A_Valid_4_delay_11_37;
    io_A_Valid_4_delay_13_35 <= io_A_Valid_4_delay_12_36;
    io_A_Valid_4_delay_14_34 <= io_A_Valid_4_delay_13_35;
    io_A_Valid_4_delay_15_33 <= io_A_Valid_4_delay_14_34;
    io_A_Valid_4_delay_16_32 <= io_A_Valid_4_delay_15_33;
    io_A_Valid_4_delay_17_31 <= io_A_Valid_4_delay_16_32;
    io_A_Valid_4_delay_18_30 <= io_A_Valid_4_delay_17_31;
    io_A_Valid_4_delay_19_29 <= io_A_Valid_4_delay_18_30;
    io_A_Valid_4_delay_20_28 <= io_A_Valid_4_delay_19_29;
    io_A_Valid_4_delay_21_27 <= io_A_Valid_4_delay_20_28;
    io_A_Valid_4_delay_22_26 <= io_A_Valid_4_delay_21_27;
    io_A_Valid_4_delay_23_25 <= io_A_Valid_4_delay_22_26;
    io_A_Valid_4_delay_24_24 <= io_A_Valid_4_delay_23_25;
    io_A_Valid_4_delay_25_23 <= io_A_Valid_4_delay_24_24;
    io_A_Valid_4_delay_26_22 <= io_A_Valid_4_delay_25_23;
    io_A_Valid_4_delay_27_21 <= io_A_Valid_4_delay_26_22;
    io_A_Valid_4_delay_28_20 <= io_A_Valid_4_delay_27_21;
    io_A_Valid_4_delay_29_19 <= io_A_Valid_4_delay_28_20;
    io_A_Valid_4_delay_30_18 <= io_A_Valid_4_delay_29_19;
    io_A_Valid_4_delay_31_17 <= io_A_Valid_4_delay_30_18;
    io_A_Valid_4_delay_32_16 <= io_A_Valid_4_delay_31_17;
    io_A_Valid_4_delay_33_15 <= io_A_Valid_4_delay_32_16;
    io_A_Valid_4_delay_34_14 <= io_A_Valid_4_delay_33_15;
    io_A_Valid_4_delay_35_13 <= io_A_Valid_4_delay_34_14;
    io_A_Valid_4_delay_36_12 <= io_A_Valid_4_delay_35_13;
    io_A_Valid_4_delay_37_11 <= io_A_Valid_4_delay_36_12;
    io_A_Valid_4_delay_38_10 <= io_A_Valid_4_delay_37_11;
    io_A_Valid_4_delay_39_9 <= io_A_Valid_4_delay_38_10;
    io_A_Valid_4_delay_40_8 <= io_A_Valid_4_delay_39_9;
    io_A_Valid_4_delay_41_7 <= io_A_Valid_4_delay_40_8;
    io_A_Valid_4_delay_42_6 <= io_A_Valid_4_delay_41_7;
    io_A_Valid_4_delay_43_5 <= io_A_Valid_4_delay_42_6;
    io_A_Valid_4_delay_44_4 <= io_A_Valid_4_delay_43_5;
    io_A_Valid_4_delay_45_3 <= io_A_Valid_4_delay_44_4;
    io_A_Valid_4_delay_46_2 <= io_A_Valid_4_delay_45_3;
    io_A_Valid_4_delay_47_1 <= io_A_Valid_4_delay_46_2;
    io_A_Valid_4_delay_48 <= io_A_Valid_4_delay_47_1;
    io_B_Valid_48_delay_1_3 <= io_B_Valid_48;
    io_B_Valid_48_delay_2_2 <= io_B_Valid_48_delay_1_3;
    io_B_Valid_48_delay_3_1 <= io_B_Valid_48_delay_2_2;
    io_B_Valid_48_delay_4 <= io_B_Valid_48_delay_3_1;
    io_A_Valid_4_delay_1_48 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_47 <= io_A_Valid_4_delay_1_48;
    io_A_Valid_4_delay_3_46 <= io_A_Valid_4_delay_2_47;
    io_A_Valid_4_delay_4_45 <= io_A_Valid_4_delay_3_46;
    io_A_Valid_4_delay_5_44 <= io_A_Valid_4_delay_4_45;
    io_A_Valid_4_delay_6_43 <= io_A_Valid_4_delay_5_44;
    io_A_Valid_4_delay_7_42 <= io_A_Valid_4_delay_6_43;
    io_A_Valid_4_delay_8_41 <= io_A_Valid_4_delay_7_42;
    io_A_Valid_4_delay_9_40 <= io_A_Valid_4_delay_8_41;
    io_A_Valid_4_delay_10_39 <= io_A_Valid_4_delay_9_40;
    io_A_Valid_4_delay_11_38 <= io_A_Valid_4_delay_10_39;
    io_A_Valid_4_delay_12_37 <= io_A_Valid_4_delay_11_38;
    io_A_Valid_4_delay_13_36 <= io_A_Valid_4_delay_12_37;
    io_A_Valid_4_delay_14_35 <= io_A_Valid_4_delay_13_36;
    io_A_Valid_4_delay_15_34 <= io_A_Valid_4_delay_14_35;
    io_A_Valid_4_delay_16_33 <= io_A_Valid_4_delay_15_34;
    io_A_Valid_4_delay_17_32 <= io_A_Valid_4_delay_16_33;
    io_A_Valid_4_delay_18_31 <= io_A_Valid_4_delay_17_32;
    io_A_Valid_4_delay_19_30 <= io_A_Valid_4_delay_18_31;
    io_A_Valid_4_delay_20_29 <= io_A_Valid_4_delay_19_30;
    io_A_Valid_4_delay_21_28 <= io_A_Valid_4_delay_20_29;
    io_A_Valid_4_delay_22_27 <= io_A_Valid_4_delay_21_28;
    io_A_Valid_4_delay_23_26 <= io_A_Valid_4_delay_22_27;
    io_A_Valid_4_delay_24_25 <= io_A_Valid_4_delay_23_26;
    io_A_Valid_4_delay_25_24 <= io_A_Valid_4_delay_24_25;
    io_A_Valid_4_delay_26_23 <= io_A_Valid_4_delay_25_24;
    io_A_Valid_4_delay_27_22 <= io_A_Valid_4_delay_26_23;
    io_A_Valid_4_delay_28_21 <= io_A_Valid_4_delay_27_22;
    io_A_Valid_4_delay_29_20 <= io_A_Valid_4_delay_28_21;
    io_A_Valid_4_delay_30_19 <= io_A_Valid_4_delay_29_20;
    io_A_Valid_4_delay_31_18 <= io_A_Valid_4_delay_30_19;
    io_A_Valid_4_delay_32_17 <= io_A_Valid_4_delay_31_18;
    io_A_Valid_4_delay_33_16 <= io_A_Valid_4_delay_32_17;
    io_A_Valid_4_delay_34_15 <= io_A_Valid_4_delay_33_16;
    io_A_Valid_4_delay_35_14 <= io_A_Valid_4_delay_34_15;
    io_A_Valid_4_delay_36_13 <= io_A_Valid_4_delay_35_14;
    io_A_Valid_4_delay_37_12 <= io_A_Valid_4_delay_36_13;
    io_A_Valid_4_delay_38_11 <= io_A_Valid_4_delay_37_12;
    io_A_Valid_4_delay_39_10 <= io_A_Valid_4_delay_38_11;
    io_A_Valid_4_delay_40_9 <= io_A_Valid_4_delay_39_10;
    io_A_Valid_4_delay_41_8 <= io_A_Valid_4_delay_40_9;
    io_A_Valid_4_delay_42_7 <= io_A_Valid_4_delay_41_8;
    io_A_Valid_4_delay_43_6 <= io_A_Valid_4_delay_42_7;
    io_A_Valid_4_delay_44_5 <= io_A_Valid_4_delay_43_6;
    io_A_Valid_4_delay_45_4 <= io_A_Valid_4_delay_44_5;
    io_A_Valid_4_delay_46_3 <= io_A_Valid_4_delay_45_4;
    io_A_Valid_4_delay_47_2 <= io_A_Valid_4_delay_46_3;
    io_A_Valid_4_delay_48_1 <= io_A_Valid_4_delay_47_2;
    io_A_Valid_4_delay_49 <= io_A_Valid_4_delay_48_1;
    io_B_Valid_49_delay_1_3 <= io_B_Valid_49;
    io_B_Valid_49_delay_2_2 <= io_B_Valid_49_delay_1_3;
    io_B_Valid_49_delay_3_1 <= io_B_Valid_49_delay_2_2;
    io_B_Valid_49_delay_4 <= io_B_Valid_49_delay_3_1;
    io_A_Valid_4_delay_1_49 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_48 <= io_A_Valid_4_delay_1_49;
    io_A_Valid_4_delay_3_47 <= io_A_Valid_4_delay_2_48;
    io_A_Valid_4_delay_4_46 <= io_A_Valid_4_delay_3_47;
    io_A_Valid_4_delay_5_45 <= io_A_Valid_4_delay_4_46;
    io_A_Valid_4_delay_6_44 <= io_A_Valid_4_delay_5_45;
    io_A_Valid_4_delay_7_43 <= io_A_Valid_4_delay_6_44;
    io_A_Valid_4_delay_8_42 <= io_A_Valid_4_delay_7_43;
    io_A_Valid_4_delay_9_41 <= io_A_Valid_4_delay_8_42;
    io_A_Valid_4_delay_10_40 <= io_A_Valid_4_delay_9_41;
    io_A_Valid_4_delay_11_39 <= io_A_Valid_4_delay_10_40;
    io_A_Valid_4_delay_12_38 <= io_A_Valid_4_delay_11_39;
    io_A_Valid_4_delay_13_37 <= io_A_Valid_4_delay_12_38;
    io_A_Valid_4_delay_14_36 <= io_A_Valid_4_delay_13_37;
    io_A_Valid_4_delay_15_35 <= io_A_Valid_4_delay_14_36;
    io_A_Valid_4_delay_16_34 <= io_A_Valid_4_delay_15_35;
    io_A_Valid_4_delay_17_33 <= io_A_Valid_4_delay_16_34;
    io_A_Valid_4_delay_18_32 <= io_A_Valid_4_delay_17_33;
    io_A_Valid_4_delay_19_31 <= io_A_Valid_4_delay_18_32;
    io_A_Valid_4_delay_20_30 <= io_A_Valid_4_delay_19_31;
    io_A_Valid_4_delay_21_29 <= io_A_Valid_4_delay_20_30;
    io_A_Valid_4_delay_22_28 <= io_A_Valid_4_delay_21_29;
    io_A_Valid_4_delay_23_27 <= io_A_Valid_4_delay_22_28;
    io_A_Valid_4_delay_24_26 <= io_A_Valid_4_delay_23_27;
    io_A_Valid_4_delay_25_25 <= io_A_Valid_4_delay_24_26;
    io_A_Valid_4_delay_26_24 <= io_A_Valid_4_delay_25_25;
    io_A_Valid_4_delay_27_23 <= io_A_Valid_4_delay_26_24;
    io_A_Valid_4_delay_28_22 <= io_A_Valid_4_delay_27_23;
    io_A_Valid_4_delay_29_21 <= io_A_Valid_4_delay_28_22;
    io_A_Valid_4_delay_30_20 <= io_A_Valid_4_delay_29_21;
    io_A_Valid_4_delay_31_19 <= io_A_Valid_4_delay_30_20;
    io_A_Valid_4_delay_32_18 <= io_A_Valid_4_delay_31_19;
    io_A_Valid_4_delay_33_17 <= io_A_Valid_4_delay_32_18;
    io_A_Valid_4_delay_34_16 <= io_A_Valid_4_delay_33_17;
    io_A_Valid_4_delay_35_15 <= io_A_Valid_4_delay_34_16;
    io_A_Valid_4_delay_36_14 <= io_A_Valid_4_delay_35_15;
    io_A_Valid_4_delay_37_13 <= io_A_Valid_4_delay_36_14;
    io_A_Valid_4_delay_38_12 <= io_A_Valid_4_delay_37_13;
    io_A_Valid_4_delay_39_11 <= io_A_Valid_4_delay_38_12;
    io_A_Valid_4_delay_40_10 <= io_A_Valid_4_delay_39_11;
    io_A_Valid_4_delay_41_9 <= io_A_Valid_4_delay_40_10;
    io_A_Valid_4_delay_42_8 <= io_A_Valid_4_delay_41_9;
    io_A_Valid_4_delay_43_7 <= io_A_Valid_4_delay_42_8;
    io_A_Valid_4_delay_44_6 <= io_A_Valid_4_delay_43_7;
    io_A_Valid_4_delay_45_5 <= io_A_Valid_4_delay_44_6;
    io_A_Valid_4_delay_46_4 <= io_A_Valid_4_delay_45_5;
    io_A_Valid_4_delay_47_3 <= io_A_Valid_4_delay_46_4;
    io_A_Valid_4_delay_48_2 <= io_A_Valid_4_delay_47_3;
    io_A_Valid_4_delay_49_1 <= io_A_Valid_4_delay_48_2;
    io_A_Valid_4_delay_50 <= io_A_Valid_4_delay_49_1;
    io_B_Valid_50_delay_1_3 <= io_B_Valid_50;
    io_B_Valid_50_delay_2_2 <= io_B_Valid_50_delay_1_3;
    io_B_Valid_50_delay_3_1 <= io_B_Valid_50_delay_2_2;
    io_B_Valid_50_delay_4 <= io_B_Valid_50_delay_3_1;
    io_A_Valid_4_delay_1_50 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_49 <= io_A_Valid_4_delay_1_50;
    io_A_Valid_4_delay_3_48 <= io_A_Valid_4_delay_2_49;
    io_A_Valid_4_delay_4_47 <= io_A_Valid_4_delay_3_48;
    io_A_Valid_4_delay_5_46 <= io_A_Valid_4_delay_4_47;
    io_A_Valid_4_delay_6_45 <= io_A_Valid_4_delay_5_46;
    io_A_Valid_4_delay_7_44 <= io_A_Valid_4_delay_6_45;
    io_A_Valid_4_delay_8_43 <= io_A_Valid_4_delay_7_44;
    io_A_Valid_4_delay_9_42 <= io_A_Valid_4_delay_8_43;
    io_A_Valid_4_delay_10_41 <= io_A_Valid_4_delay_9_42;
    io_A_Valid_4_delay_11_40 <= io_A_Valid_4_delay_10_41;
    io_A_Valid_4_delay_12_39 <= io_A_Valid_4_delay_11_40;
    io_A_Valid_4_delay_13_38 <= io_A_Valid_4_delay_12_39;
    io_A_Valid_4_delay_14_37 <= io_A_Valid_4_delay_13_38;
    io_A_Valid_4_delay_15_36 <= io_A_Valid_4_delay_14_37;
    io_A_Valid_4_delay_16_35 <= io_A_Valid_4_delay_15_36;
    io_A_Valid_4_delay_17_34 <= io_A_Valid_4_delay_16_35;
    io_A_Valid_4_delay_18_33 <= io_A_Valid_4_delay_17_34;
    io_A_Valid_4_delay_19_32 <= io_A_Valid_4_delay_18_33;
    io_A_Valid_4_delay_20_31 <= io_A_Valid_4_delay_19_32;
    io_A_Valid_4_delay_21_30 <= io_A_Valid_4_delay_20_31;
    io_A_Valid_4_delay_22_29 <= io_A_Valid_4_delay_21_30;
    io_A_Valid_4_delay_23_28 <= io_A_Valid_4_delay_22_29;
    io_A_Valid_4_delay_24_27 <= io_A_Valid_4_delay_23_28;
    io_A_Valid_4_delay_25_26 <= io_A_Valid_4_delay_24_27;
    io_A_Valid_4_delay_26_25 <= io_A_Valid_4_delay_25_26;
    io_A_Valid_4_delay_27_24 <= io_A_Valid_4_delay_26_25;
    io_A_Valid_4_delay_28_23 <= io_A_Valid_4_delay_27_24;
    io_A_Valid_4_delay_29_22 <= io_A_Valid_4_delay_28_23;
    io_A_Valid_4_delay_30_21 <= io_A_Valid_4_delay_29_22;
    io_A_Valid_4_delay_31_20 <= io_A_Valid_4_delay_30_21;
    io_A_Valid_4_delay_32_19 <= io_A_Valid_4_delay_31_20;
    io_A_Valid_4_delay_33_18 <= io_A_Valid_4_delay_32_19;
    io_A_Valid_4_delay_34_17 <= io_A_Valid_4_delay_33_18;
    io_A_Valid_4_delay_35_16 <= io_A_Valid_4_delay_34_17;
    io_A_Valid_4_delay_36_15 <= io_A_Valid_4_delay_35_16;
    io_A_Valid_4_delay_37_14 <= io_A_Valid_4_delay_36_15;
    io_A_Valid_4_delay_38_13 <= io_A_Valid_4_delay_37_14;
    io_A_Valid_4_delay_39_12 <= io_A_Valid_4_delay_38_13;
    io_A_Valid_4_delay_40_11 <= io_A_Valid_4_delay_39_12;
    io_A_Valid_4_delay_41_10 <= io_A_Valid_4_delay_40_11;
    io_A_Valid_4_delay_42_9 <= io_A_Valid_4_delay_41_10;
    io_A_Valid_4_delay_43_8 <= io_A_Valid_4_delay_42_9;
    io_A_Valid_4_delay_44_7 <= io_A_Valid_4_delay_43_8;
    io_A_Valid_4_delay_45_6 <= io_A_Valid_4_delay_44_7;
    io_A_Valid_4_delay_46_5 <= io_A_Valid_4_delay_45_6;
    io_A_Valid_4_delay_47_4 <= io_A_Valid_4_delay_46_5;
    io_A_Valid_4_delay_48_3 <= io_A_Valid_4_delay_47_4;
    io_A_Valid_4_delay_49_2 <= io_A_Valid_4_delay_48_3;
    io_A_Valid_4_delay_50_1 <= io_A_Valid_4_delay_49_2;
    io_A_Valid_4_delay_51 <= io_A_Valid_4_delay_50_1;
    io_B_Valid_51_delay_1_3 <= io_B_Valid_51;
    io_B_Valid_51_delay_2_2 <= io_B_Valid_51_delay_1_3;
    io_B_Valid_51_delay_3_1 <= io_B_Valid_51_delay_2_2;
    io_B_Valid_51_delay_4 <= io_B_Valid_51_delay_3_1;
    io_A_Valid_4_delay_1_51 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_50 <= io_A_Valid_4_delay_1_51;
    io_A_Valid_4_delay_3_49 <= io_A_Valid_4_delay_2_50;
    io_A_Valid_4_delay_4_48 <= io_A_Valid_4_delay_3_49;
    io_A_Valid_4_delay_5_47 <= io_A_Valid_4_delay_4_48;
    io_A_Valid_4_delay_6_46 <= io_A_Valid_4_delay_5_47;
    io_A_Valid_4_delay_7_45 <= io_A_Valid_4_delay_6_46;
    io_A_Valid_4_delay_8_44 <= io_A_Valid_4_delay_7_45;
    io_A_Valid_4_delay_9_43 <= io_A_Valid_4_delay_8_44;
    io_A_Valid_4_delay_10_42 <= io_A_Valid_4_delay_9_43;
    io_A_Valid_4_delay_11_41 <= io_A_Valid_4_delay_10_42;
    io_A_Valid_4_delay_12_40 <= io_A_Valid_4_delay_11_41;
    io_A_Valid_4_delay_13_39 <= io_A_Valid_4_delay_12_40;
    io_A_Valid_4_delay_14_38 <= io_A_Valid_4_delay_13_39;
    io_A_Valid_4_delay_15_37 <= io_A_Valid_4_delay_14_38;
    io_A_Valid_4_delay_16_36 <= io_A_Valid_4_delay_15_37;
    io_A_Valid_4_delay_17_35 <= io_A_Valid_4_delay_16_36;
    io_A_Valid_4_delay_18_34 <= io_A_Valid_4_delay_17_35;
    io_A_Valid_4_delay_19_33 <= io_A_Valid_4_delay_18_34;
    io_A_Valid_4_delay_20_32 <= io_A_Valid_4_delay_19_33;
    io_A_Valid_4_delay_21_31 <= io_A_Valid_4_delay_20_32;
    io_A_Valid_4_delay_22_30 <= io_A_Valid_4_delay_21_31;
    io_A_Valid_4_delay_23_29 <= io_A_Valid_4_delay_22_30;
    io_A_Valid_4_delay_24_28 <= io_A_Valid_4_delay_23_29;
    io_A_Valid_4_delay_25_27 <= io_A_Valid_4_delay_24_28;
    io_A_Valid_4_delay_26_26 <= io_A_Valid_4_delay_25_27;
    io_A_Valid_4_delay_27_25 <= io_A_Valid_4_delay_26_26;
    io_A_Valid_4_delay_28_24 <= io_A_Valid_4_delay_27_25;
    io_A_Valid_4_delay_29_23 <= io_A_Valid_4_delay_28_24;
    io_A_Valid_4_delay_30_22 <= io_A_Valid_4_delay_29_23;
    io_A_Valid_4_delay_31_21 <= io_A_Valid_4_delay_30_22;
    io_A_Valid_4_delay_32_20 <= io_A_Valid_4_delay_31_21;
    io_A_Valid_4_delay_33_19 <= io_A_Valid_4_delay_32_20;
    io_A_Valid_4_delay_34_18 <= io_A_Valid_4_delay_33_19;
    io_A_Valid_4_delay_35_17 <= io_A_Valid_4_delay_34_18;
    io_A_Valid_4_delay_36_16 <= io_A_Valid_4_delay_35_17;
    io_A_Valid_4_delay_37_15 <= io_A_Valid_4_delay_36_16;
    io_A_Valid_4_delay_38_14 <= io_A_Valid_4_delay_37_15;
    io_A_Valid_4_delay_39_13 <= io_A_Valid_4_delay_38_14;
    io_A_Valid_4_delay_40_12 <= io_A_Valid_4_delay_39_13;
    io_A_Valid_4_delay_41_11 <= io_A_Valid_4_delay_40_12;
    io_A_Valid_4_delay_42_10 <= io_A_Valid_4_delay_41_11;
    io_A_Valid_4_delay_43_9 <= io_A_Valid_4_delay_42_10;
    io_A_Valid_4_delay_44_8 <= io_A_Valid_4_delay_43_9;
    io_A_Valid_4_delay_45_7 <= io_A_Valid_4_delay_44_8;
    io_A_Valid_4_delay_46_6 <= io_A_Valid_4_delay_45_7;
    io_A_Valid_4_delay_47_5 <= io_A_Valid_4_delay_46_6;
    io_A_Valid_4_delay_48_4 <= io_A_Valid_4_delay_47_5;
    io_A_Valid_4_delay_49_3 <= io_A_Valid_4_delay_48_4;
    io_A_Valid_4_delay_50_2 <= io_A_Valid_4_delay_49_3;
    io_A_Valid_4_delay_51_1 <= io_A_Valid_4_delay_50_2;
    io_A_Valid_4_delay_52 <= io_A_Valid_4_delay_51_1;
    io_B_Valid_52_delay_1_3 <= io_B_Valid_52;
    io_B_Valid_52_delay_2_2 <= io_B_Valid_52_delay_1_3;
    io_B_Valid_52_delay_3_1 <= io_B_Valid_52_delay_2_2;
    io_B_Valid_52_delay_4 <= io_B_Valid_52_delay_3_1;
    io_A_Valid_4_delay_1_52 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_51 <= io_A_Valid_4_delay_1_52;
    io_A_Valid_4_delay_3_50 <= io_A_Valid_4_delay_2_51;
    io_A_Valid_4_delay_4_49 <= io_A_Valid_4_delay_3_50;
    io_A_Valid_4_delay_5_48 <= io_A_Valid_4_delay_4_49;
    io_A_Valid_4_delay_6_47 <= io_A_Valid_4_delay_5_48;
    io_A_Valid_4_delay_7_46 <= io_A_Valid_4_delay_6_47;
    io_A_Valid_4_delay_8_45 <= io_A_Valid_4_delay_7_46;
    io_A_Valid_4_delay_9_44 <= io_A_Valid_4_delay_8_45;
    io_A_Valid_4_delay_10_43 <= io_A_Valid_4_delay_9_44;
    io_A_Valid_4_delay_11_42 <= io_A_Valid_4_delay_10_43;
    io_A_Valid_4_delay_12_41 <= io_A_Valid_4_delay_11_42;
    io_A_Valid_4_delay_13_40 <= io_A_Valid_4_delay_12_41;
    io_A_Valid_4_delay_14_39 <= io_A_Valid_4_delay_13_40;
    io_A_Valid_4_delay_15_38 <= io_A_Valid_4_delay_14_39;
    io_A_Valid_4_delay_16_37 <= io_A_Valid_4_delay_15_38;
    io_A_Valid_4_delay_17_36 <= io_A_Valid_4_delay_16_37;
    io_A_Valid_4_delay_18_35 <= io_A_Valid_4_delay_17_36;
    io_A_Valid_4_delay_19_34 <= io_A_Valid_4_delay_18_35;
    io_A_Valid_4_delay_20_33 <= io_A_Valid_4_delay_19_34;
    io_A_Valid_4_delay_21_32 <= io_A_Valid_4_delay_20_33;
    io_A_Valid_4_delay_22_31 <= io_A_Valid_4_delay_21_32;
    io_A_Valid_4_delay_23_30 <= io_A_Valid_4_delay_22_31;
    io_A_Valid_4_delay_24_29 <= io_A_Valid_4_delay_23_30;
    io_A_Valid_4_delay_25_28 <= io_A_Valid_4_delay_24_29;
    io_A_Valid_4_delay_26_27 <= io_A_Valid_4_delay_25_28;
    io_A_Valid_4_delay_27_26 <= io_A_Valid_4_delay_26_27;
    io_A_Valid_4_delay_28_25 <= io_A_Valid_4_delay_27_26;
    io_A_Valid_4_delay_29_24 <= io_A_Valid_4_delay_28_25;
    io_A_Valid_4_delay_30_23 <= io_A_Valid_4_delay_29_24;
    io_A_Valid_4_delay_31_22 <= io_A_Valid_4_delay_30_23;
    io_A_Valid_4_delay_32_21 <= io_A_Valid_4_delay_31_22;
    io_A_Valid_4_delay_33_20 <= io_A_Valid_4_delay_32_21;
    io_A_Valid_4_delay_34_19 <= io_A_Valid_4_delay_33_20;
    io_A_Valid_4_delay_35_18 <= io_A_Valid_4_delay_34_19;
    io_A_Valid_4_delay_36_17 <= io_A_Valid_4_delay_35_18;
    io_A_Valid_4_delay_37_16 <= io_A_Valid_4_delay_36_17;
    io_A_Valid_4_delay_38_15 <= io_A_Valid_4_delay_37_16;
    io_A_Valid_4_delay_39_14 <= io_A_Valid_4_delay_38_15;
    io_A_Valid_4_delay_40_13 <= io_A_Valid_4_delay_39_14;
    io_A_Valid_4_delay_41_12 <= io_A_Valid_4_delay_40_13;
    io_A_Valid_4_delay_42_11 <= io_A_Valid_4_delay_41_12;
    io_A_Valid_4_delay_43_10 <= io_A_Valid_4_delay_42_11;
    io_A_Valid_4_delay_44_9 <= io_A_Valid_4_delay_43_10;
    io_A_Valid_4_delay_45_8 <= io_A_Valid_4_delay_44_9;
    io_A_Valid_4_delay_46_7 <= io_A_Valid_4_delay_45_8;
    io_A_Valid_4_delay_47_6 <= io_A_Valid_4_delay_46_7;
    io_A_Valid_4_delay_48_5 <= io_A_Valid_4_delay_47_6;
    io_A_Valid_4_delay_49_4 <= io_A_Valid_4_delay_48_5;
    io_A_Valid_4_delay_50_3 <= io_A_Valid_4_delay_49_4;
    io_A_Valid_4_delay_51_2 <= io_A_Valid_4_delay_50_3;
    io_A_Valid_4_delay_52_1 <= io_A_Valid_4_delay_51_2;
    io_A_Valid_4_delay_53 <= io_A_Valid_4_delay_52_1;
    io_B_Valid_53_delay_1_3 <= io_B_Valid_53;
    io_B_Valid_53_delay_2_2 <= io_B_Valid_53_delay_1_3;
    io_B_Valid_53_delay_3_1 <= io_B_Valid_53_delay_2_2;
    io_B_Valid_53_delay_4 <= io_B_Valid_53_delay_3_1;
    io_A_Valid_4_delay_1_53 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_52 <= io_A_Valid_4_delay_1_53;
    io_A_Valid_4_delay_3_51 <= io_A_Valid_4_delay_2_52;
    io_A_Valid_4_delay_4_50 <= io_A_Valid_4_delay_3_51;
    io_A_Valid_4_delay_5_49 <= io_A_Valid_4_delay_4_50;
    io_A_Valid_4_delay_6_48 <= io_A_Valid_4_delay_5_49;
    io_A_Valid_4_delay_7_47 <= io_A_Valid_4_delay_6_48;
    io_A_Valid_4_delay_8_46 <= io_A_Valid_4_delay_7_47;
    io_A_Valid_4_delay_9_45 <= io_A_Valid_4_delay_8_46;
    io_A_Valid_4_delay_10_44 <= io_A_Valid_4_delay_9_45;
    io_A_Valid_4_delay_11_43 <= io_A_Valid_4_delay_10_44;
    io_A_Valid_4_delay_12_42 <= io_A_Valid_4_delay_11_43;
    io_A_Valid_4_delay_13_41 <= io_A_Valid_4_delay_12_42;
    io_A_Valid_4_delay_14_40 <= io_A_Valid_4_delay_13_41;
    io_A_Valid_4_delay_15_39 <= io_A_Valid_4_delay_14_40;
    io_A_Valid_4_delay_16_38 <= io_A_Valid_4_delay_15_39;
    io_A_Valid_4_delay_17_37 <= io_A_Valid_4_delay_16_38;
    io_A_Valid_4_delay_18_36 <= io_A_Valid_4_delay_17_37;
    io_A_Valid_4_delay_19_35 <= io_A_Valid_4_delay_18_36;
    io_A_Valid_4_delay_20_34 <= io_A_Valid_4_delay_19_35;
    io_A_Valid_4_delay_21_33 <= io_A_Valid_4_delay_20_34;
    io_A_Valid_4_delay_22_32 <= io_A_Valid_4_delay_21_33;
    io_A_Valid_4_delay_23_31 <= io_A_Valid_4_delay_22_32;
    io_A_Valid_4_delay_24_30 <= io_A_Valid_4_delay_23_31;
    io_A_Valid_4_delay_25_29 <= io_A_Valid_4_delay_24_30;
    io_A_Valid_4_delay_26_28 <= io_A_Valid_4_delay_25_29;
    io_A_Valid_4_delay_27_27 <= io_A_Valid_4_delay_26_28;
    io_A_Valid_4_delay_28_26 <= io_A_Valid_4_delay_27_27;
    io_A_Valid_4_delay_29_25 <= io_A_Valid_4_delay_28_26;
    io_A_Valid_4_delay_30_24 <= io_A_Valid_4_delay_29_25;
    io_A_Valid_4_delay_31_23 <= io_A_Valid_4_delay_30_24;
    io_A_Valid_4_delay_32_22 <= io_A_Valid_4_delay_31_23;
    io_A_Valid_4_delay_33_21 <= io_A_Valid_4_delay_32_22;
    io_A_Valid_4_delay_34_20 <= io_A_Valid_4_delay_33_21;
    io_A_Valid_4_delay_35_19 <= io_A_Valid_4_delay_34_20;
    io_A_Valid_4_delay_36_18 <= io_A_Valid_4_delay_35_19;
    io_A_Valid_4_delay_37_17 <= io_A_Valid_4_delay_36_18;
    io_A_Valid_4_delay_38_16 <= io_A_Valid_4_delay_37_17;
    io_A_Valid_4_delay_39_15 <= io_A_Valid_4_delay_38_16;
    io_A_Valid_4_delay_40_14 <= io_A_Valid_4_delay_39_15;
    io_A_Valid_4_delay_41_13 <= io_A_Valid_4_delay_40_14;
    io_A_Valid_4_delay_42_12 <= io_A_Valid_4_delay_41_13;
    io_A_Valid_4_delay_43_11 <= io_A_Valid_4_delay_42_12;
    io_A_Valid_4_delay_44_10 <= io_A_Valid_4_delay_43_11;
    io_A_Valid_4_delay_45_9 <= io_A_Valid_4_delay_44_10;
    io_A_Valid_4_delay_46_8 <= io_A_Valid_4_delay_45_9;
    io_A_Valid_4_delay_47_7 <= io_A_Valid_4_delay_46_8;
    io_A_Valid_4_delay_48_6 <= io_A_Valid_4_delay_47_7;
    io_A_Valid_4_delay_49_5 <= io_A_Valid_4_delay_48_6;
    io_A_Valid_4_delay_50_4 <= io_A_Valid_4_delay_49_5;
    io_A_Valid_4_delay_51_3 <= io_A_Valid_4_delay_50_4;
    io_A_Valid_4_delay_52_2 <= io_A_Valid_4_delay_51_3;
    io_A_Valid_4_delay_53_1 <= io_A_Valid_4_delay_52_2;
    io_A_Valid_4_delay_54 <= io_A_Valid_4_delay_53_1;
    io_B_Valid_54_delay_1_3 <= io_B_Valid_54;
    io_B_Valid_54_delay_2_2 <= io_B_Valid_54_delay_1_3;
    io_B_Valid_54_delay_3_1 <= io_B_Valid_54_delay_2_2;
    io_B_Valid_54_delay_4 <= io_B_Valid_54_delay_3_1;
    io_A_Valid_4_delay_1_54 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_53 <= io_A_Valid_4_delay_1_54;
    io_A_Valid_4_delay_3_52 <= io_A_Valid_4_delay_2_53;
    io_A_Valid_4_delay_4_51 <= io_A_Valid_4_delay_3_52;
    io_A_Valid_4_delay_5_50 <= io_A_Valid_4_delay_4_51;
    io_A_Valid_4_delay_6_49 <= io_A_Valid_4_delay_5_50;
    io_A_Valid_4_delay_7_48 <= io_A_Valid_4_delay_6_49;
    io_A_Valid_4_delay_8_47 <= io_A_Valid_4_delay_7_48;
    io_A_Valid_4_delay_9_46 <= io_A_Valid_4_delay_8_47;
    io_A_Valid_4_delay_10_45 <= io_A_Valid_4_delay_9_46;
    io_A_Valid_4_delay_11_44 <= io_A_Valid_4_delay_10_45;
    io_A_Valid_4_delay_12_43 <= io_A_Valid_4_delay_11_44;
    io_A_Valid_4_delay_13_42 <= io_A_Valid_4_delay_12_43;
    io_A_Valid_4_delay_14_41 <= io_A_Valid_4_delay_13_42;
    io_A_Valid_4_delay_15_40 <= io_A_Valid_4_delay_14_41;
    io_A_Valid_4_delay_16_39 <= io_A_Valid_4_delay_15_40;
    io_A_Valid_4_delay_17_38 <= io_A_Valid_4_delay_16_39;
    io_A_Valid_4_delay_18_37 <= io_A_Valid_4_delay_17_38;
    io_A_Valid_4_delay_19_36 <= io_A_Valid_4_delay_18_37;
    io_A_Valid_4_delay_20_35 <= io_A_Valid_4_delay_19_36;
    io_A_Valid_4_delay_21_34 <= io_A_Valid_4_delay_20_35;
    io_A_Valid_4_delay_22_33 <= io_A_Valid_4_delay_21_34;
    io_A_Valid_4_delay_23_32 <= io_A_Valid_4_delay_22_33;
    io_A_Valid_4_delay_24_31 <= io_A_Valid_4_delay_23_32;
    io_A_Valid_4_delay_25_30 <= io_A_Valid_4_delay_24_31;
    io_A_Valid_4_delay_26_29 <= io_A_Valid_4_delay_25_30;
    io_A_Valid_4_delay_27_28 <= io_A_Valid_4_delay_26_29;
    io_A_Valid_4_delay_28_27 <= io_A_Valid_4_delay_27_28;
    io_A_Valid_4_delay_29_26 <= io_A_Valid_4_delay_28_27;
    io_A_Valid_4_delay_30_25 <= io_A_Valid_4_delay_29_26;
    io_A_Valid_4_delay_31_24 <= io_A_Valid_4_delay_30_25;
    io_A_Valid_4_delay_32_23 <= io_A_Valid_4_delay_31_24;
    io_A_Valid_4_delay_33_22 <= io_A_Valid_4_delay_32_23;
    io_A_Valid_4_delay_34_21 <= io_A_Valid_4_delay_33_22;
    io_A_Valid_4_delay_35_20 <= io_A_Valid_4_delay_34_21;
    io_A_Valid_4_delay_36_19 <= io_A_Valid_4_delay_35_20;
    io_A_Valid_4_delay_37_18 <= io_A_Valid_4_delay_36_19;
    io_A_Valid_4_delay_38_17 <= io_A_Valid_4_delay_37_18;
    io_A_Valid_4_delay_39_16 <= io_A_Valid_4_delay_38_17;
    io_A_Valid_4_delay_40_15 <= io_A_Valid_4_delay_39_16;
    io_A_Valid_4_delay_41_14 <= io_A_Valid_4_delay_40_15;
    io_A_Valid_4_delay_42_13 <= io_A_Valid_4_delay_41_14;
    io_A_Valid_4_delay_43_12 <= io_A_Valid_4_delay_42_13;
    io_A_Valid_4_delay_44_11 <= io_A_Valid_4_delay_43_12;
    io_A_Valid_4_delay_45_10 <= io_A_Valid_4_delay_44_11;
    io_A_Valid_4_delay_46_9 <= io_A_Valid_4_delay_45_10;
    io_A_Valid_4_delay_47_8 <= io_A_Valid_4_delay_46_9;
    io_A_Valid_4_delay_48_7 <= io_A_Valid_4_delay_47_8;
    io_A_Valid_4_delay_49_6 <= io_A_Valid_4_delay_48_7;
    io_A_Valid_4_delay_50_5 <= io_A_Valid_4_delay_49_6;
    io_A_Valid_4_delay_51_4 <= io_A_Valid_4_delay_50_5;
    io_A_Valid_4_delay_52_3 <= io_A_Valid_4_delay_51_4;
    io_A_Valid_4_delay_53_2 <= io_A_Valid_4_delay_52_3;
    io_A_Valid_4_delay_54_1 <= io_A_Valid_4_delay_53_2;
    io_A_Valid_4_delay_55 <= io_A_Valid_4_delay_54_1;
    io_B_Valid_55_delay_1_3 <= io_B_Valid_55;
    io_B_Valid_55_delay_2_2 <= io_B_Valid_55_delay_1_3;
    io_B_Valid_55_delay_3_1 <= io_B_Valid_55_delay_2_2;
    io_B_Valid_55_delay_4 <= io_B_Valid_55_delay_3_1;
    io_A_Valid_4_delay_1_55 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_54 <= io_A_Valid_4_delay_1_55;
    io_A_Valid_4_delay_3_53 <= io_A_Valid_4_delay_2_54;
    io_A_Valid_4_delay_4_52 <= io_A_Valid_4_delay_3_53;
    io_A_Valid_4_delay_5_51 <= io_A_Valid_4_delay_4_52;
    io_A_Valid_4_delay_6_50 <= io_A_Valid_4_delay_5_51;
    io_A_Valid_4_delay_7_49 <= io_A_Valid_4_delay_6_50;
    io_A_Valid_4_delay_8_48 <= io_A_Valid_4_delay_7_49;
    io_A_Valid_4_delay_9_47 <= io_A_Valid_4_delay_8_48;
    io_A_Valid_4_delay_10_46 <= io_A_Valid_4_delay_9_47;
    io_A_Valid_4_delay_11_45 <= io_A_Valid_4_delay_10_46;
    io_A_Valid_4_delay_12_44 <= io_A_Valid_4_delay_11_45;
    io_A_Valid_4_delay_13_43 <= io_A_Valid_4_delay_12_44;
    io_A_Valid_4_delay_14_42 <= io_A_Valid_4_delay_13_43;
    io_A_Valid_4_delay_15_41 <= io_A_Valid_4_delay_14_42;
    io_A_Valid_4_delay_16_40 <= io_A_Valid_4_delay_15_41;
    io_A_Valid_4_delay_17_39 <= io_A_Valid_4_delay_16_40;
    io_A_Valid_4_delay_18_38 <= io_A_Valid_4_delay_17_39;
    io_A_Valid_4_delay_19_37 <= io_A_Valid_4_delay_18_38;
    io_A_Valid_4_delay_20_36 <= io_A_Valid_4_delay_19_37;
    io_A_Valid_4_delay_21_35 <= io_A_Valid_4_delay_20_36;
    io_A_Valid_4_delay_22_34 <= io_A_Valid_4_delay_21_35;
    io_A_Valid_4_delay_23_33 <= io_A_Valid_4_delay_22_34;
    io_A_Valid_4_delay_24_32 <= io_A_Valid_4_delay_23_33;
    io_A_Valid_4_delay_25_31 <= io_A_Valid_4_delay_24_32;
    io_A_Valid_4_delay_26_30 <= io_A_Valid_4_delay_25_31;
    io_A_Valid_4_delay_27_29 <= io_A_Valid_4_delay_26_30;
    io_A_Valid_4_delay_28_28 <= io_A_Valid_4_delay_27_29;
    io_A_Valid_4_delay_29_27 <= io_A_Valid_4_delay_28_28;
    io_A_Valid_4_delay_30_26 <= io_A_Valid_4_delay_29_27;
    io_A_Valid_4_delay_31_25 <= io_A_Valid_4_delay_30_26;
    io_A_Valid_4_delay_32_24 <= io_A_Valid_4_delay_31_25;
    io_A_Valid_4_delay_33_23 <= io_A_Valid_4_delay_32_24;
    io_A_Valid_4_delay_34_22 <= io_A_Valid_4_delay_33_23;
    io_A_Valid_4_delay_35_21 <= io_A_Valid_4_delay_34_22;
    io_A_Valid_4_delay_36_20 <= io_A_Valid_4_delay_35_21;
    io_A_Valid_4_delay_37_19 <= io_A_Valid_4_delay_36_20;
    io_A_Valid_4_delay_38_18 <= io_A_Valid_4_delay_37_19;
    io_A_Valid_4_delay_39_17 <= io_A_Valid_4_delay_38_18;
    io_A_Valid_4_delay_40_16 <= io_A_Valid_4_delay_39_17;
    io_A_Valid_4_delay_41_15 <= io_A_Valid_4_delay_40_16;
    io_A_Valid_4_delay_42_14 <= io_A_Valid_4_delay_41_15;
    io_A_Valid_4_delay_43_13 <= io_A_Valid_4_delay_42_14;
    io_A_Valid_4_delay_44_12 <= io_A_Valid_4_delay_43_13;
    io_A_Valid_4_delay_45_11 <= io_A_Valid_4_delay_44_12;
    io_A_Valid_4_delay_46_10 <= io_A_Valid_4_delay_45_11;
    io_A_Valid_4_delay_47_9 <= io_A_Valid_4_delay_46_10;
    io_A_Valid_4_delay_48_8 <= io_A_Valid_4_delay_47_9;
    io_A_Valid_4_delay_49_7 <= io_A_Valid_4_delay_48_8;
    io_A_Valid_4_delay_50_6 <= io_A_Valid_4_delay_49_7;
    io_A_Valid_4_delay_51_5 <= io_A_Valid_4_delay_50_6;
    io_A_Valid_4_delay_52_4 <= io_A_Valid_4_delay_51_5;
    io_A_Valid_4_delay_53_3 <= io_A_Valid_4_delay_52_4;
    io_A_Valid_4_delay_54_2 <= io_A_Valid_4_delay_53_3;
    io_A_Valid_4_delay_55_1 <= io_A_Valid_4_delay_54_2;
    io_A_Valid_4_delay_56 <= io_A_Valid_4_delay_55_1;
    io_B_Valid_56_delay_1_3 <= io_B_Valid_56;
    io_B_Valid_56_delay_2_2 <= io_B_Valid_56_delay_1_3;
    io_B_Valid_56_delay_3_1 <= io_B_Valid_56_delay_2_2;
    io_B_Valid_56_delay_4 <= io_B_Valid_56_delay_3_1;
    io_A_Valid_4_delay_1_56 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_55 <= io_A_Valid_4_delay_1_56;
    io_A_Valid_4_delay_3_54 <= io_A_Valid_4_delay_2_55;
    io_A_Valid_4_delay_4_53 <= io_A_Valid_4_delay_3_54;
    io_A_Valid_4_delay_5_52 <= io_A_Valid_4_delay_4_53;
    io_A_Valid_4_delay_6_51 <= io_A_Valid_4_delay_5_52;
    io_A_Valid_4_delay_7_50 <= io_A_Valid_4_delay_6_51;
    io_A_Valid_4_delay_8_49 <= io_A_Valid_4_delay_7_50;
    io_A_Valid_4_delay_9_48 <= io_A_Valid_4_delay_8_49;
    io_A_Valid_4_delay_10_47 <= io_A_Valid_4_delay_9_48;
    io_A_Valid_4_delay_11_46 <= io_A_Valid_4_delay_10_47;
    io_A_Valid_4_delay_12_45 <= io_A_Valid_4_delay_11_46;
    io_A_Valid_4_delay_13_44 <= io_A_Valid_4_delay_12_45;
    io_A_Valid_4_delay_14_43 <= io_A_Valid_4_delay_13_44;
    io_A_Valid_4_delay_15_42 <= io_A_Valid_4_delay_14_43;
    io_A_Valid_4_delay_16_41 <= io_A_Valid_4_delay_15_42;
    io_A_Valid_4_delay_17_40 <= io_A_Valid_4_delay_16_41;
    io_A_Valid_4_delay_18_39 <= io_A_Valid_4_delay_17_40;
    io_A_Valid_4_delay_19_38 <= io_A_Valid_4_delay_18_39;
    io_A_Valid_4_delay_20_37 <= io_A_Valid_4_delay_19_38;
    io_A_Valid_4_delay_21_36 <= io_A_Valid_4_delay_20_37;
    io_A_Valid_4_delay_22_35 <= io_A_Valid_4_delay_21_36;
    io_A_Valid_4_delay_23_34 <= io_A_Valid_4_delay_22_35;
    io_A_Valid_4_delay_24_33 <= io_A_Valid_4_delay_23_34;
    io_A_Valid_4_delay_25_32 <= io_A_Valid_4_delay_24_33;
    io_A_Valid_4_delay_26_31 <= io_A_Valid_4_delay_25_32;
    io_A_Valid_4_delay_27_30 <= io_A_Valid_4_delay_26_31;
    io_A_Valid_4_delay_28_29 <= io_A_Valid_4_delay_27_30;
    io_A_Valid_4_delay_29_28 <= io_A_Valid_4_delay_28_29;
    io_A_Valid_4_delay_30_27 <= io_A_Valid_4_delay_29_28;
    io_A_Valid_4_delay_31_26 <= io_A_Valid_4_delay_30_27;
    io_A_Valid_4_delay_32_25 <= io_A_Valid_4_delay_31_26;
    io_A_Valid_4_delay_33_24 <= io_A_Valid_4_delay_32_25;
    io_A_Valid_4_delay_34_23 <= io_A_Valid_4_delay_33_24;
    io_A_Valid_4_delay_35_22 <= io_A_Valid_4_delay_34_23;
    io_A_Valid_4_delay_36_21 <= io_A_Valid_4_delay_35_22;
    io_A_Valid_4_delay_37_20 <= io_A_Valid_4_delay_36_21;
    io_A_Valid_4_delay_38_19 <= io_A_Valid_4_delay_37_20;
    io_A_Valid_4_delay_39_18 <= io_A_Valid_4_delay_38_19;
    io_A_Valid_4_delay_40_17 <= io_A_Valid_4_delay_39_18;
    io_A_Valid_4_delay_41_16 <= io_A_Valid_4_delay_40_17;
    io_A_Valid_4_delay_42_15 <= io_A_Valid_4_delay_41_16;
    io_A_Valid_4_delay_43_14 <= io_A_Valid_4_delay_42_15;
    io_A_Valid_4_delay_44_13 <= io_A_Valid_4_delay_43_14;
    io_A_Valid_4_delay_45_12 <= io_A_Valid_4_delay_44_13;
    io_A_Valid_4_delay_46_11 <= io_A_Valid_4_delay_45_12;
    io_A_Valid_4_delay_47_10 <= io_A_Valid_4_delay_46_11;
    io_A_Valid_4_delay_48_9 <= io_A_Valid_4_delay_47_10;
    io_A_Valid_4_delay_49_8 <= io_A_Valid_4_delay_48_9;
    io_A_Valid_4_delay_50_7 <= io_A_Valid_4_delay_49_8;
    io_A_Valid_4_delay_51_6 <= io_A_Valid_4_delay_50_7;
    io_A_Valid_4_delay_52_5 <= io_A_Valid_4_delay_51_6;
    io_A_Valid_4_delay_53_4 <= io_A_Valid_4_delay_52_5;
    io_A_Valid_4_delay_54_3 <= io_A_Valid_4_delay_53_4;
    io_A_Valid_4_delay_55_2 <= io_A_Valid_4_delay_54_3;
    io_A_Valid_4_delay_56_1 <= io_A_Valid_4_delay_55_2;
    io_A_Valid_4_delay_57 <= io_A_Valid_4_delay_56_1;
    io_B_Valid_57_delay_1_3 <= io_B_Valid_57;
    io_B_Valid_57_delay_2_2 <= io_B_Valid_57_delay_1_3;
    io_B_Valid_57_delay_3_1 <= io_B_Valid_57_delay_2_2;
    io_B_Valid_57_delay_4 <= io_B_Valid_57_delay_3_1;
    io_A_Valid_4_delay_1_57 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_56 <= io_A_Valid_4_delay_1_57;
    io_A_Valid_4_delay_3_55 <= io_A_Valid_4_delay_2_56;
    io_A_Valid_4_delay_4_54 <= io_A_Valid_4_delay_3_55;
    io_A_Valid_4_delay_5_53 <= io_A_Valid_4_delay_4_54;
    io_A_Valid_4_delay_6_52 <= io_A_Valid_4_delay_5_53;
    io_A_Valid_4_delay_7_51 <= io_A_Valid_4_delay_6_52;
    io_A_Valid_4_delay_8_50 <= io_A_Valid_4_delay_7_51;
    io_A_Valid_4_delay_9_49 <= io_A_Valid_4_delay_8_50;
    io_A_Valid_4_delay_10_48 <= io_A_Valid_4_delay_9_49;
    io_A_Valid_4_delay_11_47 <= io_A_Valid_4_delay_10_48;
    io_A_Valid_4_delay_12_46 <= io_A_Valid_4_delay_11_47;
    io_A_Valid_4_delay_13_45 <= io_A_Valid_4_delay_12_46;
    io_A_Valid_4_delay_14_44 <= io_A_Valid_4_delay_13_45;
    io_A_Valid_4_delay_15_43 <= io_A_Valid_4_delay_14_44;
    io_A_Valid_4_delay_16_42 <= io_A_Valid_4_delay_15_43;
    io_A_Valid_4_delay_17_41 <= io_A_Valid_4_delay_16_42;
    io_A_Valid_4_delay_18_40 <= io_A_Valid_4_delay_17_41;
    io_A_Valid_4_delay_19_39 <= io_A_Valid_4_delay_18_40;
    io_A_Valid_4_delay_20_38 <= io_A_Valid_4_delay_19_39;
    io_A_Valid_4_delay_21_37 <= io_A_Valid_4_delay_20_38;
    io_A_Valid_4_delay_22_36 <= io_A_Valid_4_delay_21_37;
    io_A_Valid_4_delay_23_35 <= io_A_Valid_4_delay_22_36;
    io_A_Valid_4_delay_24_34 <= io_A_Valid_4_delay_23_35;
    io_A_Valid_4_delay_25_33 <= io_A_Valid_4_delay_24_34;
    io_A_Valid_4_delay_26_32 <= io_A_Valid_4_delay_25_33;
    io_A_Valid_4_delay_27_31 <= io_A_Valid_4_delay_26_32;
    io_A_Valid_4_delay_28_30 <= io_A_Valid_4_delay_27_31;
    io_A_Valid_4_delay_29_29 <= io_A_Valid_4_delay_28_30;
    io_A_Valid_4_delay_30_28 <= io_A_Valid_4_delay_29_29;
    io_A_Valid_4_delay_31_27 <= io_A_Valid_4_delay_30_28;
    io_A_Valid_4_delay_32_26 <= io_A_Valid_4_delay_31_27;
    io_A_Valid_4_delay_33_25 <= io_A_Valid_4_delay_32_26;
    io_A_Valid_4_delay_34_24 <= io_A_Valid_4_delay_33_25;
    io_A_Valid_4_delay_35_23 <= io_A_Valid_4_delay_34_24;
    io_A_Valid_4_delay_36_22 <= io_A_Valid_4_delay_35_23;
    io_A_Valid_4_delay_37_21 <= io_A_Valid_4_delay_36_22;
    io_A_Valid_4_delay_38_20 <= io_A_Valid_4_delay_37_21;
    io_A_Valid_4_delay_39_19 <= io_A_Valid_4_delay_38_20;
    io_A_Valid_4_delay_40_18 <= io_A_Valid_4_delay_39_19;
    io_A_Valid_4_delay_41_17 <= io_A_Valid_4_delay_40_18;
    io_A_Valid_4_delay_42_16 <= io_A_Valid_4_delay_41_17;
    io_A_Valid_4_delay_43_15 <= io_A_Valid_4_delay_42_16;
    io_A_Valid_4_delay_44_14 <= io_A_Valid_4_delay_43_15;
    io_A_Valid_4_delay_45_13 <= io_A_Valid_4_delay_44_14;
    io_A_Valid_4_delay_46_12 <= io_A_Valid_4_delay_45_13;
    io_A_Valid_4_delay_47_11 <= io_A_Valid_4_delay_46_12;
    io_A_Valid_4_delay_48_10 <= io_A_Valid_4_delay_47_11;
    io_A_Valid_4_delay_49_9 <= io_A_Valid_4_delay_48_10;
    io_A_Valid_4_delay_50_8 <= io_A_Valid_4_delay_49_9;
    io_A_Valid_4_delay_51_7 <= io_A_Valid_4_delay_50_8;
    io_A_Valid_4_delay_52_6 <= io_A_Valid_4_delay_51_7;
    io_A_Valid_4_delay_53_5 <= io_A_Valid_4_delay_52_6;
    io_A_Valid_4_delay_54_4 <= io_A_Valid_4_delay_53_5;
    io_A_Valid_4_delay_55_3 <= io_A_Valid_4_delay_54_4;
    io_A_Valid_4_delay_56_2 <= io_A_Valid_4_delay_55_3;
    io_A_Valid_4_delay_57_1 <= io_A_Valid_4_delay_56_2;
    io_A_Valid_4_delay_58 <= io_A_Valid_4_delay_57_1;
    io_B_Valid_58_delay_1_3 <= io_B_Valid_58;
    io_B_Valid_58_delay_2_2 <= io_B_Valid_58_delay_1_3;
    io_B_Valid_58_delay_3_1 <= io_B_Valid_58_delay_2_2;
    io_B_Valid_58_delay_4 <= io_B_Valid_58_delay_3_1;
    io_A_Valid_4_delay_1_58 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_57 <= io_A_Valid_4_delay_1_58;
    io_A_Valid_4_delay_3_56 <= io_A_Valid_4_delay_2_57;
    io_A_Valid_4_delay_4_55 <= io_A_Valid_4_delay_3_56;
    io_A_Valid_4_delay_5_54 <= io_A_Valid_4_delay_4_55;
    io_A_Valid_4_delay_6_53 <= io_A_Valid_4_delay_5_54;
    io_A_Valid_4_delay_7_52 <= io_A_Valid_4_delay_6_53;
    io_A_Valid_4_delay_8_51 <= io_A_Valid_4_delay_7_52;
    io_A_Valid_4_delay_9_50 <= io_A_Valid_4_delay_8_51;
    io_A_Valid_4_delay_10_49 <= io_A_Valid_4_delay_9_50;
    io_A_Valid_4_delay_11_48 <= io_A_Valid_4_delay_10_49;
    io_A_Valid_4_delay_12_47 <= io_A_Valid_4_delay_11_48;
    io_A_Valid_4_delay_13_46 <= io_A_Valid_4_delay_12_47;
    io_A_Valid_4_delay_14_45 <= io_A_Valid_4_delay_13_46;
    io_A_Valid_4_delay_15_44 <= io_A_Valid_4_delay_14_45;
    io_A_Valid_4_delay_16_43 <= io_A_Valid_4_delay_15_44;
    io_A_Valid_4_delay_17_42 <= io_A_Valid_4_delay_16_43;
    io_A_Valid_4_delay_18_41 <= io_A_Valid_4_delay_17_42;
    io_A_Valid_4_delay_19_40 <= io_A_Valid_4_delay_18_41;
    io_A_Valid_4_delay_20_39 <= io_A_Valid_4_delay_19_40;
    io_A_Valid_4_delay_21_38 <= io_A_Valid_4_delay_20_39;
    io_A_Valid_4_delay_22_37 <= io_A_Valid_4_delay_21_38;
    io_A_Valid_4_delay_23_36 <= io_A_Valid_4_delay_22_37;
    io_A_Valid_4_delay_24_35 <= io_A_Valid_4_delay_23_36;
    io_A_Valid_4_delay_25_34 <= io_A_Valid_4_delay_24_35;
    io_A_Valid_4_delay_26_33 <= io_A_Valid_4_delay_25_34;
    io_A_Valid_4_delay_27_32 <= io_A_Valid_4_delay_26_33;
    io_A_Valid_4_delay_28_31 <= io_A_Valid_4_delay_27_32;
    io_A_Valid_4_delay_29_30 <= io_A_Valid_4_delay_28_31;
    io_A_Valid_4_delay_30_29 <= io_A_Valid_4_delay_29_30;
    io_A_Valid_4_delay_31_28 <= io_A_Valid_4_delay_30_29;
    io_A_Valid_4_delay_32_27 <= io_A_Valid_4_delay_31_28;
    io_A_Valid_4_delay_33_26 <= io_A_Valid_4_delay_32_27;
    io_A_Valid_4_delay_34_25 <= io_A_Valid_4_delay_33_26;
    io_A_Valid_4_delay_35_24 <= io_A_Valid_4_delay_34_25;
    io_A_Valid_4_delay_36_23 <= io_A_Valid_4_delay_35_24;
    io_A_Valid_4_delay_37_22 <= io_A_Valid_4_delay_36_23;
    io_A_Valid_4_delay_38_21 <= io_A_Valid_4_delay_37_22;
    io_A_Valid_4_delay_39_20 <= io_A_Valid_4_delay_38_21;
    io_A_Valid_4_delay_40_19 <= io_A_Valid_4_delay_39_20;
    io_A_Valid_4_delay_41_18 <= io_A_Valid_4_delay_40_19;
    io_A_Valid_4_delay_42_17 <= io_A_Valid_4_delay_41_18;
    io_A_Valid_4_delay_43_16 <= io_A_Valid_4_delay_42_17;
    io_A_Valid_4_delay_44_15 <= io_A_Valid_4_delay_43_16;
    io_A_Valid_4_delay_45_14 <= io_A_Valid_4_delay_44_15;
    io_A_Valid_4_delay_46_13 <= io_A_Valid_4_delay_45_14;
    io_A_Valid_4_delay_47_12 <= io_A_Valid_4_delay_46_13;
    io_A_Valid_4_delay_48_11 <= io_A_Valid_4_delay_47_12;
    io_A_Valid_4_delay_49_10 <= io_A_Valid_4_delay_48_11;
    io_A_Valid_4_delay_50_9 <= io_A_Valid_4_delay_49_10;
    io_A_Valid_4_delay_51_8 <= io_A_Valid_4_delay_50_9;
    io_A_Valid_4_delay_52_7 <= io_A_Valid_4_delay_51_8;
    io_A_Valid_4_delay_53_6 <= io_A_Valid_4_delay_52_7;
    io_A_Valid_4_delay_54_5 <= io_A_Valid_4_delay_53_6;
    io_A_Valid_4_delay_55_4 <= io_A_Valid_4_delay_54_5;
    io_A_Valid_4_delay_56_3 <= io_A_Valid_4_delay_55_4;
    io_A_Valid_4_delay_57_2 <= io_A_Valid_4_delay_56_3;
    io_A_Valid_4_delay_58_1 <= io_A_Valid_4_delay_57_2;
    io_A_Valid_4_delay_59 <= io_A_Valid_4_delay_58_1;
    io_B_Valid_59_delay_1_3 <= io_B_Valid_59;
    io_B_Valid_59_delay_2_2 <= io_B_Valid_59_delay_1_3;
    io_B_Valid_59_delay_3_1 <= io_B_Valid_59_delay_2_2;
    io_B_Valid_59_delay_4 <= io_B_Valid_59_delay_3_1;
    io_A_Valid_4_delay_1_59 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_58 <= io_A_Valid_4_delay_1_59;
    io_A_Valid_4_delay_3_57 <= io_A_Valid_4_delay_2_58;
    io_A_Valid_4_delay_4_56 <= io_A_Valid_4_delay_3_57;
    io_A_Valid_4_delay_5_55 <= io_A_Valid_4_delay_4_56;
    io_A_Valid_4_delay_6_54 <= io_A_Valid_4_delay_5_55;
    io_A_Valid_4_delay_7_53 <= io_A_Valid_4_delay_6_54;
    io_A_Valid_4_delay_8_52 <= io_A_Valid_4_delay_7_53;
    io_A_Valid_4_delay_9_51 <= io_A_Valid_4_delay_8_52;
    io_A_Valid_4_delay_10_50 <= io_A_Valid_4_delay_9_51;
    io_A_Valid_4_delay_11_49 <= io_A_Valid_4_delay_10_50;
    io_A_Valid_4_delay_12_48 <= io_A_Valid_4_delay_11_49;
    io_A_Valid_4_delay_13_47 <= io_A_Valid_4_delay_12_48;
    io_A_Valid_4_delay_14_46 <= io_A_Valid_4_delay_13_47;
    io_A_Valid_4_delay_15_45 <= io_A_Valid_4_delay_14_46;
    io_A_Valid_4_delay_16_44 <= io_A_Valid_4_delay_15_45;
    io_A_Valid_4_delay_17_43 <= io_A_Valid_4_delay_16_44;
    io_A_Valid_4_delay_18_42 <= io_A_Valid_4_delay_17_43;
    io_A_Valid_4_delay_19_41 <= io_A_Valid_4_delay_18_42;
    io_A_Valid_4_delay_20_40 <= io_A_Valid_4_delay_19_41;
    io_A_Valid_4_delay_21_39 <= io_A_Valid_4_delay_20_40;
    io_A_Valid_4_delay_22_38 <= io_A_Valid_4_delay_21_39;
    io_A_Valid_4_delay_23_37 <= io_A_Valid_4_delay_22_38;
    io_A_Valid_4_delay_24_36 <= io_A_Valid_4_delay_23_37;
    io_A_Valid_4_delay_25_35 <= io_A_Valid_4_delay_24_36;
    io_A_Valid_4_delay_26_34 <= io_A_Valid_4_delay_25_35;
    io_A_Valid_4_delay_27_33 <= io_A_Valid_4_delay_26_34;
    io_A_Valid_4_delay_28_32 <= io_A_Valid_4_delay_27_33;
    io_A_Valid_4_delay_29_31 <= io_A_Valid_4_delay_28_32;
    io_A_Valid_4_delay_30_30 <= io_A_Valid_4_delay_29_31;
    io_A_Valid_4_delay_31_29 <= io_A_Valid_4_delay_30_30;
    io_A_Valid_4_delay_32_28 <= io_A_Valid_4_delay_31_29;
    io_A_Valid_4_delay_33_27 <= io_A_Valid_4_delay_32_28;
    io_A_Valid_4_delay_34_26 <= io_A_Valid_4_delay_33_27;
    io_A_Valid_4_delay_35_25 <= io_A_Valid_4_delay_34_26;
    io_A_Valid_4_delay_36_24 <= io_A_Valid_4_delay_35_25;
    io_A_Valid_4_delay_37_23 <= io_A_Valid_4_delay_36_24;
    io_A_Valid_4_delay_38_22 <= io_A_Valid_4_delay_37_23;
    io_A_Valid_4_delay_39_21 <= io_A_Valid_4_delay_38_22;
    io_A_Valid_4_delay_40_20 <= io_A_Valid_4_delay_39_21;
    io_A_Valid_4_delay_41_19 <= io_A_Valid_4_delay_40_20;
    io_A_Valid_4_delay_42_18 <= io_A_Valid_4_delay_41_19;
    io_A_Valid_4_delay_43_17 <= io_A_Valid_4_delay_42_18;
    io_A_Valid_4_delay_44_16 <= io_A_Valid_4_delay_43_17;
    io_A_Valid_4_delay_45_15 <= io_A_Valid_4_delay_44_16;
    io_A_Valid_4_delay_46_14 <= io_A_Valid_4_delay_45_15;
    io_A_Valid_4_delay_47_13 <= io_A_Valid_4_delay_46_14;
    io_A_Valid_4_delay_48_12 <= io_A_Valid_4_delay_47_13;
    io_A_Valid_4_delay_49_11 <= io_A_Valid_4_delay_48_12;
    io_A_Valid_4_delay_50_10 <= io_A_Valid_4_delay_49_11;
    io_A_Valid_4_delay_51_9 <= io_A_Valid_4_delay_50_10;
    io_A_Valid_4_delay_52_8 <= io_A_Valid_4_delay_51_9;
    io_A_Valid_4_delay_53_7 <= io_A_Valid_4_delay_52_8;
    io_A_Valid_4_delay_54_6 <= io_A_Valid_4_delay_53_7;
    io_A_Valid_4_delay_55_5 <= io_A_Valid_4_delay_54_6;
    io_A_Valid_4_delay_56_4 <= io_A_Valid_4_delay_55_5;
    io_A_Valid_4_delay_57_3 <= io_A_Valid_4_delay_56_4;
    io_A_Valid_4_delay_58_2 <= io_A_Valid_4_delay_57_3;
    io_A_Valid_4_delay_59_1 <= io_A_Valid_4_delay_58_2;
    io_A_Valid_4_delay_60 <= io_A_Valid_4_delay_59_1;
    io_B_Valid_60_delay_1_3 <= io_B_Valid_60;
    io_B_Valid_60_delay_2_2 <= io_B_Valid_60_delay_1_3;
    io_B_Valid_60_delay_3_1 <= io_B_Valid_60_delay_2_2;
    io_B_Valid_60_delay_4 <= io_B_Valid_60_delay_3_1;
    io_A_Valid_4_delay_1_60 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_59 <= io_A_Valid_4_delay_1_60;
    io_A_Valid_4_delay_3_58 <= io_A_Valid_4_delay_2_59;
    io_A_Valid_4_delay_4_57 <= io_A_Valid_4_delay_3_58;
    io_A_Valid_4_delay_5_56 <= io_A_Valid_4_delay_4_57;
    io_A_Valid_4_delay_6_55 <= io_A_Valid_4_delay_5_56;
    io_A_Valid_4_delay_7_54 <= io_A_Valid_4_delay_6_55;
    io_A_Valid_4_delay_8_53 <= io_A_Valid_4_delay_7_54;
    io_A_Valid_4_delay_9_52 <= io_A_Valid_4_delay_8_53;
    io_A_Valid_4_delay_10_51 <= io_A_Valid_4_delay_9_52;
    io_A_Valid_4_delay_11_50 <= io_A_Valid_4_delay_10_51;
    io_A_Valid_4_delay_12_49 <= io_A_Valid_4_delay_11_50;
    io_A_Valid_4_delay_13_48 <= io_A_Valid_4_delay_12_49;
    io_A_Valid_4_delay_14_47 <= io_A_Valid_4_delay_13_48;
    io_A_Valid_4_delay_15_46 <= io_A_Valid_4_delay_14_47;
    io_A_Valid_4_delay_16_45 <= io_A_Valid_4_delay_15_46;
    io_A_Valid_4_delay_17_44 <= io_A_Valid_4_delay_16_45;
    io_A_Valid_4_delay_18_43 <= io_A_Valid_4_delay_17_44;
    io_A_Valid_4_delay_19_42 <= io_A_Valid_4_delay_18_43;
    io_A_Valid_4_delay_20_41 <= io_A_Valid_4_delay_19_42;
    io_A_Valid_4_delay_21_40 <= io_A_Valid_4_delay_20_41;
    io_A_Valid_4_delay_22_39 <= io_A_Valid_4_delay_21_40;
    io_A_Valid_4_delay_23_38 <= io_A_Valid_4_delay_22_39;
    io_A_Valid_4_delay_24_37 <= io_A_Valid_4_delay_23_38;
    io_A_Valid_4_delay_25_36 <= io_A_Valid_4_delay_24_37;
    io_A_Valid_4_delay_26_35 <= io_A_Valid_4_delay_25_36;
    io_A_Valid_4_delay_27_34 <= io_A_Valid_4_delay_26_35;
    io_A_Valid_4_delay_28_33 <= io_A_Valid_4_delay_27_34;
    io_A_Valid_4_delay_29_32 <= io_A_Valid_4_delay_28_33;
    io_A_Valid_4_delay_30_31 <= io_A_Valid_4_delay_29_32;
    io_A_Valid_4_delay_31_30 <= io_A_Valid_4_delay_30_31;
    io_A_Valid_4_delay_32_29 <= io_A_Valid_4_delay_31_30;
    io_A_Valid_4_delay_33_28 <= io_A_Valid_4_delay_32_29;
    io_A_Valid_4_delay_34_27 <= io_A_Valid_4_delay_33_28;
    io_A_Valid_4_delay_35_26 <= io_A_Valid_4_delay_34_27;
    io_A_Valid_4_delay_36_25 <= io_A_Valid_4_delay_35_26;
    io_A_Valid_4_delay_37_24 <= io_A_Valid_4_delay_36_25;
    io_A_Valid_4_delay_38_23 <= io_A_Valid_4_delay_37_24;
    io_A_Valid_4_delay_39_22 <= io_A_Valid_4_delay_38_23;
    io_A_Valid_4_delay_40_21 <= io_A_Valid_4_delay_39_22;
    io_A_Valid_4_delay_41_20 <= io_A_Valid_4_delay_40_21;
    io_A_Valid_4_delay_42_19 <= io_A_Valid_4_delay_41_20;
    io_A_Valid_4_delay_43_18 <= io_A_Valid_4_delay_42_19;
    io_A_Valid_4_delay_44_17 <= io_A_Valid_4_delay_43_18;
    io_A_Valid_4_delay_45_16 <= io_A_Valid_4_delay_44_17;
    io_A_Valid_4_delay_46_15 <= io_A_Valid_4_delay_45_16;
    io_A_Valid_4_delay_47_14 <= io_A_Valid_4_delay_46_15;
    io_A_Valid_4_delay_48_13 <= io_A_Valid_4_delay_47_14;
    io_A_Valid_4_delay_49_12 <= io_A_Valid_4_delay_48_13;
    io_A_Valid_4_delay_50_11 <= io_A_Valid_4_delay_49_12;
    io_A_Valid_4_delay_51_10 <= io_A_Valid_4_delay_50_11;
    io_A_Valid_4_delay_52_9 <= io_A_Valid_4_delay_51_10;
    io_A_Valid_4_delay_53_8 <= io_A_Valid_4_delay_52_9;
    io_A_Valid_4_delay_54_7 <= io_A_Valid_4_delay_53_8;
    io_A_Valid_4_delay_55_6 <= io_A_Valid_4_delay_54_7;
    io_A_Valid_4_delay_56_5 <= io_A_Valid_4_delay_55_6;
    io_A_Valid_4_delay_57_4 <= io_A_Valid_4_delay_56_5;
    io_A_Valid_4_delay_58_3 <= io_A_Valid_4_delay_57_4;
    io_A_Valid_4_delay_59_2 <= io_A_Valid_4_delay_58_3;
    io_A_Valid_4_delay_60_1 <= io_A_Valid_4_delay_59_2;
    io_A_Valid_4_delay_61 <= io_A_Valid_4_delay_60_1;
    io_B_Valid_61_delay_1_3 <= io_B_Valid_61;
    io_B_Valid_61_delay_2_2 <= io_B_Valid_61_delay_1_3;
    io_B_Valid_61_delay_3_1 <= io_B_Valid_61_delay_2_2;
    io_B_Valid_61_delay_4 <= io_B_Valid_61_delay_3_1;
    io_A_Valid_4_delay_1_61 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_60 <= io_A_Valid_4_delay_1_61;
    io_A_Valid_4_delay_3_59 <= io_A_Valid_4_delay_2_60;
    io_A_Valid_4_delay_4_58 <= io_A_Valid_4_delay_3_59;
    io_A_Valid_4_delay_5_57 <= io_A_Valid_4_delay_4_58;
    io_A_Valid_4_delay_6_56 <= io_A_Valid_4_delay_5_57;
    io_A_Valid_4_delay_7_55 <= io_A_Valid_4_delay_6_56;
    io_A_Valid_4_delay_8_54 <= io_A_Valid_4_delay_7_55;
    io_A_Valid_4_delay_9_53 <= io_A_Valid_4_delay_8_54;
    io_A_Valid_4_delay_10_52 <= io_A_Valid_4_delay_9_53;
    io_A_Valid_4_delay_11_51 <= io_A_Valid_4_delay_10_52;
    io_A_Valid_4_delay_12_50 <= io_A_Valid_4_delay_11_51;
    io_A_Valid_4_delay_13_49 <= io_A_Valid_4_delay_12_50;
    io_A_Valid_4_delay_14_48 <= io_A_Valid_4_delay_13_49;
    io_A_Valid_4_delay_15_47 <= io_A_Valid_4_delay_14_48;
    io_A_Valid_4_delay_16_46 <= io_A_Valid_4_delay_15_47;
    io_A_Valid_4_delay_17_45 <= io_A_Valid_4_delay_16_46;
    io_A_Valid_4_delay_18_44 <= io_A_Valid_4_delay_17_45;
    io_A_Valid_4_delay_19_43 <= io_A_Valid_4_delay_18_44;
    io_A_Valid_4_delay_20_42 <= io_A_Valid_4_delay_19_43;
    io_A_Valid_4_delay_21_41 <= io_A_Valid_4_delay_20_42;
    io_A_Valid_4_delay_22_40 <= io_A_Valid_4_delay_21_41;
    io_A_Valid_4_delay_23_39 <= io_A_Valid_4_delay_22_40;
    io_A_Valid_4_delay_24_38 <= io_A_Valid_4_delay_23_39;
    io_A_Valid_4_delay_25_37 <= io_A_Valid_4_delay_24_38;
    io_A_Valid_4_delay_26_36 <= io_A_Valid_4_delay_25_37;
    io_A_Valid_4_delay_27_35 <= io_A_Valid_4_delay_26_36;
    io_A_Valid_4_delay_28_34 <= io_A_Valid_4_delay_27_35;
    io_A_Valid_4_delay_29_33 <= io_A_Valid_4_delay_28_34;
    io_A_Valid_4_delay_30_32 <= io_A_Valid_4_delay_29_33;
    io_A_Valid_4_delay_31_31 <= io_A_Valid_4_delay_30_32;
    io_A_Valid_4_delay_32_30 <= io_A_Valid_4_delay_31_31;
    io_A_Valid_4_delay_33_29 <= io_A_Valid_4_delay_32_30;
    io_A_Valid_4_delay_34_28 <= io_A_Valid_4_delay_33_29;
    io_A_Valid_4_delay_35_27 <= io_A_Valid_4_delay_34_28;
    io_A_Valid_4_delay_36_26 <= io_A_Valid_4_delay_35_27;
    io_A_Valid_4_delay_37_25 <= io_A_Valid_4_delay_36_26;
    io_A_Valid_4_delay_38_24 <= io_A_Valid_4_delay_37_25;
    io_A_Valid_4_delay_39_23 <= io_A_Valid_4_delay_38_24;
    io_A_Valid_4_delay_40_22 <= io_A_Valid_4_delay_39_23;
    io_A_Valid_4_delay_41_21 <= io_A_Valid_4_delay_40_22;
    io_A_Valid_4_delay_42_20 <= io_A_Valid_4_delay_41_21;
    io_A_Valid_4_delay_43_19 <= io_A_Valid_4_delay_42_20;
    io_A_Valid_4_delay_44_18 <= io_A_Valid_4_delay_43_19;
    io_A_Valid_4_delay_45_17 <= io_A_Valid_4_delay_44_18;
    io_A_Valid_4_delay_46_16 <= io_A_Valid_4_delay_45_17;
    io_A_Valid_4_delay_47_15 <= io_A_Valid_4_delay_46_16;
    io_A_Valid_4_delay_48_14 <= io_A_Valid_4_delay_47_15;
    io_A_Valid_4_delay_49_13 <= io_A_Valid_4_delay_48_14;
    io_A_Valid_4_delay_50_12 <= io_A_Valid_4_delay_49_13;
    io_A_Valid_4_delay_51_11 <= io_A_Valid_4_delay_50_12;
    io_A_Valid_4_delay_52_10 <= io_A_Valid_4_delay_51_11;
    io_A_Valid_4_delay_53_9 <= io_A_Valid_4_delay_52_10;
    io_A_Valid_4_delay_54_8 <= io_A_Valid_4_delay_53_9;
    io_A_Valid_4_delay_55_7 <= io_A_Valid_4_delay_54_8;
    io_A_Valid_4_delay_56_6 <= io_A_Valid_4_delay_55_7;
    io_A_Valid_4_delay_57_5 <= io_A_Valid_4_delay_56_6;
    io_A_Valid_4_delay_58_4 <= io_A_Valid_4_delay_57_5;
    io_A_Valid_4_delay_59_3 <= io_A_Valid_4_delay_58_4;
    io_A_Valid_4_delay_60_2 <= io_A_Valid_4_delay_59_3;
    io_A_Valid_4_delay_61_1 <= io_A_Valid_4_delay_60_2;
    io_A_Valid_4_delay_62 <= io_A_Valid_4_delay_61_1;
    io_B_Valid_62_delay_1_3 <= io_B_Valid_62;
    io_B_Valid_62_delay_2_2 <= io_B_Valid_62_delay_1_3;
    io_B_Valid_62_delay_3_1 <= io_B_Valid_62_delay_2_2;
    io_B_Valid_62_delay_4 <= io_B_Valid_62_delay_3_1;
    io_A_Valid_4_delay_1_62 <= io_A_Valid_4;
    io_A_Valid_4_delay_2_61 <= io_A_Valid_4_delay_1_62;
    io_A_Valid_4_delay_3_60 <= io_A_Valid_4_delay_2_61;
    io_A_Valid_4_delay_4_59 <= io_A_Valid_4_delay_3_60;
    io_A_Valid_4_delay_5_58 <= io_A_Valid_4_delay_4_59;
    io_A_Valid_4_delay_6_57 <= io_A_Valid_4_delay_5_58;
    io_A_Valid_4_delay_7_56 <= io_A_Valid_4_delay_6_57;
    io_A_Valid_4_delay_8_55 <= io_A_Valid_4_delay_7_56;
    io_A_Valid_4_delay_9_54 <= io_A_Valid_4_delay_8_55;
    io_A_Valid_4_delay_10_53 <= io_A_Valid_4_delay_9_54;
    io_A_Valid_4_delay_11_52 <= io_A_Valid_4_delay_10_53;
    io_A_Valid_4_delay_12_51 <= io_A_Valid_4_delay_11_52;
    io_A_Valid_4_delay_13_50 <= io_A_Valid_4_delay_12_51;
    io_A_Valid_4_delay_14_49 <= io_A_Valid_4_delay_13_50;
    io_A_Valid_4_delay_15_48 <= io_A_Valid_4_delay_14_49;
    io_A_Valid_4_delay_16_47 <= io_A_Valid_4_delay_15_48;
    io_A_Valid_4_delay_17_46 <= io_A_Valid_4_delay_16_47;
    io_A_Valid_4_delay_18_45 <= io_A_Valid_4_delay_17_46;
    io_A_Valid_4_delay_19_44 <= io_A_Valid_4_delay_18_45;
    io_A_Valid_4_delay_20_43 <= io_A_Valid_4_delay_19_44;
    io_A_Valid_4_delay_21_42 <= io_A_Valid_4_delay_20_43;
    io_A_Valid_4_delay_22_41 <= io_A_Valid_4_delay_21_42;
    io_A_Valid_4_delay_23_40 <= io_A_Valid_4_delay_22_41;
    io_A_Valid_4_delay_24_39 <= io_A_Valid_4_delay_23_40;
    io_A_Valid_4_delay_25_38 <= io_A_Valid_4_delay_24_39;
    io_A_Valid_4_delay_26_37 <= io_A_Valid_4_delay_25_38;
    io_A_Valid_4_delay_27_36 <= io_A_Valid_4_delay_26_37;
    io_A_Valid_4_delay_28_35 <= io_A_Valid_4_delay_27_36;
    io_A_Valid_4_delay_29_34 <= io_A_Valid_4_delay_28_35;
    io_A_Valid_4_delay_30_33 <= io_A_Valid_4_delay_29_34;
    io_A_Valid_4_delay_31_32 <= io_A_Valid_4_delay_30_33;
    io_A_Valid_4_delay_32_31 <= io_A_Valid_4_delay_31_32;
    io_A_Valid_4_delay_33_30 <= io_A_Valid_4_delay_32_31;
    io_A_Valid_4_delay_34_29 <= io_A_Valid_4_delay_33_30;
    io_A_Valid_4_delay_35_28 <= io_A_Valid_4_delay_34_29;
    io_A_Valid_4_delay_36_27 <= io_A_Valid_4_delay_35_28;
    io_A_Valid_4_delay_37_26 <= io_A_Valid_4_delay_36_27;
    io_A_Valid_4_delay_38_25 <= io_A_Valid_4_delay_37_26;
    io_A_Valid_4_delay_39_24 <= io_A_Valid_4_delay_38_25;
    io_A_Valid_4_delay_40_23 <= io_A_Valid_4_delay_39_24;
    io_A_Valid_4_delay_41_22 <= io_A_Valid_4_delay_40_23;
    io_A_Valid_4_delay_42_21 <= io_A_Valid_4_delay_41_22;
    io_A_Valid_4_delay_43_20 <= io_A_Valid_4_delay_42_21;
    io_A_Valid_4_delay_44_19 <= io_A_Valid_4_delay_43_20;
    io_A_Valid_4_delay_45_18 <= io_A_Valid_4_delay_44_19;
    io_A_Valid_4_delay_46_17 <= io_A_Valid_4_delay_45_18;
    io_A_Valid_4_delay_47_16 <= io_A_Valid_4_delay_46_17;
    io_A_Valid_4_delay_48_15 <= io_A_Valid_4_delay_47_16;
    io_A_Valid_4_delay_49_14 <= io_A_Valid_4_delay_48_15;
    io_A_Valid_4_delay_50_13 <= io_A_Valid_4_delay_49_14;
    io_A_Valid_4_delay_51_12 <= io_A_Valid_4_delay_50_13;
    io_A_Valid_4_delay_52_11 <= io_A_Valid_4_delay_51_12;
    io_A_Valid_4_delay_53_10 <= io_A_Valid_4_delay_52_11;
    io_A_Valid_4_delay_54_9 <= io_A_Valid_4_delay_53_10;
    io_A_Valid_4_delay_55_8 <= io_A_Valid_4_delay_54_9;
    io_A_Valid_4_delay_56_7 <= io_A_Valid_4_delay_55_8;
    io_A_Valid_4_delay_57_6 <= io_A_Valid_4_delay_56_7;
    io_A_Valid_4_delay_58_5 <= io_A_Valid_4_delay_57_6;
    io_A_Valid_4_delay_59_4 <= io_A_Valid_4_delay_58_5;
    io_A_Valid_4_delay_60_3 <= io_A_Valid_4_delay_59_4;
    io_A_Valid_4_delay_61_2 <= io_A_Valid_4_delay_60_3;
    io_A_Valid_4_delay_62_1 <= io_A_Valid_4_delay_61_2;
    io_A_Valid_4_delay_63 <= io_A_Valid_4_delay_62_1;
    io_B_Valid_63_delay_1_3 <= io_B_Valid_63;
    io_B_Valid_63_delay_2_2 <= io_B_Valid_63_delay_1_3;
    io_B_Valid_63_delay_3_1 <= io_B_Valid_63_delay_2_2;
    io_B_Valid_63_delay_4 <= io_B_Valid_63_delay_3_1;
    io_B_Valid_0_delay_1_4 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_3 <= io_B_Valid_0_delay_1_4;
    io_B_Valid_0_delay_3_2 <= io_B_Valid_0_delay_2_3;
    io_B_Valid_0_delay_4_1 <= io_B_Valid_0_delay_3_2;
    io_B_Valid_0_delay_5 <= io_B_Valid_0_delay_4_1;
    io_A_Valid_5_delay_1 <= io_A_Valid_5;
    io_B_Valid_1_delay_1_4 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_3 <= io_B_Valid_1_delay_1_4;
    io_B_Valid_1_delay_3_2 <= io_B_Valid_1_delay_2_3;
    io_B_Valid_1_delay_4_1 <= io_B_Valid_1_delay_3_2;
    io_B_Valid_1_delay_5 <= io_B_Valid_1_delay_4_1;
    io_A_Valid_5_delay_1_1 <= io_A_Valid_5;
    io_A_Valid_5_delay_2 <= io_A_Valid_5_delay_1_1;
    io_B_Valid_2_delay_1_4 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_3 <= io_B_Valid_2_delay_1_4;
    io_B_Valid_2_delay_3_2 <= io_B_Valid_2_delay_2_3;
    io_B_Valid_2_delay_4_1 <= io_B_Valid_2_delay_3_2;
    io_B_Valid_2_delay_5 <= io_B_Valid_2_delay_4_1;
    io_A_Valid_5_delay_1_2 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_1 <= io_A_Valid_5_delay_1_2;
    io_A_Valid_5_delay_3 <= io_A_Valid_5_delay_2_1;
    io_B_Valid_3_delay_1_4 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_3 <= io_B_Valid_3_delay_1_4;
    io_B_Valid_3_delay_3_2 <= io_B_Valid_3_delay_2_3;
    io_B_Valid_3_delay_4_1 <= io_B_Valid_3_delay_3_2;
    io_B_Valid_3_delay_5 <= io_B_Valid_3_delay_4_1;
    io_A_Valid_5_delay_1_3 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_2 <= io_A_Valid_5_delay_1_3;
    io_A_Valid_5_delay_3_1 <= io_A_Valid_5_delay_2_2;
    io_A_Valid_5_delay_4 <= io_A_Valid_5_delay_3_1;
    io_B_Valid_4_delay_1_4 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_3 <= io_B_Valid_4_delay_1_4;
    io_B_Valid_4_delay_3_2 <= io_B_Valid_4_delay_2_3;
    io_B_Valid_4_delay_4_1 <= io_B_Valid_4_delay_3_2;
    io_B_Valid_4_delay_5 <= io_B_Valid_4_delay_4_1;
    io_A_Valid_5_delay_1_4 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_3 <= io_A_Valid_5_delay_1_4;
    io_A_Valid_5_delay_3_2 <= io_A_Valid_5_delay_2_3;
    io_A_Valid_5_delay_4_1 <= io_A_Valid_5_delay_3_2;
    io_A_Valid_5_delay_5 <= io_A_Valid_5_delay_4_1;
    io_B_Valid_5_delay_1_4 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_3 <= io_B_Valid_5_delay_1_4;
    io_B_Valid_5_delay_3_2 <= io_B_Valid_5_delay_2_3;
    io_B_Valid_5_delay_4_1 <= io_B_Valid_5_delay_3_2;
    io_B_Valid_5_delay_5 <= io_B_Valid_5_delay_4_1;
    io_A_Valid_5_delay_1_5 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_4 <= io_A_Valid_5_delay_1_5;
    io_A_Valid_5_delay_3_3 <= io_A_Valid_5_delay_2_4;
    io_A_Valid_5_delay_4_2 <= io_A_Valid_5_delay_3_3;
    io_A_Valid_5_delay_5_1 <= io_A_Valid_5_delay_4_2;
    io_A_Valid_5_delay_6 <= io_A_Valid_5_delay_5_1;
    io_B_Valid_6_delay_1_4 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_3 <= io_B_Valid_6_delay_1_4;
    io_B_Valid_6_delay_3_2 <= io_B_Valid_6_delay_2_3;
    io_B_Valid_6_delay_4_1 <= io_B_Valid_6_delay_3_2;
    io_B_Valid_6_delay_5 <= io_B_Valid_6_delay_4_1;
    io_A_Valid_5_delay_1_6 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_5 <= io_A_Valid_5_delay_1_6;
    io_A_Valid_5_delay_3_4 <= io_A_Valid_5_delay_2_5;
    io_A_Valid_5_delay_4_3 <= io_A_Valid_5_delay_3_4;
    io_A_Valid_5_delay_5_2 <= io_A_Valid_5_delay_4_3;
    io_A_Valid_5_delay_6_1 <= io_A_Valid_5_delay_5_2;
    io_A_Valid_5_delay_7 <= io_A_Valid_5_delay_6_1;
    io_B_Valid_7_delay_1_4 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_3 <= io_B_Valid_7_delay_1_4;
    io_B_Valid_7_delay_3_2 <= io_B_Valid_7_delay_2_3;
    io_B_Valid_7_delay_4_1 <= io_B_Valid_7_delay_3_2;
    io_B_Valid_7_delay_5 <= io_B_Valid_7_delay_4_1;
    io_A_Valid_5_delay_1_7 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_6 <= io_A_Valid_5_delay_1_7;
    io_A_Valid_5_delay_3_5 <= io_A_Valid_5_delay_2_6;
    io_A_Valid_5_delay_4_4 <= io_A_Valid_5_delay_3_5;
    io_A_Valid_5_delay_5_3 <= io_A_Valid_5_delay_4_4;
    io_A_Valid_5_delay_6_2 <= io_A_Valid_5_delay_5_3;
    io_A_Valid_5_delay_7_1 <= io_A_Valid_5_delay_6_2;
    io_A_Valid_5_delay_8 <= io_A_Valid_5_delay_7_1;
    io_B_Valid_8_delay_1_4 <= io_B_Valid_8;
    io_B_Valid_8_delay_2_3 <= io_B_Valid_8_delay_1_4;
    io_B_Valid_8_delay_3_2 <= io_B_Valid_8_delay_2_3;
    io_B_Valid_8_delay_4_1 <= io_B_Valid_8_delay_3_2;
    io_B_Valid_8_delay_5 <= io_B_Valid_8_delay_4_1;
    io_A_Valid_5_delay_1_8 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_7 <= io_A_Valid_5_delay_1_8;
    io_A_Valid_5_delay_3_6 <= io_A_Valid_5_delay_2_7;
    io_A_Valid_5_delay_4_5 <= io_A_Valid_5_delay_3_6;
    io_A_Valid_5_delay_5_4 <= io_A_Valid_5_delay_4_5;
    io_A_Valid_5_delay_6_3 <= io_A_Valid_5_delay_5_4;
    io_A_Valid_5_delay_7_2 <= io_A_Valid_5_delay_6_3;
    io_A_Valid_5_delay_8_1 <= io_A_Valid_5_delay_7_2;
    io_A_Valid_5_delay_9 <= io_A_Valid_5_delay_8_1;
    io_B_Valid_9_delay_1_4 <= io_B_Valid_9;
    io_B_Valid_9_delay_2_3 <= io_B_Valid_9_delay_1_4;
    io_B_Valid_9_delay_3_2 <= io_B_Valid_9_delay_2_3;
    io_B_Valid_9_delay_4_1 <= io_B_Valid_9_delay_3_2;
    io_B_Valid_9_delay_5 <= io_B_Valid_9_delay_4_1;
    io_A_Valid_5_delay_1_9 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_8 <= io_A_Valid_5_delay_1_9;
    io_A_Valid_5_delay_3_7 <= io_A_Valid_5_delay_2_8;
    io_A_Valid_5_delay_4_6 <= io_A_Valid_5_delay_3_7;
    io_A_Valid_5_delay_5_5 <= io_A_Valid_5_delay_4_6;
    io_A_Valid_5_delay_6_4 <= io_A_Valid_5_delay_5_5;
    io_A_Valid_5_delay_7_3 <= io_A_Valid_5_delay_6_4;
    io_A_Valid_5_delay_8_2 <= io_A_Valid_5_delay_7_3;
    io_A_Valid_5_delay_9_1 <= io_A_Valid_5_delay_8_2;
    io_A_Valid_5_delay_10 <= io_A_Valid_5_delay_9_1;
    io_B_Valid_10_delay_1_4 <= io_B_Valid_10;
    io_B_Valid_10_delay_2_3 <= io_B_Valid_10_delay_1_4;
    io_B_Valid_10_delay_3_2 <= io_B_Valid_10_delay_2_3;
    io_B_Valid_10_delay_4_1 <= io_B_Valid_10_delay_3_2;
    io_B_Valid_10_delay_5 <= io_B_Valid_10_delay_4_1;
    io_A_Valid_5_delay_1_10 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_9 <= io_A_Valid_5_delay_1_10;
    io_A_Valid_5_delay_3_8 <= io_A_Valid_5_delay_2_9;
    io_A_Valid_5_delay_4_7 <= io_A_Valid_5_delay_3_8;
    io_A_Valid_5_delay_5_6 <= io_A_Valid_5_delay_4_7;
    io_A_Valid_5_delay_6_5 <= io_A_Valid_5_delay_5_6;
    io_A_Valid_5_delay_7_4 <= io_A_Valid_5_delay_6_5;
    io_A_Valid_5_delay_8_3 <= io_A_Valid_5_delay_7_4;
    io_A_Valid_5_delay_9_2 <= io_A_Valid_5_delay_8_3;
    io_A_Valid_5_delay_10_1 <= io_A_Valid_5_delay_9_2;
    io_A_Valid_5_delay_11 <= io_A_Valid_5_delay_10_1;
    io_B_Valid_11_delay_1_4 <= io_B_Valid_11;
    io_B_Valid_11_delay_2_3 <= io_B_Valid_11_delay_1_4;
    io_B_Valid_11_delay_3_2 <= io_B_Valid_11_delay_2_3;
    io_B_Valid_11_delay_4_1 <= io_B_Valid_11_delay_3_2;
    io_B_Valid_11_delay_5 <= io_B_Valid_11_delay_4_1;
    io_A_Valid_5_delay_1_11 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_10 <= io_A_Valid_5_delay_1_11;
    io_A_Valid_5_delay_3_9 <= io_A_Valid_5_delay_2_10;
    io_A_Valid_5_delay_4_8 <= io_A_Valid_5_delay_3_9;
    io_A_Valid_5_delay_5_7 <= io_A_Valid_5_delay_4_8;
    io_A_Valid_5_delay_6_6 <= io_A_Valid_5_delay_5_7;
    io_A_Valid_5_delay_7_5 <= io_A_Valid_5_delay_6_6;
    io_A_Valid_5_delay_8_4 <= io_A_Valid_5_delay_7_5;
    io_A_Valid_5_delay_9_3 <= io_A_Valid_5_delay_8_4;
    io_A_Valid_5_delay_10_2 <= io_A_Valid_5_delay_9_3;
    io_A_Valid_5_delay_11_1 <= io_A_Valid_5_delay_10_2;
    io_A_Valid_5_delay_12 <= io_A_Valid_5_delay_11_1;
    io_B_Valid_12_delay_1_4 <= io_B_Valid_12;
    io_B_Valid_12_delay_2_3 <= io_B_Valid_12_delay_1_4;
    io_B_Valid_12_delay_3_2 <= io_B_Valid_12_delay_2_3;
    io_B_Valid_12_delay_4_1 <= io_B_Valid_12_delay_3_2;
    io_B_Valid_12_delay_5 <= io_B_Valid_12_delay_4_1;
    io_A_Valid_5_delay_1_12 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_11 <= io_A_Valid_5_delay_1_12;
    io_A_Valid_5_delay_3_10 <= io_A_Valid_5_delay_2_11;
    io_A_Valid_5_delay_4_9 <= io_A_Valid_5_delay_3_10;
    io_A_Valid_5_delay_5_8 <= io_A_Valid_5_delay_4_9;
    io_A_Valid_5_delay_6_7 <= io_A_Valid_5_delay_5_8;
    io_A_Valid_5_delay_7_6 <= io_A_Valid_5_delay_6_7;
    io_A_Valid_5_delay_8_5 <= io_A_Valid_5_delay_7_6;
    io_A_Valid_5_delay_9_4 <= io_A_Valid_5_delay_8_5;
    io_A_Valid_5_delay_10_3 <= io_A_Valid_5_delay_9_4;
    io_A_Valid_5_delay_11_2 <= io_A_Valid_5_delay_10_3;
    io_A_Valid_5_delay_12_1 <= io_A_Valid_5_delay_11_2;
    io_A_Valid_5_delay_13 <= io_A_Valid_5_delay_12_1;
    io_B_Valid_13_delay_1_4 <= io_B_Valid_13;
    io_B_Valid_13_delay_2_3 <= io_B_Valid_13_delay_1_4;
    io_B_Valid_13_delay_3_2 <= io_B_Valid_13_delay_2_3;
    io_B_Valid_13_delay_4_1 <= io_B_Valid_13_delay_3_2;
    io_B_Valid_13_delay_5 <= io_B_Valid_13_delay_4_1;
    io_A_Valid_5_delay_1_13 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_12 <= io_A_Valid_5_delay_1_13;
    io_A_Valid_5_delay_3_11 <= io_A_Valid_5_delay_2_12;
    io_A_Valid_5_delay_4_10 <= io_A_Valid_5_delay_3_11;
    io_A_Valid_5_delay_5_9 <= io_A_Valid_5_delay_4_10;
    io_A_Valid_5_delay_6_8 <= io_A_Valid_5_delay_5_9;
    io_A_Valid_5_delay_7_7 <= io_A_Valid_5_delay_6_8;
    io_A_Valid_5_delay_8_6 <= io_A_Valid_5_delay_7_7;
    io_A_Valid_5_delay_9_5 <= io_A_Valid_5_delay_8_6;
    io_A_Valid_5_delay_10_4 <= io_A_Valid_5_delay_9_5;
    io_A_Valid_5_delay_11_3 <= io_A_Valid_5_delay_10_4;
    io_A_Valid_5_delay_12_2 <= io_A_Valid_5_delay_11_3;
    io_A_Valid_5_delay_13_1 <= io_A_Valid_5_delay_12_2;
    io_A_Valid_5_delay_14 <= io_A_Valid_5_delay_13_1;
    io_B_Valid_14_delay_1_4 <= io_B_Valid_14;
    io_B_Valid_14_delay_2_3 <= io_B_Valid_14_delay_1_4;
    io_B_Valid_14_delay_3_2 <= io_B_Valid_14_delay_2_3;
    io_B_Valid_14_delay_4_1 <= io_B_Valid_14_delay_3_2;
    io_B_Valid_14_delay_5 <= io_B_Valid_14_delay_4_1;
    io_A_Valid_5_delay_1_14 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_13 <= io_A_Valid_5_delay_1_14;
    io_A_Valid_5_delay_3_12 <= io_A_Valid_5_delay_2_13;
    io_A_Valid_5_delay_4_11 <= io_A_Valid_5_delay_3_12;
    io_A_Valid_5_delay_5_10 <= io_A_Valid_5_delay_4_11;
    io_A_Valid_5_delay_6_9 <= io_A_Valid_5_delay_5_10;
    io_A_Valid_5_delay_7_8 <= io_A_Valid_5_delay_6_9;
    io_A_Valid_5_delay_8_7 <= io_A_Valid_5_delay_7_8;
    io_A_Valid_5_delay_9_6 <= io_A_Valid_5_delay_8_7;
    io_A_Valid_5_delay_10_5 <= io_A_Valid_5_delay_9_6;
    io_A_Valid_5_delay_11_4 <= io_A_Valid_5_delay_10_5;
    io_A_Valid_5_delay_12_3 <= io_A_Valid_5_delay_11_4;
    io_A_Valid_5_delay_13_2 <= io_A_Valid_5_delay_12_3;
    io_A_Valid_5_delay_14_1 <= io_A_Valid_5_delay_13_2;
    io_A_Valid_5_delay_15 <= io_A_Valid_5_delay_14_1;
    io_B_Valid_15_delay_1_4 <= io_B_Valid_15;
    io_B_Valid_15_delay_2_3 <= io_B_Valid_15_delay_1_4;
    io_B_Valid_15_delay_3_2 <= io_B_Valid_15_delay_2_3;
    io_B_Valid_15_delay_4_1 <= io_B_Valid_15_delay_3_2;
    io_B_Valid_15_delay_5 <= io_B_Valid_15_delay_4_1;
    io_A_Valid_5_delay_1_15 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_14 <= io_A_Valid_5_delay_1_15;
    io_A_Valid_5_delay_3_13 <= io_A_Valid_5_delay_2_14;
    io_A_Valid_5_delay_4_12 <= io_A_Valid_5_delay_3_13;
    io_A_Valid_5_delay_5_11 <= io_A_Valid_5_delay_4_12;
    io_A_Valid_5_delay_6_10 <= io_A_Valid_5_delay_5_11;
    io_A_Valid_5_delay_7_9 <= io_A_Valid_5_delay_6_10;
    io_A_Valid_5_delay_8_8 <= io_A_Valid_5_delay_7_9;
    io_A_Valid_5_delay_9_7 <= io_A_Valid_5_delay_8_8;
    io_A_Valid_5_delay_10_6 <= io_A_Valid_5_delay_9_7;
    io_A_Valid_5_delay_11_5 <= io_A_Valid_5_delay_10_6;
    io_A_Valid_5_delay_12_4 <= io_A_Valid_5_delay_11_5;
    io_A_Valid_5_delay_13_3 <= io_A_Valid_5_delay_12_4;
    io_A_Valid_5_delay_14_2 <= io_A_Valid_5_delay_13_3;
    io_A_Valid_5_delay_15_1 <= io_A_Valid_5_delay_14_2;
    io_A_Valid_5_delay_16 <= io_A_Valid_5_delay_15_1;
    io_B_Valid_16_delay_1_4 <= io_B_Valid_16;
    io_B_Valid_16_delay_2_3 <= io_B_Valid_16_delay_1_4;
    io_B_Valid_16_delay_3_2 <= io_B_Valid_16_delay_2_3;
    io_B_Valid_16_delay_4_1 <= io_B_Valid_16_delay_3_2;
    io_B_Valid_16_delay_5 <= io_B_Valid_16_delay_4_1;
    io_A_Valid_5_delay_1_16 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_15 <= io_A_Valid_5_delay_1_16;
    io_A_Valid_5_delay_3_14 <= io_A_Valid_5_delay_2_15;
    io_A_Valid_5_delay_4_13 <= io_A_Valid_5_delay_3_14;
    io_A_Valid_5_delay_5_12 <= io_A_Valid_5_delay_4_13;
    io_A_Valid_5_delay_6_11 <= io_A_Valid_5_delay_5_12;
    io_A_Valid_5_delay_7_10 <= io_A_Valid_5_delay_6_11;
    io_A_Valid_5_delay_8_9 <= io_A_Valid_5_delay_7_10;
    io_A_Valid_5_delay_9_8 <= io_A_Valid_5_delay_8_9;
    io_A_Valid_5_delay_10_7 <= io_A_Valid_5_delay_9_8;
    io_A_Valid_5_delay_11_6 <= io_A_Valid_5_delay_10_7;
    io_A_Valid_5_delay_12_5 <= io_A_Valid_5_delay_11_6;
    io_A_Valid_5_delay_13_4 <= io_A_Valid_5_delay_12_5;
    io_A_Valid_5_delay_14_3 <= io_A_Valid_5_delay_13_4;
    io_A_Valid_5_delay_15_2 <= io_A_Valid_5_delay_14_3;
    io_A_Valid_5_delay_16_1 <= io_A_Valid_5_delay_15_2;
    io_A_Valid_5_delay_17 <= io_A_Valid_5_delay_16_1;
    io_B_Valid_17_delay_1_4 <= io_B_Valid_17;
    io_B_Valid_17_delay_2_3 <= io_B_Valid_17_delay_1_4;
    io_B_Valid_17_delay_3_2 <= io_B_Valid_17_delay_2_3;
    io_B_Valid_17_delay_4_1 <= io_B_Valid_17_delay_3_2;
    io_B_Valid_17_delay_5 <= io_B_Valid_17_delay_4_1;
    io_A_Valid_5_delay_1_17 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_16 <= io_A_Valid_5_delay_1_17;
    io_A_Valid_5_delay_3_15 <= io_A_Valid_5_delay_2_16;
    io_A_Valid_5_delay_4_14 <= io_A_Valid_5_delay_3_15;
    io_A_Valid_5_delay_5_13 <= io_A_Valid_5_delay_4_14;
    io_A_Valid_5_delay_6_12 <= io_A_Valid_5_delay_5_13;
    io_A_Valid_5_delay_7_11 <= io_A_Valid_5_delay_6_12;
    io_A_Valid_5_delay_8_10 <= io_A_Valid_5_delay_7_11;
    io_A_Valid_5_delay_9_9 <= io_A_Valid_5_delay_8_10;
    io_A_Valid_5_delay_10_8 <= io_A_Valid_5_delay_9_9;
    io_A_Valid_5_delay_11_7 <= io_A_Valid_5_delay_10_8;
    io_A_Valid_5_delay_12_6 <= io_A_Valid_5_delay_11_7;
    io_A_Valid_5_delay_13_5 <= io_A_Valid_5_delay_12_6;
    io_A_Valid_5_delay_14_4 <= io_A_Valid_5_delay_13_5;
    io_A_Valid_5_delay_15_3 <= io_A_Valid_5_delay_14_4;
    io_A_Valid_5_delay_16_2 <= io_A_Valid_5_delay_15_3;
    io_A_Valid_5_delay_17_1 <= io_A_Valid_5_delay_16_2;
    io_A_Valid_5_delay_18 <= io_A_Valid_5_delay_17_1;
    io_B_Valid_18_delay_1_4 <= io_B_Valid_18;
    io_B_Valid_18_delay_2_3 <= io_B_Valid_18_delay_1_4;
    io_B_Valid_18_delay_3_2 <= io_B_Valid_18_delay_2_3;
    io_B_Valid_18_delay_4_1 <= io_B_Valid_18_delay_3_2;
    io_B_Valid_18_delay_5 <= io_B_Valid_18_delay_4_1;
    io_A_Valid_5_delay_1_18 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_17 <= io_A_Valid_5_delay_1_18;
    io_A_Valid_5_delay_3_16 <= io_A_Valid_5_delay_2_17;
    io_A_Valid_5_delay_4_15 <= io_A_Valid_5_delay_3_16;
    io_A_Valid_5_delay_5_14 <= io_A_Valid_5_delay_4_15;
    io_A_Valid_5_delay_6_13 <= io_A_Valid_5_delay_5_14;
    io_A_Valid_5_delay_7_12 <= io_A_Valid_5_delay_6_13;
    io_A_Valid_5_delay_8_11 <= io_A_Valid_5_delay_7_12;
    io_A_Valid_5_delay_9_10 <= io_A_Valid_5_delay_8_11;
    io_A_Valid_5_delay_10_9 <= io_A_Valid_5_delay_9_10;
    io_A_Valid_5_delay_11_8 <= io_A_Valid_5_delay_10_9;
    io_A_Valid_5_delay_12_7 <= io_A_Valid_5_delay_11_8;
    io_A_Valid_5_delay_13_6 <= io_A_Valid_5_delay_12_7;
    io_A_Valid_5_delay_14_5 <= io_A_Valid_5_delay_13_6;
    io_A_Valid_5_delay_15_4 <= io_A_Valid_5_delay_14_5;
    io_A_Valid_5_delay_16_3 <= io_A_Valid_5_delay_15_4;
    io_A_Valid_5_delay_17_2 <= io_A_Valid_5_delay_16_3;
    io_A_Valid_5_delay_18_1 <= io_A_Valid_5_delay_17_2;
    io_A_Valid_5_delay_19 <= io_A_Valid_5_delay_18_1;
    io_B_Valid_19_delay_1_4 <= io_B_Valid_19;
    io_B_Valid_19_delay_2_3 <= io_B_Valid_19_delay_1_4;
    io_B_Valid_19_delay_3_2 <= io_B_Valid_19_delay_2_3;
    io_B_Valid_19_delay_4_1 <= io_B_Valid_19_delay_3_2;
    io_B_Valid_19_delay_5 <= io_B_Valid_19_delay_4_1;
    io_A_Valid_5_delay_1_19 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_18 <= io_A_Valid_5_delay_1_19;
    io_A_Valid_5_delay_3_17 <= io_A_Valid_5_delay_2_18;
    io_A_Valid_5_delay_4_16 <= io_A_Valid_5_delay_3_17;
    io_A_Valid_5_delay_5_15 <= io_A_Valid_5_delay_4_16;
    io_A_Valid_5_delay_6_14 <= io_A_Valid_5_delay_5_15;
    io_A_Valid_5_delay_7_13 <= io_A_Valid_5_delay_6_14;
    io_A_Valid_5_delay_8_12 <= io_A_Valid_5_delay_7_13;
    io_A_Valid_5_delay_9_11 <= io_A_Valid_5_delay_8_12;
    io_A_Valid_5_delay_10_10 <= io_A_Valid_5_delay_9_11;
    io_A_Valid_5_delay_11_9 <= io_A_Valid_5_delay_10_10;
    io_A_Valid_5_delay_12_8 <= io_A_Valid_5_delay_11_9;
    io_A_Valid_5_delay_13_7 <= io_A_Valid_5_delay_12_8;
    io_A_Valid_5_delay_14_6 <= io_A_Valid_5_delay_13_7;
    io_A_Valid_5_delay_15_5 <= io_A_Valid_5_delay_14_6;
    io_A_Valid_5_delay_16_4 <= io_A_Valid_5_delay_15_5;
    io_A_Valid_5_delay_17_3 <= io_A_Valid_5_delay_16_4;
    io_A_Valid_5_delay_18_2 <= io_A_Valid_5_delay_17_3;
    io_A_Valid_5_delay_19_1 <= io_A_Valid_5_delay_18_2;
    io_A_Valid_5_delay_20 <= io_A_Valid_5_delay_19_1;
    io_B_Valid_20_delay_1_4 <= io_B_Valid_20;
    io_B_Valid_20_delay_2_3 <= io_B_Valid_20_delay_1_4;
    io_B_Valid_20_delay_3_2 <= io_B_Valid_20_delay_2_3;
    io_B_Valid_20_delay_4_1 <= io_B_Valid_20_delay_3_2;
    io_B_Valid_20_delay_5 <= io_B_Valid_20_delay_4_1;
    io_A_Valid_5_delay_1_20 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_19 <= io_A_Valid_5_delay_1_20;
    io_A_Valid_5_delay_3_18 <= io_A_Valid_5_delay_2_19;
    io_A_Valid_5_delay_4_17 <= io_A_Valid_5_delay_3_18;
    io_A_Valid_5_delay_5_16 <= io_A_Valid_5_delay_4_17;
    io_A_Valid_5_delay_6_15 <= io_A_Valid_5_delay_5_16;
    io_A_Valid_5_delay_7_14 <= io_A_Valid_5_delay_6_15;
    io_A_Valid_5_delay_8_13 <= io_A_Valid_5_delay_7_14;
    io_A_Valid_5_delay_9_12 <= io_A_Valid_5_delay_8_13;
    io_A_Valid_5_delay_10_11 <= io_A_Valid_5_delay_9_12;
    io_A_Valid_5_delay_11_10 <= io_A_Valid_5_delay_10_11;
    io_A_Valid_5_delay_12_9 <= io_A_Valid_5_delay_11_10;
    io_A_Valid_5_delay_13_8 <= io_A_Valid_5_delay_12_9;
    io_A_Valid_5_delay_14_7 <= io_A_Valid_5_delay_13_8;
    io_A_Valid_5_delay_15_6 <= io_A_Valid_5_delay_14_7;
    io_A_Valid_5_delay_16_5 <= io_A_Valid_5_delay_15_6;
    io_A_Valid_5_delay_17_4 <= io_A_Valid_5_delay_16_5;
    io_A_Valid_5_delay_18_3 <= io_A_Valid_5_delay_17_4;
    io_A_Valid_5_delay_19_2 <= io_A_Valid_5_delay_18_3;
    io_A_Valid_5_delay_20_1 <= io_A_Valid_5_delay_19_2;
    io_A_Valid_5_delay_21 <= io_A_Valid_5_delay_20_1;
    io_B_Valid_21_delay_1_4 <= io_B_Valid_21;
    io_B_Valid_21_delay_2_3 <= io_B_Valid_21_delay_1_4;
    io_B_Valid_21_delay_3_2 <= io_B_Valid_21_delay_2_3;
    io_B_Valid_21_delay_4_1 <= io_B_Valid_21_delay_3_2;
    io_B_Valid_21_delay_5 <= io_B_Valid_21_delay_4_1;
    io_A_Valid_5_delay_1_21 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_20 <= io_A_Valid_5_delay_1_21;
    io_A_Valid_5_delay_3_19 <= io_A_Valid_5_delay_2_20;
    io_A_Valid_5_delay_4_18 <= io_A_Valid_5_delay_3_19;
    io_A_Valid_5_delay_5_17 <= io_A_Valid_5_delay_4_18;
    io_A_Valid_5_delay_6_16 <= io_A_Valid_5_delay_5_17;
    io_A_Valid_5_delay_7_15 <= io_A_Valid_5_delay_6_16;
    io_A_Valid_5_delay_8_14 <= io_A_Valid_5_delay_7_15;
    io_A_Valid_5_delay_9_13 <= io_A_Valid_5_delay_8_14;
    io_A_Valid_5_delay_10_12 <= io_A_Valid_5_delay_9_13;
    io_A_Valid_5_delay_11_11 <= io_A_Valid_5_delay_10_12;
    io_A_Valid_5_delay_12_10 <= io_A_Valid_5_delay_11_11;
    io_A_Valid_5_delay_13_9 <= io_A_Valid_5_delay_12_10;
    io_A_Valid_5_delay_14_8 <= io_A_Valid_5_delay_13_9;
    io_A_Valid_5_delay_15_7 <= io_A_Valid_5_delay_14_8;
    io_A_Valid_5_delay_16_6 <= io_A_Valid_5_delay_15_7;
    io_A_Valid_5_delay_17_5 <= io_A_Valid_5_delay_16_6;
    io_A_Valid_5_delay_18_4 <= io_A_Valid_5_delay_17_5;
    io_A_Valid_5_delay_19_3 <= io_A_Valid_5_delay_18_4;
    io_A_Valid_5_delay_20_2 <= io_A_Valid_5_delay_19_3;
    io_A_Valid_5_delay_21_1 <= io_A_Valid_5_delay_20_2;
    io_A_Valid_5_delay_22 <= io_A_Valid_5_delay_21_1;
    io_B_Valid_22_delay_1_4 <= io_B_Valid_22;
    io_B_Valid_22_delay_2_3 <= io_B_Valid_22_delay_1_4;
    io_B_Valid_22_delay_3_2 <= io_B_Valid_22_delay_2_3;
    io_B_Valid_22_delay_4_1 <= io_B_Valid_22_delay_3_2;
    io_B_Valid_22_delay_5 <= io_B_Valid_22_delay_4_1;
    io_A_Valid_5_delay_1_22 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_21 <= io_A_Valid_5_delay_1_22;
    io_A_Valid_5_delay_3_20 <= io_A_Valid_5_delay_2_21;
    io_A_Valid_5_delay_4_19 <= io_A_Valid_5_delay_3_20;
    io_A_Valid_5_delay_5_18 <= io_A_Valid_5_delay_4_19;
    io_A_Valid_5_delay_6_17 <= io_A_Valid_5_delay_5_18;
    io_A_Valid_5_delay_7_16 <= io_A_Valid_5_delay_6_17;
    io_A_Valid_5_delay_8_15 <= io_A_Valid_5_delay_7_16;
    io_A_Valid_5_delay_9_14 <= io_A_Valid_5_delay_8_15;
    io_A_Valid_5_delay_10_13 <= io_A_Valid_5_delay_9_14;
    io_A_Valid_5_delay_11_12 <= io_A_Valid_5_delay_10_13;
    io_A_Valid_5_delay_12_11 <= io_A_Valid_5_delay_11_12;
    io_A_Valid_5_delay_13_10 <= io_A_Valid_5_delay_12_11;
    io_A_Valid_5_delay_14_9 <= io_A_Valid_5_delay_13_10;
    io_A_Valid_5_delay_15_8 <= io_A_Valid_5_delay_14_9;
    io_A_Valid_5_delay_16_7 <= io_A_Valid_5_delay_15_8;
    io_A_Valid_5_delay_17_6 <= io_A_Valid_5_delay_16_7;
    io_A_Valid_5_delay_18_5 <= io_A_Valid_5_delay_17_6;
    io_A_Valid_5_delay_19_4 <= io_A_Valid_5_delay_18_5;
    io_A_Valid_5_delay_20_3 <= io_A_Valid_5_delay_19_4;
    io_A_Valid_5_delay_21_2 <= io_A_Valid_5_delay_20_3;
    io_A_Valid_5_delay_22_1 <= io_A_Valid_5_delay_21_2;
    io_A_Valid_5_delay_23 <= io_A_Valid_5_delay_22_1;
    io_B_Valid_23_delay_1_4 <= io_B_Valid_23;
    io_B_Valid_23_delay_2_3 <= io_B_Valid_23_delay_1_4;
    io_B_Valid_23_delay_3_2 <= io_B_Valid_23_delay_2_3;
    io_B_Valid_23_delay_4_1 <= io_B_Valid_23_delay_3_2;
    io_B_Valid_23_delay_5 <= io_B_Valid_23_delay_4_1;
    io_A_Valid_5_delay_1_23 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_22 <= io_A_Valid_5_delay_1_23;
    io_A_Valid_5_delay_3_21 <= io_A_Valid_5_delay_2_22;
    io_A_Valid_5_delay_4_20 <= io_A_Valid_5_delay_3_21;
    io_A_Valid_5_delay_5_19 <= io_A_Valid_5_delay_4_20;
    io_A_Valid_5_delay_6_18 <= io_A_Valid_5_delay_5_19;
    io_A_Valid_5_delay_7_17 <= io_A_Valid_5_delay_6_18;
    io_A_Valid_5_delay_8_16 <= io_A_Valid_5_delay_7_17;
    io_A_Valid_5_delay_9_15 <= io_A_Valid_5_delay_8_16;
    io_A_Valid_5_delay_10_14 <= io_A_Valid_5_delay_9_15;
    io_A_Valid_5_delay_11_13 <= io_A_Valid_5_delay_10_14;
    io_A_Valid_5_delay_12_12 <= io_A_Valid_5_delay_11_13;
    io_A_Valid_5_delay_13_11 <= io_A_Valid_5_delay_12_12;
    io_A_Valid_5_delay_14_10 <= io_A_Valid_5_delay_13_11;
    io_A_Valid_5_delay_15_9 <= io_A_Valid_5_delay_14_10;
    io_A_Valid_5_delay_16_8 <= io_A_Valid_5_delay_15_9;
    io_A_Valid_5_delay_17_7 <= io_A_Valid_5_delay_16_8;
    io_A_Valid_5_delay_18_6 <= io_A_Valid_5_delay_17_7;
    io_A_Valid_5_delay_19_5 <= io_A_Valid_5_delay_18_6;
    io_A_Valid_5_delay_20_4 <= io_A_Valid_5_delay_19_5;
    io_A_Valid_5_delay_21_3 <= io_A_Valid_5_delay_20_4;
    io_A_Valid_5_delay_22_2 <= io_A_Valid_5_delay_21_3;
    io_A_Valid_5_delay_23_1 <= io_A_Valid_5_delay_22_2;
    io_A_Valid_5_delay_24 <= io_A_Valid_5_delay_23_1;
    io_B_Valid_24_delay_1_4 <= io_B_Valid_24;
    io_B_Valid_24_delay_2_3 <= io_B_Valid_24_delay_1_4;
    io_B_Valid_24_delay_3_2 <= io_B_Valid_24_delay_2_3;
    io_B_Valid_24_delay_4_1 <= io_B_Valid_24_delay_3_2;
    io_B_Valid_24_delay_5 <= io_B_Valid_24_delay_4_1;
    io_A_Valid_5_delay_1_24 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_23 <= io_A_Valid_5_delay_1_24;
    io_A_Valid_5_delay_3_22 <= io_A_Valid_5_delay_2_23;
    io_A_Valid_5_delay_4_21 <= io_A_Valid_5_delay_3_22;
    io_A_Valid_5_delay_5_20 <= io_A_Valid_5_delay_4_21;
    io_A_Valid_5_delay_6_19 <= io_A_Valid_5_delay_5_20;
    io_A_Valid_5_delay_7_18 <= io_A_Valid_5_delay_6_19;
    io_A_Valid_5_delay_8_17 <= io_A_Valid_5_delay_7_18;
    io_A_Valid_5_delay_9_16 <= io_A_Valid_5_delay_8_17;
    io_A_Valid_5_delay_10_15 <= io_A_Valid_5_delay_9_16;
    io_A_Valid_5_delay_11_14 <= io_A_Valid_5_delay_10_15;
    io_A_Valid_5_delay_12_13 <= io_A_Valid_5_delay_11_14;
    io_A_Valid_5_delay_13_12 <= io_A_Valid_5_delay_12_13;
    io_A_Valid_5_delay_14_11 <= io_A_Valid_5_delay_13_12;
    io_A_Valid_5_delay_15_10 <= io_A_Valid_5_delay_14_11;
    io_A_Valid_5_delay_16_9 <= io_A_Valid_5_delay_15_10;
    io_A_Valid_5_delay_17_8 <= io_A_Valid_5_delay_16_9;
    io_A_Valid_5_delay_18_7 <= io_A_Valid_5_delay_17_8;
    io_A_Valid_5_delay_19_6 <= io_A_Valid_5_delay_18_7;
    io_A_Valid_5_delay_20_5 <= io_A_Valid_5_delay_19_6;
    io_A_Valid_5_delay_21_4 <= io_A_Valid_5_delay_20_5;
    io_A_Valid_5_delay_22_3 <= io_A_Valid_5_delay_21_4;
    io_A_Valid_5_delay_23_2 <= io_A_Valid_5_delay_22_3;
    io_A_Valid_5_delay_24_1 <= io_A_Valid_5_delay_23_2;
    io_A_Valid_5_delay_25 <= io_A_Valid_5_delay_24_1;
    io_B_Valid_25_delay_1_4 <= io_B_Valid_25;
    io_B_Valid_25_delay_2_3 <= io_B_Valid_25_delay_1_4;
    io_B_Valid_25_delay_3_2 <= io_B_Valid_25_delay_2_3;
    io_B_Valid_25_delay_4_1 <= io_B_Valid_25_delay_3_2;
    io_B_Valid_25_delay_5 <= io_B_Valid_25_delay_4_1;
    io_A_Valid_5_delay_1_25 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_24 <= io_A_Valid_5_delay_1_25;
    io_A_Valid_5_delay_3_23 <= io_A_Valid_5_delay_2_24;
    io_A_Valid_5_delay_4_22 <= io_A_Valid_5_delay_3_23;
    io_A_Valid_5_delay_5_21 <= io_A_Valid_5_delay_4_22;
    io_A_Valid_5_delay_6_20 <= io_A_Valid_5_delay_5_21;
    io_A_Valid_5_delay_7_19 <= io_A_Valid_5_delay_6_20;
    io_A_Valid_5_delay_8_18 <= io_A_Valid_5_delay_7_19;
    io_A_Valid_5_delay_9_17 <= io_A_Valid_5_delay_8_18;
    io_A_Valid_5_delay_10_16 <= io_A_Valid_5_delay_9_17;
    io_A_Valid_5_delay_11_15 <= io_A_Valid_5_delay_10_16;
    io_A_Valid_5_delay_12_14 <= io_A_Valid_5_delay_11_15;
    io_A_Valid_5_delay_13_13 <= io_A_Valid_5_delay_12_14;
    io_A_Valid_5_delay_14_12 <= io_A_Valid_5_delay_13_13;
    io_A_Valid_5_delay_15_11 <= io_A_Valid_5_delay_14_12;
    io_A_Valid_5_delay_16_10 <= io_A_Valid_5_delay_15_11;
    io_A_Valid_5_delay_17_9 <= io_A_Valid_5_delay_16_10;
    io_A_Valid_5_delay_18_8 <= io_A_Valid_5_delay_17_9;
    io_A_Valid_5_delay_19_7 <= io_A_Valid_5_delay_18_8;
    io_A_Valid_5_delay_20_6 <= io_A_Valid_5_delay_19_7;
    io_A_Valid_5_delay_21_5 <= io_A_Valid_5_delay_20_6;
    io_A_Valid_5_delay_22_4 <= io_A_Valid_5_delay_21_5;
    io_A_Valid_5_delay_23_3 <= io_A_Valid_5_delay_22_4;
    io_A_Valid_5_delay_24_2 <= io_A_Valid_5_delay_23_3;
    io_A_Valid_5_delay_25_1 <= io_A_Valid_5_delay_24_2;
    io_A_Valid_5_delay_26 <= io_A_Valid_5_delay_25_1;
    io_B_Valid_26_delay_1_4 <= io_B_Valid_26;
    io_B_Valid_26_delay_2_3 <= io_B_Valid_26_delay_1_4;
    io_B_Valid_26_delay_3_2 <= io_B_Valid_26_delay_2_3;
    io_B_Valid_26_delay_4_1 <= io_B_Valid_26_delay_3_2;
    io_B_Valid_26_delay_5 <= io_B_Valid_26_delay_4_1;
    io_A_Valid_5_delay_1_26 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_25 <= io_A_Valid_5_delay_1_26;
    io_A_Valid_5_delay_3_24 <= io_A_Valid_5_delay_2_25;
    io_A_Valid_5_delay_4_23 <= io_A_Valid_5_delay_3_24;
    io_A_Valid_5_delay_5_22 <= io_A_Valid_5_delay_4_23;
    io_A_Valid_5_delay_6_21 <= io_A_Valid_5_delay_5_22;
    io_A_Valid_5_delay_7_20 <= io_A_Valid_5_delay_6_21;
    io_A_Valid_5_delay_8_19 <= io_A_Valid_5_delay_7_20;
    io_A_Valid_5_delay_9_18 <= io_A_Valid_5_delay_8_19;
    io_A_Valid_5_delay_10_17 <= io_A_Valid_5_delay_9_18;
    io_A_Valid_5_delay_11_16 <= io_A_Valid_5_delay_10_17;
    io_A_Valid_5_delay_12_15 <= io_A_Valid_5_delay_11_16;
    io_A_Valid_5_delay_13_14 <= io_A_Valid_5_delay_12_15;
    io_A_Valid_5_delay_14_13 <= io_A_Valid_5_delay_13_14;
    io_A_Valid_5_delay_15_12 <= io_A_Valid_5_delay_14_13;
    io_A_Valid_5_delay_16_11 <= io_A_Valid_5_delay_15_12;
    io_A_Valid_5_delay_17_10 <= io_A_Valid_5_delay_16_11;
    io_A_Valid_5_delay_18_9 <= io_A_Valid_5_delay_17_10;
    io_A_Valid_5_delay_19_8 <= io_A_Valid_5_delay_18_9;
    io_A_Valid_5_delay_20_7 <= io_A_Valid_5_delay_19_8;
    io_A_Valid_5_delay_21_6 <= io_A_Valid_5_delay_20_7;
    io_A_Valid_5_delay_22_5 <= io_A_Valid_5_delay_21_6;
    io_A_Valid_5_delay_23_4 <= io_A_Valid_5_delay_22_5;
    io_A_Valid_5_delay_24_3 <= io_A_Valid_5_delay_23_4;
    io_A_Valid_5_delay_25_2 <= io_A_Valid_5_delay_24_3;
    io_A_Valid_5_delay_26_1 <= io_A_Valid_5_delay_25_2;
    io_A_Valid_5_delay_27 <= io_A_Valid_5_delay_26_1;
    io_B_Valid_27_delay_1_4 <= io_B_Valid_27;
    io_B_Valid_27_delay_2_3 <= io_B_Valid_27_delay_1_4;
    io_B_Valid_27_delay_3_2 <= io_B_Valid_27_delay_2_3;
    io_B_Valid_27_delay_4_1 <= io_B_Valid_27_delay_3_2;
    io_B_Valid_27_delay_5 <= io_B_Valid_27_delay_4_1;
    io_A_Valid_5_delay_1_27 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_26 <= io_A_Valid_5_delay_1_27;
    io_A_Valid_5_delay_3_25 <= io_A_Valid_5_delay_2_26;
    io_A_Valid_5_delay_4_24 <= io_A_Valid_5_delay_3_25;
    io_A_Valid_5_delay_5_23 <= io_A_Valid_5_delay_4_24;
    io_A_Valid_5_delay_6_22 <= io_A_Valid_5_delay_5_23;
    io_A_Valid_5_delay_7_21 <= io_A_Valid_5_delay_6_22;
    io_A_Valid_5_delay_8_20 <= io_A_Valid_5_delay_7_21;
    io_A_Valid_5_delay_9_19 <= io_A_Valid_5_delay_8_20;
    io_A_Valid_5_delay_10_18 <= io_A_Valid_5_delay_9_19;
    io_A_Valid_5_delay_11_17 <= io_A_Valid_5_delay_10_18;
    io_A_Valid_5_delay_12_16 <= io_A_Valid_5_delay_11_17;
    io_A_Valid_5_delay_13_15 <= io_A_Valid_5_delay_12_16;
    io_A_Valid_5_delay_14_14 <= io_A_Valid_5_delay_13_15;
    io_A_Valid_5_delay_15_13 <= io_A_Valid_5_delay_14_14;
    io_A_Valid_5_delay_16_12 <= io_A_Valid_5_delay_15_13;
    io_A_Valid_5_delay_17_11 <= io_A_Valid_5_delay_16_12;
    io_A_Valid_5_delay_18_10 <= io_A_Valid_5_delay_17_11;
    io_A_Valid_5_delay_19_9 <= io_A_Valid_5_delay_18_10;
    io_A_Valid_5_delay_20_8 <= io_A_Valid_5_delay_19_9;
    io_A_Valid_5_delay_21_7 <= io_A_Valid_5_delay_20_8;
    io_A_Valid_5_delay_22_6 <= io_A_Valid_5_delay_21_7;
    io_A_Valid_5_delay_23_5 <= io_A_Valid_5_delay_22_6;
    io_A_Valid_5_delay_24_4 <= io_A_Valid_5_delay_23_5;
    io_A_Valid_5_delay_25_3 <= io_A_Valid_5_delay_24_4;
    io_A_Valid_5_delay_26_2 <= io_A_Valid_5_delay_25_3;
    io_A_Valid_5_delay_27_1 <= io_A_Valid_5_delay_26_2;
    io_A_Valid_5_delay_28 <= io_A_Valid_5_delay_27_1;
    io_B_Valid_28_delay_1_4 <= io_B_Valid_28;
    io_B_Valid_28_delay_2_3 <= io_B_Valid_28_delay_1_4;
    io_B_Valid_28_delay_3_2 <= io_B_Valid_28_delay_2_3;
    io_B_Valid_28_delay_4_1 <= io_B_Valid_28_delay_3_2;
    io_B_Valid_28_delay_5 <= io_B_Valid_28_delay_4_1;
    io_A_Valid_5_delay_1_28 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_27 <= io_A_Valid_5_delay_1_28;
    io_A_Valid_5_delay_3_26 <= io_A_Valid_5_delay_2_27;
    io_A_Valid_5_delay_4_25 <= io_A_Valid_5_delay_3_26;
    io_A_Valid_5_delay_5_24 <= io_A_Valid_5_delay_4_25;
    io_A_Valid_5_delay_6_23 <= io_A_Valid_5_delay_5_24;
    io_A_Valid_5_delay_7_22 <= io_A_Valid_5_delay_6_23;
    io_A_Valid_5_delay_8_21 <= io_A_Valid_5_delay_7_22;
    io_A_Valid_5_delay_9_20 <= io_A_Valid_5_delay_8_21;
    io_A_Valid_5_delay_10_19 <= io_A_Valid_5_delay_9_20;
    io_A_Valid_5_delay_11_18 <= io_A_Valid_5_delay_10_19;
    io_A_Valid_5_delay_12_17 <= io_A_Valid_5_delay_11_18;
    io_A_Valid_5_delay_13_16 <= io_A_Valid_5_delay_12_17;
    io_A_Valid_5_delay_14_15 <= io_A_Valid_5_delay_13_16;
    io_A_Valid_5_delay_15_14 <= io_A_Valid_5_delay_14_15;
    io_A_Valid_5_delay_16_13 <= io_A_Valid_5_delay_15_14;
    io_A_Valid_5_delay_17_12 <= io_A_Valid_5_delay_16_13;
    io_A_Valid_5_delay_18_11 <= io_A_Valid_5_delay_17_12;
    io_A_Valid_5_delay_19_10 <= io_A_Valid_5_delay_18_11;
    io_A_Valid_5_delay_20_9 <= io_A_Valid_5_delay_19_10;
    io_A_Valid_5_delay_21_8 <= io_A_Valid_5_delay_20_9;
    io_A_Valid_5_delay_22_7 <= io_A_Valid_5_delay_21_8;
    io_A_Valid_5_delay_23_6 <= io_A_Valid_5_delay_22_7;
    io_A_Valid_5_delay_24_5 <= io_A_Valid_5_delay_23_6;
    io_A_Valid_5_delay_25_4 <= io_A_Valid_5_delay_24_5;
    io_A_Valid_5_delay_26_3 <= io_A_Valid_5_delay_25_4;
    io_A_Valid_5_delay_27_2 <= io_A_Valid_5_delay_26_3;
    io_A_Valid_5_delay_28_1 <= io_A_Valid_5_delay_27_2;
    io_A_Valid_5_delay_29 <= io_A_Valid_5_delay_28_1;
    io_B_Valid_29_delay_1_4 <= io_B_Valid_29;
    io_B_Valid_29_delay_2_3 <= io_B_Valid_29_delay_1_4;
    io_B_Valid_29_delay_3_2 <= io_B_Valid_29_delay_2_3;
    io_B_Valid_29_delay_4_1 <= io_B_Valid_29_delay_3_2;
    io_B_Valid_29_delay_5 <= io_B_Valid_29_delay_4_1;
    io_A_Valid_5_delay_1_29 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_28 <= io_A_Valid_5_delay_1_29;
    io_A_Valid_5_delay_3_27 <= io_A_Valid_5_delay_2_28;
    io_A_Valid_5_delay_4_26 <= io_A_Valid_5_delay_3_27;
    io_A_Valid_5_delay_5_25 <= io_A_Valid_5_delay_4_26;
    io_A_Valid_5_delay_6_24 <= io_A_Valid_5_delay_5_25;
    io_A_Valid_5_delay_7_23 <= io_A_Valid_5_delay_6_24;
    io_A_Valid_5_delay_8_22 <= io_A_Valid_5_delay_7_23;
    io_A_Valid_5_delay_9_21 <= io_A_Valid_5_delay_8_22;
    io_A_Valid_5_delay_10_20 <= io_A_Valid_5_delay_9_21;
    io_A_Valid_5_delay_11_19 <= io_A_Valid_5_delay_10_20;
    io_A_Valid_5_delay_12_18 <= io_A_Valid_5_delay_11_19;
    io_A_Valid_5_delay_13_17 <= io_A_Valid_5_delay_12_18;
    io_A_Valid_5_delay_14_16 <= io_A_Valid_5_delay_13_17;
    io_A_Valid_5_delay_15_15 <= io_A_Valid_5_delay_14_16;
    io_A_Valid_5_delay_16_14 <= io_A_Valid_5_delay_15_15;
    io_A_Valid_5_delay_17_13 <= io_A_Valid_5_delay_16_14;
    io_A_Valid_5_delay_18_12 <= io_A_Valid_5_delay_17_13;
    io_A_Valid_5_delay_19_11 <= io_A_Valid_5_delay_18_12;
    io_A_Valid_5_delay_20_10 <= io_A_Valid_5_delay_19_11;
    io_A_Valid_5_delay_21_9 <= io_A_Valid_5_delay_20_10;
    io_A_Valid_5_delay_22_8 <= io_A_Valid_5_delay_21_9;
    io_A_Valid_5_delay_23_7 <= io_A_Valid_5_delay_22_8;
    io_A_Valid_5_delay_24_6 <= io_A_Valid_5_delay_23_7;
    io_A_Valid_5_delay_25_5 <= io_A_Valid_5_delay_24_6;
    io_A_Valid_5_delay_26_4 <= io_A_Valid_5_delay_25_5;
    io_A_Valid_5_delay_27_3 <= io_A_Valid_5_delay_26_4;
    io_A_Valid_5_delay_28_2 <= io_A_Valid_5_delay_27_3;
    io_A_Valid_5_delay_29_1 <= io_A_Valid_5_delay_28_2;
    io_A_Valid_5_delay_30 <= io_A_Valid_5_delay_29_1;
    io_B_Valid_30_delay_1_4 <= io_B_Valid_30;
    io_B_Valid_30_delay_2_3 <= io_B_Valid_30_delay_1_4;
    io_B_Valid_30_delay_3_2 <= io_B_Valid_30_delay_2_3;
    io_B_Valid_30_delay_4_1 <= io_B_Valid_30_delay_3_2;
    io_B_Valid_30_delay_5 <= io_B_Valid_30_delay_4_1;
    io_A_Valid_5_delay_1_30 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_29 <= io_A_Valid_5_delay_1_30;
    io_A_Valid_5_delay_3_28 <= io_A_Valid_5_delay_2_29;
    io_A_Valid_5_delay_4_27 <= io_A_Valid_5_delay_3_28;
    io_A_Valid_5_delay_5_26 <= io_A_Valid_5_delay_4_27;
    io_A_Valid_5_delay_6_25 <= io_A_Valid_5_delay_5_26;
    io_A_Valid_5_delay_7_24 <= io_A_Valid_5_delay_6_25;
    io_A_Valid_5_delay_8_23 <= io_A_Valid_5_delay_7_24;
    io_A_Valid_5_delay_9_22 <= io_A_Valid_5_delay_8_23;
    io_A_Valid_5_delay_10_21 <= io_A_Valid_5_delay_9_22;
    io_A_Valid_5_delay_11_20 <= io_A_Valid_5_delay_10_21;
    io_A_Valid_5_delay_12_19 <= io_A_Valid_5_delay_11_20;
    io_A_Valid_5_delay_13_18 <= io_A_Valid_5_delay_12_19;
    io_A_Valid_5_delay_14_17 <= io_A_Valid_5_delay_13_18;
    io_A_Valid_5_delay_15_16 <= io_A_Valid_5_delay_14_17;
    io_A_Valid_5_delay_16_15 <= io_A_Valid_5_delay_15_16;
    io_A_Valid_5_delay_17_14 <= io_A_Valid_5_delay_16_15;
    io_A_Valid_5_delay_18_13 <= io_A_Valid_5_delay_17_14;
    io_A_Valid_5_delay_19_12 <= io_A_Valid_5_delay_18_13;
    io_A_Valid_5_delay_20_11 <= io_A_Valid_5_delay_19_12;
    io_A_Valid_5_delay_21_10 <= io_A_Valid_5_delay_20_11;
    io_A_Valid_5_delay_22_9 <= io_A_Valid_5_delay_21_10;
    io_A_Valid_5_delay_23_8 <= io_A_Valid_5_delay_22_9;
    io_A_Valid_5_delay_24_7 <= io_A_Valid_5_delay_23_8;
    io_A_Valid_5_delay_25_6 <= io_A_Valid_5_delay_24_7;
    io_A_Valid_5_delay_26_5 <= io_A_Valid_5_delay_25_6;
    io_A_Valid_5_delay_27_4 <= io_A_Valid_5_delay_26_5;
    io_A_Valid_5_delay_28_3 <= io_A_Valid_5_delay_27_4;
    io_A_Valid_5_delay_29_2 <= io_A_Valid_5_delay_28_3;
    io_A_Valid_5_delay_30_1 <= io_A_Valid_5_delay_29_2;
    io_A_Valid_5_delay_31 <= io_A_Valid_5_delay_30_1;
    io_B_Valid_31_delay_1_4 <= io_B_Valid_31;
    io_B_Valid_31_delay_2_3 <= io_B_Valid_31_delay_1_4;
    io_B_Valid_31_delay_3_2 <= io_B_Valid_31_delay_2_3;
    io_B_Valid_31_delay_4_1 <= io_B_Valid_31_delay_3_2;
    io_B_Valid_31_delay_5 <= io_B_Valid_31_delay_4_1;
    io_A_Valid_5_delay_1_31 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_30 <= io_A_Valid_5_delay_1_31;
    io_A_Valid_5_delay_3_29 <= io_A_Valid_5_delay_2_30;
    io_A_Valid_5_delay_4_28 <= io_A_Valid_5_delay_3_29;
    io_A_Valid_5_delay_5_27 <= io_A_Valid_5_delay_4_28;
    io_A_Valid_5_delay_6_26 <= io_A_Valid_5_delay_5_27;
    io_A_Valid_5_delay_7_25 <= io_A_Valid_5_delay_6_26;
    io_A_Valid_5_delay_8_24 <= io_A_Valid_5_delay_7_25;
    io_A_Valid_5_delay_9_23 <= io_A_Valid_5_delay_8_24;
    io_A_Valid_5_delay_10_22 <= io_A_Valid_5_delay_9_23;
    io_A_Valid_5_delay_11_21 <= io_A_Valid_5_delay_10_22;
    io_A_Valid_5_delay_12_20 <= io_A_Valid_5_delay_11_21;
    io_A_Valid_5_delay_13_19 <= io_A_Valid_5_delay_12_20;
    io_A_Valid_5_delay_14_18 <= io_A_Valid_5_delay_13_19;
    io_A_Valid_5_delay_15_17 <= io_A_Valid_5_delay_14_18;
    io_A_Valid_5_delay_16_16 <= io_A_Valid_5_delay_15_17;
    io_A_Valid_5_delay_17_15 <= io_A_Valid_5_delay_16_16;
    io_A_Valid_5_delay_18_14 <= io_A_Valid_5_delay_17_15;
    io_A_Valid_5_delay_19_13 <= io_A_Valid_5_delay_18_14;
    io_A_Valid_5_delay_20_12 <= io_A_Valid_5_delay_19_13;
    io_A_Valid_5_delay_21_11 <= io_A_Valid_5_delay_20_12;
    io_A_Valid_5_delay_22_10 <= io_A_Valid_5_delay_21_11;
    io_A_Valid_5_delay_23_9 <= io_A_Valid_5_delay_22_10;
    io_A_Valid_5_delay_24_8 <= io_A_Valid_5_delay_23_9;
    io_A_Valid_5_delay_25_7 <= io_A_Valid_5_delay_24_8;
    io_A_Valid_5_delay_26_6 <= io_A_Valid_5_delay_25_7;
    io_A_Valid_5_delay_27_5 <= io_A_Valid_5_delay_26_6;
    io_A_Valid_5_delay_28_4 <= io_A_Valid_5_delay_27_5;
    io_A_Valid_5_delay_29_3 <= io_A_Valid_5_delay_28_4;
    io_A_Valid_5_delay_30_2 <= io_A_Valid_5_delay_29_3;
    io_A_Valid_5_delay_31_1 <= io_A_Valid_5_delay_30_2;
    io_A_Valid_5_delay_32 <= io_A_Valid_5_delay_31_1;
    io_B_Valid_32_delay_1_4 <= io_B_Valid_32;
    io_B_Valid_32_delay_2_3 <= io_B_Valid_32_delay_1_4;
    io_B_Valid_32_delay_3_2 <= io_B_Valid_32_delay_2_3;
    io_B_Valid_32_delay_4_1 <= io_B_Valid_32_delay_3_2;
    io_B_Valid_32_delay_5 <= io_B_Valid_32_delay_4_1;
    io_A_Valid_5_delay_1_32 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_31 <= io_A_Valid_5_delay_1_32;
    io_A_Valid_5_delay_3_30 <= io_A_Valid_5_delay_2_31;
    io_A_Valid_5_delay_4_29 <= io_A_Valid_5_delay_3_30;
    io_A_Valid_5_delay_5_28 <= io_A_Valid_5_delay_4_29;
    io_A_Valid_5_delay_6_27 <= io_A_Valid_5_delay_5_28;
    io_A_Valid_5_delay_7_26 <= io_A_Valid_5_delay_6_27;
    io_A_Valid_5_delay_8_25 <= io_A_Valid_5_delay_7_26;
    io_A_Valid_5_delay_9_24 <= io_A_Valid_5_delay_8_25;
    io_A_Valid_5_delay_10_23 <= io_A_Valid_5_delay_9_24;
    io_A_Valid_5_delay_11_22 <= io_A_Valid_5_delay_10_23;
    io_A_Valid_5_delay_12_21 <= io_A_Valid_5_delay_11_22;
    io_A_Valid_5_delay_13_20 <= io_A_Valid_5_delay_12_21;
    io_A_Valid_5_delay_14_19 <= io_A_Valid_5_delay_13_20;
    io_A_Valid_5_delay_15_18 <= io_A_Valid_5_delay_14_19;
    io_A_Valid_5_delay_16_17 <= io_A_Valid_5_delay_15_18;
    io_A_Valid_5_delay_17_16 <= io_A_Valid_5_delay_16_17;
    io_A_Valid_5_delay_18_15 <= io_A_Valid_5_delay_17_16;
    io_A_Valid_5_delay_19_14 <= io_A_Valid_5_delay_18_15;
    io_A_Valid_5_delay_20_13 <= io_A_Valid_5_delay_19_14;
    io_A_Valid_5_delay_21_12 <= io_A_Valid_5_delay_20_13;
    io_A_Valid_5_delay_22_11 <= io_A_Valid_5_delay_21_12;
    io_A_Valid_5_delay_23_10 <= io_A_Valid_5_delay_22_11;
    io_A_Valid_5_delay_24_9 <= io_A_Valid_5_delay_23_10;
    io_A_Valid_5_delay_25_8 <= io_A_Valid_5_delay_24_9;
    io_A_Valid_5_delay_26_7 <= io_A_Valid_5_delay_25_8;
    io_A_Valid_5_delay_27_6 <= io_A_Valid_5_delay_26_7;
    io_A_Valid_5_delay_28_5 <= io_A_Valid_5_delay_27_6;
    io_A_Valid_5_delay_29_4 <= io_A_Valid_5_delay_28_5;
    io_A_Valid_5_delay_30_3 <= io_A_Valid_5_delay_29_4;
    io_A_Valid_5_delay_31_2 <= io_A_Valid_5_delay_30_3;
    io_A_Valid_5_delay_32_1 <= io_A_Valid_5_delay_31_2;
    io_A_Valid_5_delay_33 <= io_A_Valid_5_delay_32_1;
    io_B_Valid_33_delay_1_4 <= io_B_Valid_33;
    io_B_Valid_33_delay_2_3 <= io_B_Valid_33_delay_1_4;
    io_B_Valid_33_delay_3_2 <= io_B_Valid_33_delay_2_3;
    io_B_Valid_33_delay_4_1 <= io_B_Valid_33_delay_3_2;
    io_B_Valid_33_delay_5 <= io_B_Valid_33_delay_4_1;
    io_A_Valid_5_delay_1_33 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_32 <= io_A_Valid_5_delay_1_33;
    io_A_Valid_5_delay_3_31 <= io_A_Valid_5_delay_2_32;
    io_A_Valid_5_delay_4_30 <= io_A_Valid_5_delay_3_31;
    io_A_Valid_5_delay_5_29 <= io_A_Valid_5_delay_4_30;
    io_A_Valid_5_delay_6_28 <= io_A_Valid_5_delay_5_29;
    io_A_Valid_5_delay_7_27 <= io_A_Valid_5_delay_6_28;
    io_A_Valid_5_delay_8_26 <= io_A_Valid_5_delay_7_27;
    io_A_Valid_5_delay_9_25 <= io_A_Valid_5_delay_8_26;
    io_A_Valid_5_delay_10_24 <= io_A_Valid_5_delay_9_25;
    io_A_Valid_5_delay_11_23 <= io_A_Valid_5_delay_10_24;
    io_A_Valid_5_delay_12_22 <= io_A_Valid_5_delay_11_23;
    io_A_Valid_5_delay_13_21 <= io_A_Valid_5_delay_12_22;
    io_A_Valid_5_delay_14_20 <= io_A_Valid_5_delay_13_21;
    io_A_Valid_5_delay_15_19 <= io_A_Valid_5_delay_14_20;
    io_A_Valid_5_delay_16_18 <= io_A_Valid_5_delay_15_19;
    io_A_Valid_5_delay_17_17 <= io_A_Valid_5_delay_16_18;
    io_A_Valid_5_delay_18_16 <= io_A_Valid_5_delay_17_17;
    io_A_Valid_5_delay_19_15 <= io_A_Valid_5_delay_18_16;
    io_A_Valid_5_delay_20_14 <= io_A_Valid_5_delay_19_15;
    io_A_Valid_5_delay_21_13 <= io_A_Valid_5_delay_20_14;
    io_A_Valid_5_delay_22_12 <= io_A_Valid_5_delay_21_13;
    io_A_Valid_5_delay_23_11 <= io_A_Valid_5_delay_22_12;
    io_A_Valid_5_delay_24_10 <= io_A_Valid_5_delay_23_11;
    io_A_Valid_5_delay_25_9 <= io_A_Valid_5_delay_24_10;
    io_A_Valid_5_delay_26_8 <= io_A_Valid_5_delay_25_9;
    io_A_Valid_5_delay_27_7 <= io_A_Valid_5_delay_26_8;
    io_A_Valid_5_delay_28_6 <= io_A_Valid_5_delay_27_7;
    io_A_Valid_5_delay_29_5 <= io_A_Valid_5_delay_28_6;
    io_A_Valid_5_delay_30_4 <= io_A_Valid_5_delay_29_5;
    io_A_Valid_5_delay_31_3 <= io_A_Valid_5_delay_30_4;
    io_A_Valid_5_delay_32_2 <= io_A_Valid_5_delay_31_3;
    io_A_Valid_5_delay_33_1 <= io_A_Valid_5_delay_32_2;
    io_A_Valid_5_delay_34 <= io_A_Valid_5_delay_33_1;
    io_B_Valid_34_delay_1_4 <= io_B_Valid_34;
    io_B_Valid_34_delay_2_3 <= io_B_Valid_34_delay_1_4;
    io_B_Valid_34_delay_3_2 <= io_B_Valid_34_delay_2_3;
    io_B_Valid_34_delay_4_1 <= io_B_Valid_34_delay_3_2;
    io_B_Valid_34_delay_5 <= io_B_Valid_34_delay_4_1;
    io_A_Valid_5_delay_1_34 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_33 <= io_A_Valid_5_delay_1_34;
    io_A_Valid_5_delay_3_32 <= io_A_Valid_5_delay_2_33;
    io_A_Valid_5_delay_4_31 <= io_A_Valid_5_delay_3_32;
    io_A_Valid_5_delay_5_30 <= io_A_Valid_5_delay_4_31;
    io_A_Valid_5_delay_6_29 <= io_A_Valid_5_delay_5_30;
    io_A_Valid_5_delay_7_28 <= io_A_Valid_5_delay_6_29;
    io_A_Valid_5_delay_8_27 <= io_A_Valid_5_delay_7_28;
    io_A_Valid_5_delay_9_26 <= io_A_Valid_5_delay_8_27;
    io_A_Valid_5_delay_10_25 <= io_A_Valid_5_delay_9_26;
    io_A_Valid_5_delay_11_24 <= io_A_Valid_5_delay_10_25;
    io_A_Valid_5_delay_12_23 <= io_A_Valid_5_delay_11_24;
    io_A_Valid_5_delay_13_22 <= io_A_Valid_5_delay_12_23;
    io_A_Valid_5_delay_14_21 <= io_A_Valid_5_delay_13_22;
    io_A_Valid_5_delay_15_20 <= io_A_Valid_5_delay_14_21;
    io_A_Valid_5_delay_16_19 <= io_A_Valid_5_delay_15_20;
    io_A_Valid_5_delay_17_18 <= io_A_Valid_5_delay_16_19;
    io_A_Valid_5_delay_18_17 <= io_A_Valid_5_delay_17_18;
    io_A_Valid_5_delay_19_16 <= io_A_Valid_5_delay_18_17;
    io_A_Valid_5_delay_20_15 <= io_A_Valid_5_delay_19_16;
    io_A_Valid_5_delay_21_14 <= io_A_Valid_5_delay_20_15;
    io_A_Valid_5_delay_22_13 <= io_A_Valid_5_delay_21_14;
    io_A_Valid_5_delay_23_12 <= io_A_Valid_5_delay_22_13;
    io_A_Valid_5_delay_24_11 <= io_A_Valid_5_delay_23_12;
    io_A_Valid_5_delay_25_10 <= io_A_Valid_5_delay_24_11;
    io_A_Valid_5_delay_26_9 <= io_A_Valid_5_delay_25_10;
    io_A_Valid_5_delay_27_8 <= io_A_Valid_5_delay_26_9;
    io_A_Valid_5_delay_28_7 <= io_A_Valid_5_delay_27_8;
    io_A_Valid_5_delay_29_6 <= io_A_Valid_5_delay_28_7;
    io_A_Valid_5_delay_30_5 <= io_A_Valid_5_delay_29_6;
    io_A_Valid_5_delay_31_4 <= io_A_Valid_5_delay_30_5;
    io_A_Valid_5_delay_32_3 <= io_A_Valid_5_delay_31_4;
    io_A_Valid_5_delay_33_2 <= io_A_Valid_5_delay_32_3;
    io_A_Valid_5_delay_34_1 <= io_A_Valid_5_delay_33_2;
    io_A_Valid_5_delay_35 <= io_A_Valid_5_delay_34_1;
    io_B_Valid_35_delay_1_4 <= io_B_Valid_35;
    io_B_Valid_35_delay_2_3 <= io_B_Valid_35_delay_1_4;
    io_B_Valid_35_delay_3_2 <= io_B_Valid_35_delay_2_3;
    io_B_Valid_35_delay_4_1 <= io_B_Valid_35_delay_3_2;
    io_B_Valid_35_delay_5 <= io_B_Valid_35_delay_4_1;
    io_A_Valid_5_delay_1_35 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_34 <= io_A_Valid_5_delay_1_35;
    io_A_Valid_5_delay_3_33 <= io_A_Valid_5_delay_2_34;
    io_A_Valid_5_delay_4_32 <= io_A_Valid_5_delay_3_33;
    io_A_Valid_5_delay_5_31 <= io_A_Valid_5_delay_4_32;
    io_A_Valid_5_delay_6_30 <= io_A_Valid_5_delay_5_31;
    io_A_Valid_5_delay_7_29 <= io_A_Valid_5_delay_6_30;
    io_A_Valid_5_delay_8_28 <= io_A_Valid_5_delay_7_29;
    io_A_Valid_5_delay_9_27 <= io_A_Valid_5_delay_8_28;
    io_A_Valid_5_delay_10_26 <= io_A_Valid_5_delay_9_27;
    io_A_Valid_5_delay_11_25 <= io_A_Valid_5_delay_10_26;
    io_A_Valid_5_delay_12_24 <= io_A_Valid_5_delay_11_25;
    io_A_Valid_5_delay_13_23 <= io_A_Valid_5_delay_12_24;
    io_A_Valid_5_delay_14_22 <= io_A_Valid_5_delay_13_23;
    io_A_Valid_5_delay_15_21 <= io_A_Valid_5_delay_14_22;
    io_A_Valid_5_delay_16_20 <= io_A_Valid_5_delay_15_21;
    io_A_Valid_5_delay_17_19 <= io_A_Valid_5_delay_16_20;
    io_A_Valid_5_delay_18_18 <= io_A_Valid_5_delay_17_19;
    io_A_Valid_5_delay_19_17 <= io_A_Valid_5_delay_18_18;
    io_A_Valid_5_delay_20_16 <= io_A_Valid_5_delay_19_17;
    io_A_Valid_5_delay_21_15 <= io_A_Valid_5_delay_20_16;
    io_A_Valid_5_delay_22_14 <= io_A_Valid_5_delay_21_15;
    io_A_Valid_5_delay_23_13 <= io_A_Valid_5_delay_22_14;
    io_A_Valid_5_delay_24_12 <= io_A_Valid_5_delay_23_13;
    io_A_Valid_5_delay_25_11 <= io_A_Valid_5_delay_24_12;
    io_A_Valid_5_delay_26_10 <= io_A_Valid_5_delay_25_11;
    io_A_Valid_5_delay_27_9 <= io_A_Valid_5_delay_26_10;
    io_A_Valid_5_delay_28_8 <= io_A_Valid_5_delay_27_9;
    io_A_Valid_5_delay_29_7 <= io_A_Valid_5_delay_28_8;
    io_A_Valid_5_delay_30_6 <= io_A_Valid_5_delay_29_7;
    io_A_Valid_5_delay_31_5 <= io_A_Valid_5_delay_30_6;
    io_A_Valid_5_delay_32_4 <= io_A_Valid_5_delay_31_5;
    io_A_Valid_5_delay_33_3 <= io_A_Valid_5_delay_32_4;
    io_A_Valid_5_delay_34_2 <= io_A_Valid_5_delay_33_3;
    io_A_Valid_5_delay_35_1 <= io_A_Valid_5_delay_34_2;
    io_A_Valid_5_delay_36 <= io_A_Valid_5_delay_35_1;
    io_B_Valid_36_delay_1_4 <= io_B_Valid_36;
    io_B_Valid_36_delay_2_3 <= io_B_Valid_36_delay_1_4;
    io_B_Valid_36_delay_3_2 <= io_B_Valid_36_delay_2_3;
    io_B_Valid_36_delay_4_1 <= io_B_Valid_36_delay_3_2;
    io_B_Valid_36_delay_5 <= io_B_Valid_36_delay_4_1;
    io_A_Valid_5_delay_1_36 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_35 <= io_A_Valid_5_delay_1_36;
    io_A_Valid_5_delay_3_34 <= io_A_Valid_5_delay_2_35;
    io_A_Valid_5_delay_4_33 <= io_A_Valid_5_delay_3_34;
    io_A_Valid_5_delay_5_32 <= io_A_Valid_5_delay_4_33;
    io_A_Valid_5_delay_6_31 <= io_A_Valid_5_delay_5_32;
    io_A_Valid_5_delay_7_30 <= io_A_Valid_5_delay_6_31;
    io_A_Valid_5_delay_8_29 <= io_A_Valid_5_delay_7_30;
    io_A_Valid_5_delay_9_28 <= io_A_Valid_5_delay_8_29;
    io_A_Valid_5_delay_10_27 <= io_A_Valid_5_delay_9_28;
    io_A_Valid_5_delay_11_26 <= io_A_Valid_5_delay_10_27;
    io_A_Valid_5_delay_12_25 <= io_A_Valid_5_delay_11_26;
    io_A_Valid_5_delay_13_24 <= io_A_Valid_5_delay_12_25;
    io_A_Valid_5_delay_14_23 <= io_A_Valid_5_delay_13_24;
    io_A_Valid_5_delay_15_22 <= io_A_Valid_5_delay_14_23;
    io_A_Valid_5_delay_16_21 <= io_A_Valid_5_delay_15_22;
    io_A_Valid_5_delay_17_20 <= io_A_Valid_5_delay_16_21;
    io_A_Valid_5_delay_18_19 <= io_A_Valid_5_delay_17_20;
    io_A_Valid_5_delay_19_18 <= io_A_Valid_5_delay_18_19;
    io_A_Valid_5_delay_20_17 <= io_A_Valid_5_delay_19_18;
    io_A_Valid_5_delay_21_16 <= io_A_Valid_5_delay_20_17;
    io_A_Valid_5_delay_22_15 <= io_A_Valid_5_delay_21_16;
    io_A_Valid_5_delay_23_14 <= io_A_Valid_5_delay_22_15;
    io_A_Valid_5_delay_24_13 <= io_A_Valid_5_delay_23_14;
    io_A_Valid_5_delay_25_12 <= io_A_Valid_5_delay_24_13;
    io_A_Valid_5_delay_26_11 <= io_A_Valid_5_delay_25_12;
    io_A_Valid_5_delay_27_10 <= io_A_Valid_5_delay_26_11;
    io_A_Valid_5_delay_28_9 <= io_A_Valid_5_delay_27_10;
    io_A_Valid_5_delay_29_8 <= io_A_Valid_5_delay_28_9;
    io_A_Valid_5_delay_30_7 <= io_A_Valid_5_delay_29_8;
    io_A_Valid_5_delay_31_6 <= io_A_Valid_5_delay_30_7;
    io_A_Valid_5_delay_32_5 <= io_A_Valid_5_delay_31_6;
    io_A_Valid_5_delay_33_4 <= io_A_Valid_5_delay_32_5;
    io_A_Valid_5_delay_34_3 <= io_A_Valid_5_delay_33_4;
    io_A_Valid_5_delay_35_2 <= io_A_Valid_5_delay_34_3;
    io_A_Valid_5_delay_36_1 <= io_A_Valid_5_delay_35_2;
    io_A_Valid_5_delay_37 <= io_A_Valid_5_delay_36_1;
    io_B_Valid_37_delay_1_4 <= io_B_Valid_37;
    io_B_Valid_37_delay_2_3 <= io_B_Valid_37_delay_1_4;
    io_B_Valid_37_delay_3_2 <= io_B_Valid_37_delay_2_3;
    io_B_Valid_37_delay_4_1 <= io_B_Valid_37_delay_3_2;
    io_B_Valid_37_delay_5 <= io_B_Valid_37_delay_4_1;
    io_A_Valid_5_delay_1_37 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_36 <= io_A_Valid_5_delay_1_37;
    io_A_Valid_5_delay_3_35 <= io_A_Valid_5_delay_2_36;
    io_A_Valid_5_delay_4_34 <= io_A_Valid_5_delay_3_35;
    io_A_Valid_5_delay_5_33 <= io_A_Valid_5_delay_4_34;
    io_A_Valid_5_delay_6_32 <= io_A_Valid_5_delay_5_33;
    io_A_Valid_5_delay_7_31 <= io_A_Valid_5_delay_6_32;
    io_A_Valid_5_delay_8_30 <= io_A_Valid_5_delay_7_31;
    io_A_Valid_5_delay_9_29 <= io_A_Valid_5_delay_8_30;
    io_A_Valid_5_delay_10_28 <= io_A_Valid_5_delay_9_29;
    io_A_Valid_5_delay_11_27 <= io_A_Valid_5_delay_10_28;
    io_A_Valid_5_delay_12_26 <= io_A_Valid_5_delay_11_27;
    io_A_Valid_5_delay_13_25 <= io_A_Valid_5_delay_12_26;
    io_A_Valid_5_delay_14_24 <= io_A_Valid_5_delay_13_25;
    io_A_Valid_5_delay_15_23 <= io_A_Valid_5_delay_14_24;
    io_A_Valid_5_delay_16_22 <= io_A_Valid_5_delay_15_23;
    io_A_Valid_5_delay_17_21 <= io_A_Valid_5_delay_16_22;
    io_A_Valid_5_delay_18_20 <= io_A_Valid_5_delay_17_21;
    io_A_Valid_5_delay_19_19 <= io_A_Valid_5_delay_18_20;
    io_A_Valid_5_delay_20_18 <= io_A_Valid_5_delay_19_19;
    io_A_Valid_5_delay_21_17 <= io_A_Valid_5_delay_20_18;
    io_A_Valid_5_delay_22_16 <= io_A_Valid_5_delay_21_17;
    io_A_Valid_5_delay_23_15 <= io_A_Valid_5_delay_22_16;
    io_A_Valid_5_delay_24_14 <= io_A_Valid_5_delay_23_15;
    io_A_Valid_5_delay_25_13 <= io_A_Valid_5_delay_24_14;
    io_A_Valid_5_delay_26_12 <= io_A_Valid_5_delay_25_13;
    io_A_Valid_5_delay_27_11 <= io_A_Valid_5_delay_26_12;
    io_A_Valid_5_delay_28_10 <= io_A_Valid_5_delay_27_11;
    io_A_Valid_5_delay_29_9 <= io_A_Valid_5_delay_28_10;
    io_A_Valid_5_delay_30_8 <= io_A_Valid_5_delay_29_9;
    io_A_Valid_5_delay_31_7 <= io_A_Valid_5_delay_30_8;
    io_A_Valid_5_delay_32_6 <= io_A_Valid_5_delay_31_7;
    io_A_Valid_5_delay_33_5 <= io_A_Valid_5_delay_32_6;
    io_A_Valid_5_delay_34_4 <= io_A_Valid_5_delay_33_5;
    io_A_Valid_5_delay_35_3 <= io_A_Valid_5_delay_34_4;
    io_A_Valid_5_delay_36_2 <= io_A_Valid_5_delay_35_3;
    io_A_Valid_5_delay_37_1 <= io_A_Valid_5_delay_36_2;
    io_A_Valid_5_delay_38 <= io_A_Valid_5_delay_37_1;
    io_B_Valid_38_delay_1_4 <= io_B_Valid_38;
    io_B_Valid_38_delay_2_3 <= io_B_Valid_38_delay_1_4;
    io_B_Valid_38_delay_3_2 <= io_B_Valid_38_delay_2_3;
    io_B_Valid_38_delay_4_1 <= io_B_Valid_38_delay_3_2;
    io_B_Valid_38_delay_5 <= io_B_Valid_38_delay_4_1;
    io_A_Valid_5_delay_1_38 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_37 <= io_A_Valid_5_delay_1_38;
    io_A_Valid_5_delay_3_36 <= io_A_Valid_5_delay_2_37;
    io_A_Valid_5_delay_4_35 <= io_A_Valid_5_delay_3_36;
    io_A_Valid_5_delay_5_34 <= io_A_Valid_5_delay_4_35;
    io_A_Valid_5_delay_6_33 <= io_A_Valid_5_delay_5_34;
    io_A_Valid_5_delay_7_32 <= io_A_Valid_5_delay_6_33;
    io_A_Valid_5_delay_8_31 <= io_A_Valid_5_delay_7_32;
    io_A_Valid_5_delay_9_30 <= io_A_Valid_5_delay_8_31;
    io_A_Valid_5_delay_10_29 <= io_A_Valid_5_delay_9_30;
    io_A_Valid_5_delay_11_28 <= io_A_Valid_5_delay_10_29;
    io_A_Valid_5_delay_12_27 <= io_A_Valid_5_delay_11_28;
    io_A_Valid_5_delay_13_26 <= io_A_Valid_5_delay_12_27;
    io_A_Valid_5_delay_14_25 <= io_A_Valid_5_delay_13_26;
    io_A_Valid_5_delay_15_24 <= io_A_Valid_5_delay_14_25;
    io_A_Valid_5_delay_16_23 <= io_A_Valid_5_delay_15_24;
    io_A_Valid_5_delay_17_22 <= io_A_Valid_5_delay_16_23;
    io_A_Valid_5_delay_18_21 <= io_A_Valid_5_delay_17_22;
    io_A_Valid_5_delay_19_20 <= io_A_Valid_5_delay_18_21;
    io_A_Valid_5_delay_20_19 <= io_A_Valid_5_delay_19_20;
    io_A_Valid_5_delay_21_18 <= io_A_Valid_5_delay_20_19;
    io_A_Valid_5_delay_22_17 <= io_A_Valid_5_delay_21_18;
    io_A_Valid_5_delay_23_16 <= io_A_Valid_5_delay_22_17;
    io_A_Valid_5_delay_24_15 <= io_A_Valid_5_delay_23_16;
    io_A_Valid_5_delay_25_14 <= io_A_Valid_5_delay_24_15;
    io_A_Valid_5_delay_26_13 <= io_A_Valid_5_delay_25_14;
    io_A_Valid_5_delay_27_12 <= io_A_Valid_5_delay_26_13;
    io_A_Valid_5_delay_28_11 <= io_A_Valid_5_delay_27_12;
    io_A_Valid_5_delay_29_10 <= io_A_Valid_5_delay_28_11;
    io_A_Valid_5_delay_30_9 <= io_A_Valid_5_delay_29_10;
    io_A_Valid_5_delay_31_8 <= io_A_Valid_5_delay_30_9;
    io_A_Valid_5_delay_32_7 <= io_A_Valid_5_delay_31_8;
    io_A_Valid_5_delay_33_6 <= io_A_Valid_5_delay_32_7;
    io_A_Valid_5_delay_34_5 <= io_A_Valid_5_delay_33_6;
    io_A_Valid_5_delay_35_4 <= io_A_Valid_5_delay_34_5;
    io_A_Valid_5_delay_36_3 <= io_A_Valid_5_delay_35_4;
    io_A_Valid_5_delay_37_2 <= io_A_Valid_5_delay_36_3;
    io_A_Valid_5_delay_38_1 <= io_A_Valid_5_delay_37_2;
    io_A_Valid_5_delay_39 <= io_A_Valid_5_delay_38_1;
    io_B_Valid_39_delay_1_4 <= io_B_Valid_39;
    io_B_Valid_39_delay_2_3 <= io_B_Valid_39_delay_1_4;
    io_B_Valid_39_delay_3_2 <= io_B_Valid_39_delay_2_3;
    io_B_Valid_39_delay_4_1 <= io_B_Valid_39_delay_3_2;
    io_B_Valid_39_delay_5 <= io_B_Valid_39_delay_4_1;
    io_A_Valid_5_delay_1_39 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_38 <= io_A_Valid_5_delay_1_39;
    io_A_Valid_5_delay_3_37 <= io_A_Valid_5_delay_2_38;
    io_A_Valid_5_delay_4_36 <= io_A_Valid_5_delay_3_37;
    io_A_Valid_5_delay_5_35 <= io_A_Valid_5_delay_4_36;
    io_A_Valid_5_delay_6_34 <= io_A_Valid_5_delay_5_35;
    io_A_Valid_5_delay_7_33 <= io_A_Valid_5_delay_6_34;
    io_A_Valid_5_delay_8_32 <= io_A_Valid_5_delay_7_33;
    io_A_Valid_5_delay_9_31 <= io_A_Valid_5_delay_8_32;
    io_A_Valid_5_delay_10_30 <= io_A_Valid_5_delay_9_31;
    io_A_Valid_5_delay_11_29 <= io_A_Valid_5_delay_10_30;
    io_A_Valid_5_delay_12_28 <= io_A_Valid_5_delay_11_29;
    io_A_Valid_5_delay_13_27 <= io_A_Valid_5_delay_12_28;
    io_A_Valid_5_delay_14_26 <= io_A_Valid_5_delay_13_27;
    io_A_Valid_5_delay_15_25 <= io_A_Valid_5_delay_14_26;
    io_A_Valid_5_delay_16_24 <= io_A_Valid_5_delay_15_25;
    io_A_Valid_5_delay_17_23 <= io_A_Valid_5_delay_16_24;
    io_A_Valid_5_delay_18_22 <= io_A_Valid_5_delay_17_23;
    io_A_Valid_5_delay_19_21 <= io_A_Valid_5_delay_18_22;
    io_A_Valid_5_delay_20_20 <= io_A_Valid_5_delay_19_21;
    io_A_Valid_5_delay_21_19 <= io_A_Valid_5_delay_20_20;
    io_A_Valid_5_delay_22_18 <= io_A_Valid_5_delay_21_19;
    io_A_Valid_5_delay_23_17 <= io_A_Valid_5_delay_22_18;
    io_A_Valid_5_delay_24_16 <= io_A_Valid_5_delay_23_17;
    io_A_Valid_5_delay_25_15 <= io_A_Valid_5_delay_24_16;
    io_A_Valid_5_delay_26_14 <= io_A_Valid_5_delay_25_15;
    io_A_Valid_5_delay_27_13 <= io_A_Valid_5_delay_26_14;
    io_A_Valid_5_delay_28_12 <= io_A_Valid_5_delay_27_13;
    io_A_Valid_5_delay_29_11 <= io_A_Valid_5_delay_28_12;
    io_A_Valid_5_delay_30_10 <= io_A_Valid_5_delay_29_11;
    io_A_Valid_5_delay_31_9 <= io_A_Valid_5_delay_30_10;
    io_A_Valid_5_delay_32_8 <= io_A_Valid_5_delay_31_9;
    io_A_Valid_5_delay_33_7 <= io_A_Valid_5_delay_32_8;
    io_A_Valid_5_delay_34_6 <= io_A_Valid_5_delay_33_7;
    io_A_Valid_5_delay_35_5 <= io_A_Valid_5_delay_34_6;
    io_A_Valid_5_delay_36_4 <= io_A_Valid_5_delay_35_5;
    io_A_Valid_5_delay_37_3 <= io_A_Valid_5_delay_36_4;
    io_A_Valid_5_delay_38_2 <= io_A_Valid_5_delay_37_3;
    io_A_Valid_5_delay_39_1 <= io_A_Valid_5_delay_38_2;
    io_A_Valid_5_delay_40 <= io_A_Valid_5_delay_39_1;
    io_B_Valid_40_delay_1_4 <= io_B_Valid_40;
    io_B_Valid_40_delay_2_3 <= io_B_Valid_40_delay_1_4;
    io_B_Valid_40_delay_3_2 <= io_B_Valid_40_delay_2_3;
    io_B_Valid_40_delay_4_1 <= io_B_Valid_40_delay_3_2;
    io_B_Valid_40_delay_5 <= io_B_Valid_40_delay_4_1;
    io_A_Valid_5_delay_1_40 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_39 <= io_A_Valid_5_delay_1_40;
    io_A_Valid_5_delay_3_38 <= io_A_Valid_5_delay_2_39;
    io_A_Valid_5_delay_4_37 <= io_A_Valid_5_delay_3_38;
    io_A_Valid_5_delay_5_36 <= io_A_Valid_5_delay_4_37;
    io_A_Valid_5_delay_6_35 <= io_A_Valid_5_delay_5_36;
    io_A_Valid_5_delay_7_34 <= io_A_Valid_5_delay_6_35;
    io_A_Valid_5_delay_8_33 <= io_A_Valid_5_delay_7_34;
    io_A_Valid_5_delay_9_32 <= io_A_Valid_5_delay_8_33;
    io_A_Valid_5_delay_10_31 <= io_A_Valid_5_delay_9_32;
    io_A_Valid_5_delay_11_30 <= io_A_Valid_5_delay_10_31;
    io_A_Valid_5_delay_12_29 <= io_A_Valid_5_delay_11_30;
    io_A_Valid_5_delay_13_28 <= io_A_Valid_5_delay_12_29;
    io_A_Valid_5_delay_14_27 <= io_A_Valid_5_delay_13_28;
    io_A_Valid_5_delay_15_26 <= io_A_Valid_5_delay_14_27;
    io_A_Valid_5_delay_16_25 <= io_A_Valid_5_delay_15_26;
    io_A_Valid_5_delay_17_24 <= io_A_Valid_5_delay_16_25;
    io_A_Valid_5_delay_18_23 <= io_A_Valid_5_delay_17_24;
    io_A_Valid_5_delay_19_22 <= io_A_Valid_5_delay_18_23;
    io_A_Valid_5_delay_20_21 <= io_A_Valid_5_delay_19_22;
    io_A_Valid_5_delay_21_20 <= io_A_Valid_5_delay_20_21;
    io_A_Valid_5_delay_22_19 <= io_A_Valid_5_delay_21_20;
    io_A_Valid_5_delay_23_18 <= io_A_Valid_5_delay_22_19;
    io_A_Valid_5_delay_24_17 <= io_A_Valid_5_delay_23_18;
    io_A_Valid_5_delay_25_16 <= io_A_Valid_5_delay_24_17;
    io_A_Valid_5_delay_26_15 <= io_A_Valid_5_delay_25_16;
    io_A_Valid_5_delay_27_14 <= io_A_Valid_5_delay_26_15;
    io_A_Valid_5_delay_28_13 <= io_A_Valid_5_delay_27_14;
    io_A_Valid_5_delay_29_12 <= io_A_Valid_5_delay_28_13;
    io_A_Valid_5_delay_30_11 <= io_A_Valid_5_delay_29_12;
    io_A_Valid_5_delay_31_10 <= io_A_Valid_5_delay_30_11;
    io_A_Valid_5_delay_32_9 <= io_A_Valid_5_delay_31_10;
    io_A_Valid_5_delay_33_8 <= io_A_Valid_5_delay_32_9;
    io_A_Valid_5_delay_34_7 <= io_A_Valid_5_delay_33_8;
    io_A_Valid_5_delay_35_6 <= io_A_Valid_5_delay_34_7;
    io_A_Valid_5_delay_36_5 <= io_A_Valid_5_delay_35_6;
    io_A_Valid_5_delay_37_4 <= io_A_Valid_5_delay_36_5;
    io_A_Valid_5_delay_38_3 <= io_A_Valid_5_delay_37_4;
    io_A_Valid_5_delay_39_2 <= io_A_Valid_5_delay_38_3;
    io_A_Valid_5_delay_40_1 <= io_A_Valid_5_delay_39_2;
    io_A_Valid_5_delay_41 <= io_A_Valid_5_delay_40_1;
    io_B_Valid_41_delay_1_4 <= io_B_Valid_41;
    io_B_Valid_41_delay_2_3 <= io_B_Valid_41_delay_1_4;
    io_B_Valid_41_delay_3_2 <= io_B_Valid_41_delay_2_3;
    io_B_Valid_41_delay_4_1 <= io_B_Valid_41_delay_3_2;
    io_B_Valid_41_delay_5 <= io_B_Valid_41_delay_4_1;
    io_A_Valid_5_delay_1_41 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_40 <= io_A_Valid_5_delay_1_41;
    io_A_Valid_5_delay_3_39 <= io_A_Valid_5_delay_2_40;
    io_A_Valid_5_delay_4_38 <= io_A_Valid_5_delay_3_39;
    io_A_Valid_5_delay_5_37 <= io_A_Valid_5_delay_4_38;
    io_A_Valid_5_delay_6_36 <= io_A_Valid_5_delay_5_37;
    io_A_Valid_5_delay_7_35 <= io_A_Valid_5_delay_6_36;
    io_A_Valid_5_delay_8_34 <= io_A_Valid_5_delay_7_35;
    io_A_Valid_5_delay_9_33 <= io_A_Valid_5_delay_8_34;
    io_A_Valid_5_delay_10_32 <= io_A_Valid_5_delay_9_33;
    io_A_Valid_5_delay_11_31 <= io_A_Valid_5_delay_10_32;
    io_A_Valid_5_delay_12_30 <= io_A_Valid_5_delay_11_31;
    io_A_Valid_5_delay_13_29 <= io_A_Valid_5_delay_12_30;
    io_A_Valid_5_delay_14_28 <= io_A_Valid_5_delay_13_29;
    io_A_Valid_5_delay_15_27 <= io_A_Valid_5_delay_14_28;
    io_A_Valid_5_delay_16_26 <= io_A_Valid_5_delay_15_27;
    io_A_Valid_5_delay_17_25 <= io_A_Valid_5_delay_16_26;
    io_A_Valid_5_delay_18_24 <= io_A_Valid_5_delay_17_25;
    io_A_Valid_5_delay_19_23 <= io_A_Valid_5_delay_18_24;
    io_A_Valid_5_delay_20_22 <= io_A_Valid_5_delay_19_23;
    io_A_Valid_5_delay_21_21 <= io_A_Valid_5_delay_20_22;
    io_A_Valid_5_delay_22_20 <= io_A_Valid_5_delay_21_21;
    io_A_Valid_5_delay_23_19 <= io_A_Valid_5_delay_22_20;
    io_A_Valid_5_delay_24_18 <= io_A_Valid_5_delay_23_19;
    io_A_Valid_5_delay_25_17 <= io_A_Valid_5_delay_24_18;
    io_A_Valid_5_delay_26_16 <= io_A_Valid_5_delay_25_17;
    io_A_Valid_5_delay_27_15 <= io_A_Valid_5_delay_26_16;
    io_A_Valid_5_delay_28_14 <= io_A_Valid_5_delay_27_15;
    io_A_Valid_5_delay_29_13 <= io_A_Valid_5_delay_28_14;
    io_A_Valid_5_delay_30_12 <= io_A_Valid_5_delay_29_13;
    io_A_Valid_5_delay_31_11 <= io_A_Valid_5_delay_30_12;
    io_A_Valid_5_delay_32_10 <= io_A_Valid_5_delay_31_11;
    io_A_Valid_5_delay_33_9 <= io_A_Valid_5_delay_32_10;
    io_A_Valid_5_delay_34_8 <= io_A_Valid_5_delay_33_9;
    io_A_Valid_5_delay_35_7 <= io_A_Valid_5_delay_34_8;
    io_A_Valid_5_delay_36_6 <= io_A_Valid_5_delay_35_7;
    io_A_Valid_5_delay_37_5 <= io_A_Valid_5_delay_36_6;
    io_A_Valid_5_delay_38_4 <= io_A_Valid_5_delay_37_5;
    io_A_Valid_5_delay_39_3 <= io_A_Valid_5_delay_38_4;
    io_A_Valid_5_delay_40_2 <= io_A_Valid_5_delay_39_3;
    io_A_Valid_5_delay_41_1 <= io_A_Valid_5_delay_40_2;
    io_A_Valid_5_delay_42 <= io_A_Valid_5_delay_41_1;
    io_B_Valid_42_delay_1_4 <= io_B_Valid_42;
    io_B_Valid_42_delay_2_3 <= io_B_Valid_42_delay_1_4;
    io_B_Valid_42_delay_3_2 <= io_B_Valid_42_delay_2_3;
    io_B_Valid_42_delay_4_1 <= io_B_Valid_42_delay_3_2;
    io_B_Valid_42_delay_5 <= io_B_Valid_42_delay_4_1;
    io_A_Valid_5_delay_1_42 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_41 <= io_A_Valid_5_delay_1_42;
    io_A_Valid_5_delay_3_40 <= io_A_Valid_5_delay_2_41;
    io_A_Valid_5_delay_4_39 <= io_A_Valid_5_delay_3_40;
    io_A_Valid_5_delay_5_38 <= io_A_Valid_5_delay_4_39;
    io_A_Valid_5_delay_6_37 <= io_A_Valid_5_delay_5_38;
    io_A_Valid_5_delay_7_36 <= io_A_Valid_5_delay_6_37;
    io_A_Valid_5_delay_8_35 <= io_A_Valid_5_delay_7_36;
    io_A_Valid_5_delay_9_34 <= io_A_Valid_5_delay_8_35;
    io_A_Valid_5_delay_10_33 <= io_A_Valid_5_delay_9_34;
    io_A_Valid_5_delay_11_32 <= io_A_Valid_5_delay_10_33;
    io_A_Valid_5_delay_12_31 <= io_A_Valid_5_delay_11_32;
    io_A_Valid_5_delay_13_30 <= io_A_Valid_5_delay_12_31;
    io_A_Valid_5_delay_14_29 <= io_A_Valid_5_delay_13_30;
    io_A_Valid_5_delay_15_28 <= io_A_Valid_5_delay_14_29;
    io_A_Valid_5_delay_16_27 <= io_A_Valid_5_delay_15_28;
    io_A_Valid_5_delay_17_26 <= io_A_Valid_5_delay_16_27;
    io_A_Valid_5_delay_18_25 <= io_A_Valid_5_delay_17_26;
    io_A_Valid_5_delay_19_24 <= io_A_Valid_5_delay_18_25;
    io_A_Valid_5_delay_20_23 <= io_A_Valid_5_delay_19_24;
    io_A_Valid_5_delay_21_22 <= io_A_Valid_5_delay_20_23;
    io_A_Valid_5_delay_22_21 <= io_A_Valid_5_delay_21_22;
    io_A_Valid_5_delay_23_20 <= io_A_Valid_5_delay_22_21;
    io_A_Valid_5_delay_24_19 <= io_A_Valid_5_delay_23_20;
    io_A_Valid_5_delay_25_18 <= io_A_Valid_5_delay_24_19;
    io_A_Valid_5_delay_26_17 <= io_A_Valid_5_delay_25_18;
    io_A_Valid_5_delay_27_16 <= io_A_Valid_5_delay_26_17;
    io_A_Valid_5_delay_28_15 <= io_A_Valid_5_delay_27_16;
    io_A_Valid_5_delay_29_14 <= io_A_Valid_5_delay_28_15;
    io_A_Valid_5_delay_30_13 <= io_A_Valid_5_delay_29_14;
    io_A_Valid_5_delay_31_12 <= io_A_Valid_5_delay_30_13;
    io_A_Valid_5_delay_32_11 <= io_A_Valid_5_delay_31_12;
    io_A_Valid_5_delay_33_10 <= io_A_Valid_5_delay_32_11;
    io_A_Valid_5_delay_34_9 <= io_A_Valid_5_delay_33_10;
    io_A_Valid_5_delay_35_8 <= io_A_Valid_5_delay_34_9;
    io_A_Valid_5_delay_36_7 <= io_A_Valid_5_delay_35_8;
    io_A_Valid_5_delay_37_6 <= io_A_Valid_5_delay_36_7;
    io_A_Valid_5_delay_38_5 <= io_A_Valid_5_delay_37_6;
    io_A_Valid_5_delay_39_4 <= io_A_Valid_5_delay_38_5;
    io_A_Valid_5_delay_40_3 <= io_A_Valid_5_delay_39_4;
    io_A_Valid_5_delay_41_2 <= io_A_Valid_5_delay_40_3;
    io_A_Valid_5_delay_42_1 <= io_A_Valid_5_delay_41_2;
    io_A_Valid_5_delay_43 <= io_A_Valid_5_delay_42_1;
    io_B_Valid_43_delay_1_4 <= io_B_Valid_43;
    io_B_Valid_43_delay_2_3 <= io_B_Valid_43_delay_1_4;
    io_B_Valid_43_delay_3_2 <= io_B_Valid_43_delay_2_3;
    io_B_Valid_43_delay_4_1 <= io_B_Valid_43_delay_3_2;
    io_B_Valid_43_delay_5 <= io_B_Valid_43_delay_4_1;
    io_A_Valid_5_delay_1_43 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_42 <= io_A_Valid_5_delay_1_43;
    io_A_Valid_5_delay_3_41 <= io_A_Valid_5_delay_2_42;
    io_A_Valid_5_delay_4_40 <= io_A_Valid_5_delay_3_41;
    io_A_Valid_5_delay_5_39 <= io_A_Valid_5_delay_4_40;
    io_A_Valid_5_delay_6_38 <= io_A_Valid_5_delay_5_39;
    io_A_Valid_5_delay_7_37 <= io_A_Valid_5_delay_6_38;
    io_A_Valid_5_delay_8_36 <= io_A_Valid_5_delay_7_37;
    io_A_Valid_5_delay_9_35 <= io_A_Valid_5_delay_8_36;
    io_A_Valid_5_delay_10_34 <= io_A_Valid_5_delay_9_35;
    io_A_Valid_5_delay_11_33 <= io_A_Valid_5_delay_10_34;
    io_A_Valid_5_delay_12_32 <= io_A_Valid_5_delay_11_33;
    io_A_Valid_5_delay_13_31 <= io_A_Valid_5_delay_12_32;
    io_A_Valid_5_delay_14_30 <= io_A_Valid_5_delay_13_31;
    io_A_Valid_5_delay_15_29 <= io_A_Valid_5_delay_14_30;
    io_A_Valid_5_delay_16_28 <= io_A_Valid_5_delay_15_29;
    io_A_Valid_5_delay_17_27 <= io_A_Valid_5_delay_16_28;
    io_A_Valid_5_delay_18_26 <= io_A_Valid_5_delay_17_27;
    io_A_Valid_5_delay_19_25 <= io_A_Valid_5_delay_18_26;
    io_A_Valid_5_delay_20_24 <= io_A_Valid_5_delay_19_25;
    io_A_Valid_5_delay_21_23 <= io_A_Valid_5_delay_20_24;
    io_A_Valid_5_delay_22_22 <= io_A_Valid_5_delay_21_23;
    io_A_Valid_5_delay_23_21 <= io_A_Valid_5_delay_22_22;
    io_A_Valid_5_delay_24_20 <= io_A_Valid_5_delay_23_21;
    io_A_Valid_5_delay_25_19 <= io_A_Valid_5_delay_24_20;
    io_A_Valid_5_delay_26_18 <= io_A_Valid_5_delay_25_19;
    io_A_Valid_5_delay_27_17 <= io_A_Valid_5_delay_26_18;
    io_A_Valid_5_delay_28_16 <= io_A_Valid_5_delay_27_17;
    io_A_Valid_5_delay_29_15 <= io_A_Valid_5_delay_28_16;
    io_A_Valid_5_delay_30_14 <= io_A_Valid_5_delay_29_15;
    io_A_Valid_5_delay_31_13 <= io_A_Valid_5_delay_30_14;
    io_A_Valid_5_delay_32_12 <= io_A_Valid_5_delay_31_13;
    io_A_Valid_5_delay_33_11 <= io_A_Valid_5_delay_32_12;
    io_A_Valid_5_delay_34_10 <= io_A_Valid_5_delay_33_11;
    io_A_Valid_5_delay_35_9 <= io_A_Valid_5_delay_34_10;
    io_A_Valid_5_delay_36_8 <= io_A_Valid_5_delay_35_9;
    io_A_Valid_5_delay_37_7 <= io_A_Valid_5_delay_36_8;
    io_A_Valid_5_delay_38_6 <= io_A_Valid_5_delay_37_7;
    io_A_Valid_5_delay_39_5 <= io_A_Valid_5_delay_38_6;
    io_A_Valid_5_delay_40_4 <= io_A_Valid_5_delay_39_5;
    io_A_Valid_5_delay_41_3 <= io_A_Valid_5_delay_40_4;
    io_A_Valid_5_delay_42_2 <= io_A_Valid_5_delay_41_3;
    io_A_Valid_5_delay_43_1 <= io_A_Valid_5_delay_42_2;
    io_A_Valid_5_delay_44 <= io_A_Valid_5_delay_43_1;
    io_B_Valid_44_delay_1_4 <= io_B_Valid_44;
    io_B_Valid_44_delay_2_3 <= io_B_Valid_44_delay_1_4;
    io_B_Valid_44_delay_3_2 <= io_B_Valid_44_delay_2_3;
    io_B_Valid_44_delay_4_1 <= io_B_Valid_44_delay_3_2;
    io_B_Valid_44_delay_5 <= io_B_Valid_44_delay_4_1;
    io_A_Valid_5_delay_1_44 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_43 <= io_A_Valid_5_delay_1_44;
    io_A_Valid_5_delay_3_42 <= io_A_Valid_5_delay_2_43;
    io_A_Valid_5_delay_4_41 <= io_A_Valid_5_delay_3_42;
    io_A_Valid_5_delay_5_40 <= io_A_Valid_5_delay_4_41;
    io_A_Valid_5_delay_6_39 <= io_A_Valid_5_delay_5_40;
    io_A_Valid_5_delay_7_38 <= io_A_Valid_5_delay_6_39;
    io_A_Valid_5_delay_8_37 <= io_A_Valid_5_delay_7_38;
    io_A_Valid_5_delay_9_36 <= io_A_Valid_5_delay_8_37;
    io_A_Valid_5_delay_10_35 <= io_A_Valid_5_delay_9_36;
    io_A_Valid_5_delay_11_34 <= io_A_Valid_5_delay_10_35;
    io_A_Valid_5_delay_12_33 <= io_A_Valid_5_delay_11_34;
    io_A_Valid_5_delay_13_32 <= io_A_Valid_5_delay_12_33;
    io_A_Valid_5_delay_14_31 <= io_A_Valid_5_delay_13_32;
    io_A_Valid_5_delay_15_30 <= io_A_Valid_5_delay_14_31;
    io_A_Valid_5_delay_16_29 <= io_A_Valid_5_delay_15_30;
    io_A_Valid_5_delay_17_28 <= io_A_Valid_5_delay_16_29;
    io_A_Valid_5_delay_18_27 <= io_A_Valid_5_delay_17_28;
    io_A_Valid_5_delay_19_26 <= io_A_Valid_5_delay_18_27;
    io_A_Valid_5_delay_20_25 <= io_A_Valid_5_delay_19_26;
    io_A_Valid_5_delay_21_24 <= io_A_Valid_5_delay_20_25;
    io_A_Valid_5_delay_22_23 <= io_A_Valid_5_delay_21_24;
    io_A_Valid_5_delay_23_22 <= io_A_Valid_5_delay_22_23;
    io_A_Valid_5_delay_24_21 <= io_A_Valid_5_delay_23_22;
    io_A_Valid_5_delay_25_20 <= io_A_Valid_5_delay_24_21;
    io_A_Valid_5_delay_26_19 <= io_A_Valid_5_delay_25_20;
    io_A_Valid_5_delay_27_18 <= io_A_Valid_5_delay_26_19;
    io_A_Valid_5_delay_28_17 <= io_A_Valid_5_delay_27_18;
    io_A_Valid_5_delay_29_16 <= io_A_Valid_5_delay_28_17;
    io_A_Valid_5_delay_30_15 <= io_A_Valid_5_delay_29_16;
    io_A_Valid_5_delay_31_14 <= io_A_Valid_5_delay_30_15;
    io_A_Valid_5_delay_32_13 <= io_A_Valid_5_delay_31_14;
    io_A_Valid_5_delay_33_12 <= io_A_Valid_5_delay_32_13;
    io_A_Valid_5_delay_34_11 <= io_A_Valid_5_delay_33_12;
    io_A_Valid_5_delay_35_10 <= io_A_Valid_5_delay_34_11;
    io_A_Valid_5_delay_36_9 <= io_A_Valid_5_delay_35_10;
    io_A_Valid_5_delay_37_8 <= io_A_Valid_5_delay_36_9;
    io_A_Valid_5_delay_38_7 <= io_A_Valid_5_delay_37_8;
    io_A_Valid_5_delay_39_6 <= io_A_Valid_5_delay_38_7;
    io_A_Valid_5_delay_40_5 <= io_A_Valid_5_delay_39_6;
    io_A_Valid_5_delay_41_4 <= io_A_Valid_5_delay_40_5;
    io_A_Valid_5_delay_42_3 <= io_A_Valid_5_delay_41_4;
    io_A_Valid_5_delay_43_2 <= io_A_Valid_5_delay_42_3;
    io_A_Valid_5_delay_44_1 <= io_A_Valid_5_delay_43_2;
    io_A_Valid_5_delay_45 <= io_A_Valid_5_delay_44_1;
    io_B_Valid_45_delay_1_4 <= io_B_Valid_45;
    io_B_Valid_45_delay_2_3 <= io_B_Valid_45_delay_1_4;
    io_B_Valid_45_delay_3_2 <= io_B_Valid_45_delay_2_3;
    io_B_Valid_45_delay_4_1 <= io_B_Valid_45_delay_3_2;
    io_B_Valid_45_delay_5 <= io_B_Valid_45_delay_4_1;
    io_A_Valid_5_delay_1_45 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_44 <= io_A_Valid_5_delay_1_45;
    io_A_Valid_5_delay_3_43 <= io_A_Valid_5_delay_2_44;
    io_A_Valid_5_delay_4_42 <= io_A_Valid_5_delay_3_43;
    io_A_Valid_5_delay_5_41 <= io_A_Valid_5_delay_4_42;
    io_A_Valid_5_delay_6_40 <= io_A_Valid_5_delay_5_41;
    io_A_Valid_5_delay_7_39 <= io_A_Valid_5_delay_6_40;
    io_A_Valid_5_delay_8_38 <= io_A_Valid_5_delay_7_39;
    io_A_Valid_5_delay_9_37 <= io_A_Valid_5_delay_8_38;
    io_A_Valid_5_delay_10_36 <= io_A_Valid_5_delay_9_37;
    io_A_Valid_5_delay_11_35 <= io_A_Valid_5_delay_10_36;
    io_A_Valid_5_delay_12_34 <= io_A_Valid_5_delay_11_35;
    io_A_Valid_5_delay_13_33 <= io_A_Valid_5_delay_12_34;
    io_A_Valid_5_delay_14_32 <= io_A_Valid_5_delay_13_33;
    io_A_Valid_5_delay_15_31 <= io_A_Valid_5_delay_14_32;
    io_A_Valid_5_delay_16_30 <= io_A_Valid_5_delay_15_31;
    io_A_Valid_5_delay_17_29 <= io_A_Valid_5_delay_16_30;
    io_A_Valid_5_delay_18_28 <= io_A_Valid_5_delay_17_29;
    io_A_Valid_5_delay_19_27 <= io_A_Valid_5_delay_18_28;
    io_A_Valid_5_delay_20_26 <= io_A_Valid_5_delay_19_27;
    io_A_Valid_5_delay_21_25 <= io_A_Valid_5_delay_20_26;
    io_A_Valid_5_delay_22_24 <= io_A_Valid_5_delay_21_25;
    io_A_Valid_5_delay_23_23 <= io_A_Valid_5_delay_22_24;
    io_A_Valid_5_delay_24_22 <= io_A_Valid_5_delay_23_23;
    io_A_Valid_5_delay_25_21 <= io_A_Valid_5_delay_24_22;
    io_A_Valid_5_delay_26_20 <= io_A_Valid_5_delay_25_21;
    io_A_Valid_5_delay_27_19 <= io_A_Valid_5_delay_26_20;
    io_A_Valid_5_delay_28_18 <= io_A_Valid_5_delay_27_19;
    io_A_Valid_5_delay_29_17 <= io_A_Valid_5_delay_28_18;
    io_A_Valid_5_delay_30_16 <= io_A_Valid_5_delay_29_17;
    io_A_Valid_5_delay_31_15 <= io_A_Valid_5_delay_30_16;
    io_A_Valid_5_delay_32_14 <= io_A_Valid_5_delay_31_15;
    io_A_Valid_5_delay_33_13 <= io_A_Valid_5_delay_32_14;
    io_A_Valid_5_delay_34_12 <= io_A_Valid_5_delay_33_13;
    io_A_Valid_5_delay_35_11 <= io_A_Valid_5_delay_34_12;
    io_A_Valid_5_delay_36_10 <= io_A_Valid_5_delay_35_11;
    io_A_Valid_5_delay_37_9 <= io_A_Valid_5_delay_36_10;
    io_A_Valid_5_delay_38_8 <= io_A_Valid_5_delay_37_9;
    io_A_Valid_5_delay_39_7 <= io_A_Valid_5_delay_38_8;
    io_A_Valid_5_delay_40_6 <= io_A_Valid_5_delay_39_7;
    io_A_Valid_5_delay_41_5 <= io_A_Valid_5_delay_40_6;
    io_A_Valid_5_delay_42_4 <= io_A_Valid_5_delay_41_5;
    io_A_Valid_5_delay_43_3 <= io_A_Valid_5_delay_42_4;
    io_A_Valid_5_delay_44_2 <= io_A_Valid_5_delay_43_3;
    io_A_Valid_5_delay_45_1 <= io_A_Valid_5_delay_44_2;
    io_A_Valid_5_delay_46 <= io_A_Valid_5_delay_45_1;
    io_B_Valid_46_delay_1_4 <= io_B_Valid_46;
    io_B_Valid_46_delay_2_3 <= io_B_Valid_46_delay_1_4;
    io_B_Valid_46_delay_3_2 <= io_B_Valid_46_delay_2_3;
    io_B_Valid_46_delay_4_1 <= io_B_Valid_46_delay_3_2;
    io_B_Valid_46_delay_5 <= io_B_Valid_46_delay_4_1;
    io_A_Valid_5_delay_1_46 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_45 <= io_A_Valid_5_delay_1_46;
    io_A_Valid_5_delay_3_44 <= io_A_Valid_5_delay_2_45;
    io_A_Valid_5_delay_4_43 <= io_A_Valid_5_delay_3_44;
    io_A_Valid_5_delay_5_42 <= io_A_Valid_5_delay_4_43;
    io_A_Valid_5_delay_6_41 <= io_A_Valid_5_delay_5_42;
    io_A_Valid_5_delay_7_40 <= io_A_Valid_5_delay_6_41;
    io_A_Valid_5_delay_8_39 <= io_A_Valid_5_delay_7_40;
    io_A_Valid_5_delay_9_38 <= io_A_Valid_5_delay_8_39;
    io_A_Valid_5_delay_10_37 <= io_A_Valid_5_delay_9_38;
    io_A_Valid_5_delay_11_36 <= io_A_Valid_5_delay_10_37;
    io_A_Valid_5_delay_12_35 <= io_A_Valid_5_delay_11_36;
    io_A_Valid_5_delay_13_34 <= io_A_Valid_5_delay_12_35;
    io_A_Valid_5_delay_14_33 <= io_A_Valid_5_delay_13_34;
    io_A_Valid_5_delay_15_32 <= io_A_Valid_5_delay_14_33;
    io_A_Valid_5_delay_16_31 <= io_A_Valid_5_delay_15_32;
    io_A_Valid_5_delay_17_30 <= io_A_Valid_5_delay_16_31;
    io_A_Valid_5_delay_18_29 <= io_A_Valid_5_delay_17_30;
    io_A_Valid_5_delay_19_28 <= io_A_Valid_5_delay_18_29;
    io_A_Valid_5_delay_20_27 <= io_A_Valid_5_delay_19_28;
    io_A_Valid_5_delay_21_26 <= io_A_Valid_5_delay_20_27;
    io_A_Valid_5_delay_22_25 <= io_A_Valid_5_delay_21_26;
    io_A_Valid_5_delay_23_24 <= io_A_Valid_5_delay_22_25;
    io_A_Valid_5_delay_24_23 <= io_A_Valid_5_delay_23_24;
    io_A_Valid_5_delay_25_22 <= io_A_Valid_5_delay_24_23;
    io_A_Valid_5_delay_26_21 <= io_A_Valid_5_delay_25_22;
    io_A_Valid_5_delay_27_20 <= io_A_Valid_5_delay_26_21;
    io_A_Valid_5_delay_28_19 <= io_A_Valid_5_delay_27_20;
    io_A_Valid_5_delay_29_18 <= io_A_Valid_5_delay_28_19;
    io_A_Valid_5_delay_30_17 <= io_A_Valid_5_delay_29_18;
    io_A_Valid_5_delay_31_16 <= io_A_Valid_5_delay_30_17;
    io_A_Valid_5_delay_32_15 <= io_A_Valid_5_delay_31_16;
    io_A_Valid_5_delay_33_14 <= io_A_Valid_5_delay_32_15;
    io_A_Valid_5_delay_34_13 <= io_A_Valid_5_delay_33_14;
    io_A_Valid_5_delay_35_12 <= io_A_Valid_5_delay_34_13;
    io_A_Valid_5_delay_36_11 <= io_A_Valid_5_delay_35_12;
    io_A_Valid_5_delay_37_10 <= io_A_Valid_5_delay_36_11;
    io_A_Valid_5_delay_38_9 <= io_A_Valid_5_delay_37_10;
    io_A_Valid_5_delay_39_8 <= io_A_Valid_5_delay_38_9;
    io_A_Valid_5_delay_40_7 <= io_A_Valid_5_delay_39_8;
    io_A_Valid_5_delay_41_6 <= io_A_Valid_5_delay_40_7;
    io_A_Valid_5_delay_42_5 <= io_A_Valid_5_delay_41_6;
    io_A_Valid_5_delay_43_4 <= io_A_Valid_5_delay_42_5;
    io_A_Valid_5_delay_44_3 <= io_A_Valid_5_delay_43_4;
    io_A_Valid_5_delay_45_2 <= io_A_Valid_5_delay_44_3;
    io_A_Valid_5_delay_46_1 <= io_A_Valid_5_delay_45_2;
    io_A_Valid_5_delay_47 <= io_A_Valid_5_delay_46_1;
    io_B_Valid_47_delay_1_4 <= io_B_Valid_47;
    io_B_Valid_47_delay_2_3 <= io_B_Valid_47_delay_1_4;
    io_B_Valid_47_delay_3_2 <= io_B_Valid_47_delay_2_3;
    io_B_Valid_47_delay_4_1 <= io_B_Valid_47_delay_3_2;
    io_B_Valid_47_delay_5 <= io_B_Valid_47_delay_4_1;
    io_A_Valid_5_delay_1_47 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_46 <= io_A_Valid_5_delay_1_47;
    io_A_Valid_5_delay_3_45 <= io_A_Valid_5_delay_2_46;
    io_A_Valid_5_delay_4_44 <= io_A_Valid_5_delay_3_45;
    io_A_Valid_5_delay_5_43 <= io_A_Valid_5_delay_4_44;
    io_A_Valid_5_delay_6_42 <= io_A_Valid_5_delay_5_43;
    io_A_Valid_5_delay_7_41 <= io_A_Valid_5_delay_6_42;
    io_A_Valid_5_delay_8_40 <= io_A_Valid_5_delay_7_41;
    io_A_Valid_5_delay_9_39 <= io_A_Valid_5_delay_8_40;
    io_A_Valid_5_delay_10_38 <= io_A_Valid_5_delay_9_39;
    io_A_Valid_5_delay_11_37 <= io_A_Valid_5_delay_10_38;
    io_A_Valid_5_delay_12_36 <= io_A_Valid_5_delay_11_37;
    io_A_Valid_5_delay_13_35 <= io_A_Valid_5_delay_12_36;
    io_A_Valid_5_delay_14_34 <= io_A_Valid_5_delay_13_35;
    io_A_Valid_5_delay_15_33 <= io_A_Valid_5_delay_14_34;
    io_A_Valid_5_delay_16_32 <= io_A_Valid_5_delay_15_33;
    io_A_Valid_5_delay_17_31 <= io_A_Valid_5_delay_16_32;
    io_A_Valid_5_delay_18_30 <= io_A_Valid_5_delay_17_31;
    io_A_Valid_5_delay_19_29 <= io_A_Valid_5_delay_18_30;
    io_A_Valid_5_delay_20_28 <= io_A_Valid_5_delay_19_29;
    io_A_Valid_5_delay_21_27 <= io_A_Valid_5_delay_20_28;
    io_A_Valid_5_delay_22_26 <= io_A_Valid_5_delay_21_27;
    io_A_Valid_5_delay_23_25 <= io_A_Valid_5_delay_22_26;
    io_A_Valid_5_delay_24_24 <= io_A_Valid_5_delay_23_25;
    io_A_Valid_5_delay_25_23 <= io_A_Valid_5_delay_24_24;
    io_A_Valid_5_delay_26_22 <= io_A_Valid_5_delay_25_23;
    io_A_Valid_5_delay_27_21 <= io_A_Valid_5_delay_26_22;
    io_A_Valid_5_delay_28_20 <= io_A_Valid_5_delay_27_21;
    io_A_Valid_5_delay_29_19 <= io_A_Valid_5_delay_28_20;
    io_A_Valid_5_delay_30_18 <= io_A_Valid_5_delay_29_19;
    io_A_Valid_5_delay_31_17 <= io_A_Valid_5_delay_30_18;
    io_A_Valid_5_delay_32_16 <= io_A_Valid_5_delay_31_17;
    io_A_Valid_5_delay_33_15 <= io_A_Valid_5_delay_32_16;
    io_A_Valid_5_delay_34_14 <= io_A_Valid_5_delay_33_15;
    io_A_Valid_5_delay_35_13 <= io_A_Valid_5_delay_34_14;
    io_A_Valid_5_delay_36_12 <= io_A_Valid_5_delay_35_13;
    io_A_Valid_5_delay_37_11 <= io_A_Valid_5_delay_36_12;
    io_A_Valid_5_delay_38_10 <= io_A_Valid_5_delay_37_11;
    io_A_Valid_5_delay_39_9 <= io_A_Valid_5_delay_38_10;
    io_A_Valid_5_delay_40_8 <= io_A_Valid_5_delay_39_9;
    io_A_Valid_5_delay_41_7 <= io_A_Valid_5_delay_40_8;
    io_A_Valid_5_delay_42_6 <= io_A_Valid_5_delay_41_7;
    io_A_Valid_5_delay_43_5 <= io_A_Valid_5_delay_42_6;
    io_A_Valid_5_delay_44_4 <= io_A_Valid_5_delay_43_5;
    io_A_Valid_5_delay_45_3 <= io_A_Valid_5_delay_44_4;
    io_A_Valid_5_delay_46_2 <= io_A_Valid_5_delay_45_3;
    io_A_Valid_5_delay_47_1 <= io_A_Valid_5_delay_46_2;
    io_A_Valid_5_delay_48 <= io_A_Valid_5_delay_47_1;
    io_B_Valid_48_delay_1_4 <= io_B_Valid_48;
    io_B_Valid_48_delay_2_3 <= io_B_Valid_48_delay_1_4;
    io_B_Valid_48_delay_3_2 <= io_B_Valid_48_delay_2_3;
    io_B_Valid_48_delay_4_1 <= io_B_Valid_48_delay_3_2;
    io_B_Valid_48_delay_5 <= io_B_Valid_48_delay_4_1;
    io_A_Valid_5_delay_1_48 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_47 <= io_A_Valid_5_delay_1_48;
    io_A_Valid_5_delay_3_46 <= io_A_Valid_5_delay_2_47;
    io_A_Valid_5_delay_4_45 <= io_A_Valid_5_delay_3_46;
    io_A_Valid_5_delay_5_44 <= io_A_Valid_5_delay_4_45;
    io_A_Valid_5_delay_6_43 <= io_A_Valid_5_delay_5_44;
    io_A_Valid_5_delay_7_42 <= io_A_Valid_5_delay_6_43;
    io_A_Valid_5_delay_8_41 <= io_A_Valid_5_delay_7_42;
    io_A_Valid_5_delay_9_40 <= io_A_Valid_5_delay_8_41;
    io_A_Valid_5_delay_10_39 <= io_A_Valid_5_delay_9_40;
    io_A_Valid_5_delay_11_38 <= io_A_Valid_5_delay_10_39;
    io_A_Valid_5_delay_12_37 <= io_A_Valid_5_delay_11_38;
    io_A_Valid_5_delay_13_36 <= io_A_Valid_5_delay_12_37;
    io_A_Valid_5_delay_14_35 <= io_A_Valid_5_delay_13_36;
    io_A_Valid_5_delay_15_34 <= io_A_Valid_5_delay_14_35;
    io_A_Valid_5_delay_16_33 <= io_A_Valid_5_delay_15_34;
    io_A_Valid_5_delay_17_32 <= io_A_Valid_5_delay_16_33;
    io_A_Valid_5_delay_18_31 <= io_A_Valid_5_delay_17_32;
    io_A_Valid_5_delay_19_30 <= io_A_Valid_5_delay_18_31;
    io_A_Valid_5_delay_20_29 <= io_A_Valid_5_delay_19_30;
    io_A_Valid_5_delay_21_28 <= io_A_Valid_5_delay_20_29;
    io_A_Valid_5_delay_22_27 <= io_A_Valid_5_delay_21_28;
    io_A_Valid_5_delay_23_26 <= io_A_Valid_5_delay_22_27;
    io_A_Valid_5_delay_24_25 <= io_A_Valid_5_delay_23_26;
    io_A_Valid_5_delay_25_24 <= io_A_Valid_5_delay_24_25;
    io_A_Valid_5_delay_26_23 <= io_A_Valid_5_delay_25_24;
    io_A_Valid_5_delay_27_22 <= io_A_Valid_5_delay_26_23;
    io_A_Valid_5_delay_28_21 <= io_A_Valid_5_delay_27_22;
    io_A_Valid_5_delay_29_20 <= io_A_Valid_5_delay_28_21;
    io_A_Valid_5_delay_30_19 <= io_A_Valid_5_delay_29_20;
    io_A_Valid_5_delay_31_18 <= io_A_Valid_5_delay_30_19;
    io_A_Valid_5_delay_32_17 <= io_A_Valid_5_delay_31_18;
    io_A_Valid_5_delay_33_16 <= io_A_Valid_5_delay_32_17;
    io_A_Valid_5_delay_34_15 <= io_A_Valid_5_delay_33_16;
    io_A_Valid_5_delay_35_14 <= io_A_Valid_5_delay_34_15;
    io_A_Valid_5_delay_36_13 <= io_A_Valid_5_delay_35_14;
    io_A_Valid_5_delay_37_12 <= io_A_Valid_5_delay_36_13;
    io_A_Valid_5_delay_38_11 <= io_A_Valid_5_delay_37_12;
    io_A_Valid_5_delay_39_10 <= io_A_Valid_5_delay_38_11;
    io_A_Valid_5_delay_40_9 <= io_A_Valid_5_delay_39_10;
    io_A_Valid_5_delay_41_8 <= io_A_Valid_5_delay_40_9;
    io_A_Valid_5_delay_42_7 <= io_A_Valid_5_delay_41_8;
    io_A_Valid_5_delay_43_6 <= io_A_Valid_5_delay_42_7;
    io_A_Valid_5_delay_44_5 <= io_A_Valid_5_delay_43_6;
    io_A_Valid_5_delay_45_4 <= io_A_Valid_5_delay_44_5;
    io_A_Valid_5_delay_46_3 <= io_A_Valid_5_delay_45_4;
    io_A_Valid_5_delay_47_2 <= io_A_Valid_5_delay_46_3;
    io_A_Valid_5_delay_48_1 <= io_A_Valid_5_delay_47_2;
    io_A_Valid_5_delay_49 <= io_A_Valid_5_delay_48_1;
    io_B_Valid_49_delay_1_4 <= io_B_Valid_49;
    io_B_Valid_49_delay_2_3 <= io_B_Valid_49_delay_1_4;
    io_B_Valid_49_delay_3_2 <= io_B_Valid_49_delay_2_3;
    io_B_Valid_49_delay_4_1 <= io_B_Valid_49_delay_3_2;
    io_B_Valid_49_delay_5 <= io_B_Valid_49_delay_4_1;
    io_A_Valid_5_delay_1_49 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_48 <= io_A_Valid_5_delay_1_49;
    io_A_Valid_5_delay_3_47 <= io_A_Valid_5_delay_2_48;
    io_A_Valid_5_delay_4_46 <= io_A_Valid_5_delay_3_47;
    io_A_Valid_5_delay_5_45 <= io_A_Valid_5_delay_4_46;
    io_A_Valid_5_delay_6_44 <= io_A_Valid_5_delay_5_45;
    io_A_Valid_5_delay_7_43 <= io_A_Valid_5_delay_6_44;
    io_A_Valid_5_delay_8_42 <= io_A_Valid_5_delay_7_43;
    io_A_Valid_5_delay_9_41 <= io_A_Valid_5_delay_8_42;
    io_A_Valid_5_delay_10_40 <= io_A_Valid_5_delay_9_41;
    io_A_Valid_5_delay_11_39 <= io_A_Valid_5_delay_10_40;
    io_A_Valid_5_delay_12_38 <= io_A_Valid_5_delay_11_39;
    io_A_Valid_5_delay_13_37 <= io_A_Valid_5_delay_12_38;
    io_A_Valid_5_delay_14_36 <= io_A_Valid_5_delay_13_37;
    io_A_Valid_5_delay_15_35 <= io_A_Valid_5_delay_14_36;
    io_A_Valid_5_delay_16_34 <= io_A_Valid_5_delay_15_35;
    io_A_Valid_5_delay_17_33 <= io_A_Valid_5_delay_16_34;
    io_A_Valid_5_delay_18_32 <= io_A_Valid_5_delay_17_33;
    io_A_Valid_5_delay_19_31 <= io_A_Valid_5_delay_18_32;
    io_A_Valid_5_delay_20_30 <= io_A_Valid_5_delay_19_31;
    io_A_Valid_5_delay_21_29 <= io_A_Valid_5_delay_20_30;
    io_A_Valid_5_delay_22_28 <= io_A_Valid_5_delay_21_29;
    io_A_Valid_5_delay_23_27 <= io_A_Valid_5_delay_22_28;
    io_A_Valid_5_delay_24_26 <= io_A_Valid_5_delay_23_27;
    io_A_Valid_5_delay_25_25 <= io_A_Valid_5_delay_24_26;
    io_A_Valid_5_delay_26_24 <= io_A_Valid_5_delay_25_25;
    io_A_Valid_5_delay_27_23 <= io_A_Valid_5_delay_26_24;
    io_A_Valid_5_delay_28_22 <= io_A_Valid_5_delay_27_23;
    io_A_Valid_5_delay_29_21 <= io_A_Valid_5_delay_28_22;
    io_A_Valid_5_delay_30_20 <= io_A_Valid_5_delay_29_21;
    io_A_Valid_5_delay_31_19 <= io_A_Valid_5_delay_30_20;
    io_A_Valid_5_delay_32_18 <= io_A_Valid_5_delay_31_19;
    io_A_Valid_5_delay_33_17 <= io_A_Valid_5_delay_32_18;
    io_A_Valid_5_delay_34_16 <= io_A_Valid_5_delay_33_17;
    io_A_Valid_5_delay_35_15 <= io_A_Valid_5_delay_34_16;
    io_A_Valid_5_delay_36_14 <= io_A_Valid_5_delay_35_15;
    io_A_Valid_5_delay_37_13 <= io_A_Valid_5_delay_36_14;
    io_A_Valid_5_delay_38_12 <= io_A_Valid_5_delay_37_13;
    io_A_Valid_5_delay_39_11 <= io_A_Valid_5_delay_38_12;
    io_A_Valid_5_delay_40_10 <= io_A_Valid_5_delay_39_11;
    io_A_Valid_5_delay_41_9 <= io_A_Valid_5_delay_40_10;
    io_A_Valid_5_delay_42_8 <= io_A_Valid_5_delay_41_9;
    io_A_Valid_5_delay_43_7 <= io_A_Valid_5_delay_42_8;
    io_A_Valid_5_delay_44_6 <= io_A_Valid_5_delay_43_7;
    io_A_Valid_5_delay_45_5 <= io_A_Valid_5_delay_44_6;
    io_A_Valid_5_delay_46_4 <= io_A_Valid_5_delay_45_5;
    io_A_Valid_5_delay_47_3 <= io_A_Valid_5_delay_46_4;
    io_A_Valid_5_delay_48_2 <= io_A_Valid_5_delay_47_3;
    io_A_Valid_5_delay_49_1 <= io_A_Valid_5_delay_48_2;
    io_A_Valid_5_delay_50 <= io_A_Valid_5_delay_49_1;
    io_B_Valid_50_delay_1_4 <= io_B_Valid_50;
    io_B_Valid_50_delay_2_3 <= io_B_Valid_50_delay_1_4;
    io_B_Valid_50_delay_3_2 <= io_B_Valid_50_delay_2_3;
    io_B_Valid_50_delay_4_1 <= io_B_Valid_50_delay_3_2;
    io_B_Valid_50_delay_5 <= io_B_Valid_50_delay_4_1;
    io_A_Valid_5_delay_1_50 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_49 <= io_A_Valid_5_delay_1_50;
    io_A_Valid_5_delay_3_48 <= io_A_Valid_5_delay_2_49;
    io_A_Valid_5_delay_4_47 <= io_A_Valid_5_delay_3_48;
    io_A_Valid_5_delay_5_46 <= io_A_Valid_5_delay_4_47;
    io_A_Valid_5_delay_6_45 <= io_A_Valid_5_delay_5_46;
    io_A_Valid_5_delay_7_44 <= io_A_Valid_5_delay_6_45;
    io_A_Valid_5_delay_8_43 <= io_A_Valid_5_delay_7_44;
    io_A_Valid_5_delay_9_42 <= io_A_Valid_5_delay_8_43;
    io_A_Valid_5_delay_10_41 <= io_A_Valid_5_delay_9_42;
    io_A_Valid_5_delay_11_40 <= io_A_Valid_5_delay_10_41;
    io_A_Valid_5_delay_12_39 <= io_A_Valid_5_delay_11_40;
    io_A_Valid_5_delay_13_38 <= io_A_Valid_5_delay_12_39;
    io_A_Valid_5_delay_14_37 <= io_A_Valid_5_delay_13_38;
    io_A_Valid_5_delay_15_36 <= io_A_Valid_5_delay_14_37;
    io_A_Valid_5_delay_16_35 <= io_A_Valid_5_delay_15_36;
    io_A_Valid_5_delay_17_34 <= io_A_Valid_5_delay_16_35;
    io_A_Valid_5_delay_18_33 <= io_A_Valid_5_delay_17_34;
    io_A_Valid_5_delay_19_32 <= io_A_Valid_5_delay_18_33;
    io_A_Valid_5_delay_20_31 <= io_A_Valid_5_delay_19_32;
    io_A_Valid_5_delay_21_30 <= io_A_Valid_5_delay_20_31;
    io_A_Valid_5_delay_22_29 <= io_A_Valid_5_delay_21_30;
    io_A_Valid_5_delay_23_28 <= io_A_Valid_5_delay_22_29;
    io_A_Valid_5_delay_24_27 <= io_A_Valid_5_delay_23_28;
    io_A_Valid_5_delay_25_26 <= io_A_Valid_5_delay_24_27;
    io_A_Valid_5_delay_26_25 <= io_A_Valid_5_delay_25_26;
    io_A_Valid_5_delay_27_24 <= io_A_Valid_5_delay_26_25;
    io_A_Valid_5_delay_28_23 <= io_A_Valid_5_delay_27_24;
    io_A_Valid_5_delay_29_22 <= io_A_Valid_5_delay_28_23;
    io_A_Valid_5_delay_30_21 <= io_A_Valid_5_delay_29_22;
    io_A_Valid_5_delay_31_20 <= io_A_Valid_5_delay_30_21;
    io_A_Valid_5_delay_32_19 <= io_A_Valid_5_delay_31_20;
    io_A_Valid_5_delay_33_18 <= io_A_Valid_5_delay_32_19;
    io_A_Valid_5_delay_34_17 <= io_A_Valid_5_delay_33_18;
    io_A_Valid_5_delay_35_16 <= io_A_Valid_5_delay_34_17;
    io_A_Valid_5_delay_36_15 <= io_A_Valid_5_delay_35_16;
    io_A_Valid_5_delay_37_14 <= io_A_Valid_5_delay_36_15;
    io_A_Valid_5_delay_38_13 <= io_A_Valid_5_delay_37_14;
    io_A_Valid_5_delay_39_12 <= io_A_Valid_5_delay_38_13;
    io_A_Valid_5_delay_40_11 <= io_A_Valid_5_delay_39_12;
    io_A_Valid_5_delay_41_10 <= io_A_Valid_5_delay_40_11;
    io_A_Valid_5_delay_42_9 <= io_A_Valid_5_delay_41_10;
    io_A_Valid_5_delay_43_8 <= io_A_Valid_5_delay_42_9;
    io_A_Valid_5_delay_44_7 <= io_A_Valid_5_delay_43_8;
    io_A_Valid_5_delay_45_6 <= io_A_Valid_5_delay_44_7;
    io_A_Valid_5_delay_46_5 <= io_A_Valid_5_delay_45_6;
    io_A_Valid_5_delay_47_4 <= io_A_Valid_5_delay_46_5;
    io_A_Valid_5_delay_48_3 <= io_A_Valid_5_delay_47_4;
    io_A_Valid_5_delay_49_2 <= io_A_Valid_5_delay_48_3;
    io_A_Valid_5_delay_50_1 <= io_A_Valid_5_delay_49_2;
    io_A_Valid_5_delay_51 <= io_A_Valid_5_delay_50_1;
    io_B_Valid_51_delay_1_4 <= io_B_Valid_51;
    io_B_Valid_51_delay_2_3 <= io_B_Valid_51_delay_1_4;
    io_B_Valid_51_delay_3_2 <= io_B_Valid_51_delay_2_3;
    io_B_Valid_51_delay_4_1 <= io_B_Valid_51_delay_3_2;
    io_B_Valid_51_delay_5 <= io_B_Valid_51_delay_4_1;
    io_A_Valid_5_delay_1_51 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_50 <= io_A_Valid_5_delay_1_51;
    io_A_Valid_5_delay_3_49 <= io_A_Valid_5_delay_2_50;
    io_A_Valid_5_delay_4_48 <= io_A_Valid_5_delay_3_49;
    io_A_Valid_5_delay_5_47 <= io_A_Valid_5_delay_4_48;
    io_A_Valid_5_delay_6_46 <= io_A_Valid_5_delay_5_47;
    io_A_Valid_5_delay_7_45 <= io_A_Valid_5_delay_6_46;
    io_A_Valid_5_delay_8_44 <= io_A_Valid_5_delay_7_45;
    io_A_Valid_5_delay_9_43 <= io_A_Valid_5_delay_8_44;
    io_A_Valid_5_delay_10_42 <= io_A_Valid_5_delay_9_43;
    io_A_Valid_5_delay_11_41 <= io_A_Valid_5_delay_10_42;
    io_A_Valid_5_delay_12_40 <= io_A_Valid_5_delay_11_41;
    io_A_Valid_5_delay_13_39 <= io_A_Valid_5_delay_12_40;
    io_A_Valid_5_delay_14_38 <= io_A_Valid_5_delay_13_39;
    io_A_Valid_5_delay_15_37 <= io_A_Valid_5_delay_14_38;
    io_A_Valid_5_delay_16_36 <= io_A_Valid_5_delay_15_37;
    io_A_Valid_5_delay_17_35 <= io_A_Valid_5_delay_16_36;
    io_A_Valid_5_delay_18_34 <= io_A_Valid_5_delay_17_35;
    io_A_Valid_5_delay_19_33 <= io_A_Valid_5_delay_18_34;
    io_A_Valid_5_delay_20_32 <= io_A_Valid_5_delay_19_33;
    io_A_Valid_5_delay_21_31 <= io_A_Valid_5_delay_20_32;
    io_A_Valid_5_delay_22_30 <= io_A_Valid_5_delay_21_31;
    io_A_Valid_5_delay_23_29 <= io_A_Valid_5_delay_22_30;
    io_A_Valid_5_delay_24_28 <= io_A_Valid_5_delay_23_29;
    io_A_Valid_5_delay_25_27 <= io_A_Valid_5_delay_24_28;
    io_A_Valid_5_delay_26_26 <= io_A_Valid_5_delay_25_27;
    io_A_Valid_5_delay_27_25 <= io_A_Valid_5_delay_26_26;
    io_A_Valid_5_delay_28_24 <= io_A_Valid_5_delay_27_25;
    io_A_Valid_5_delay_29_23 <= io_A_Valid_5_delay_28_24;
    io_A_Valid_5_delay_30_22 <= io_A_Valid_5_delay_29_23;
    io_A_Valid_5_delay_31_21 <= io_A_Valid_5_delay_30_22;
    io_A_Valid_5_delay_32_20 <= io_A_Valid_5_delay_31_21;
    io_A_Valid_5_delay_33_19 <= io_A_Valid_5_delay_32_20;
    io_A_Valid_5_delay_34_18 <= io_A_Valid_5_delay_33_19;
    io_A_Valid_5_delay_35_17 <= io_A_Valid_5_delay_34_18;
    io_A_Valid_5_delay_36_16 <= io_A_Valid_5_delay_35_17;
    io_A_Valid_5_delay_37_15 <= io_A_Valid_5_delay_36_16;
    io_A_Valid_5_delay_38_14 <= io_A_Valid_5_delay_37_15;
    io_A_Valid_5_delay_39_13 <= io_A_Valid_5_delay_38_14;
    io_A_Valid_5_delay_40_12 <= io_A_Valid_5_delay_39_13;
    io_A_Valid_5_delay_41_11 <= io_A_Valid_5_delay_40_12;
    io_A_Valid_5_delay_42_10 <= io_A_Valid_5_delay_41_11;
    io_A_Valid_5_delay_43_9 <= io_A_Valid_5_delay_42_10;
    io_A_Valid_5_delay_44_8 <= io_A_Valid_5_delay_43_9;
    io_A_Valid_5_delay_45_7 <= io_A_Valid_5_delay_44_8;
    io_A_Valid_5_delay_46_6 <= io_A_Valid_5_delay_45_7;
    io_A_Valid_5_delay_47_5 <= io_A_Valid_5_delay_46_6;
    io_A_Valid_5_delay_48_4 <= io_A_Valid_5_delay_47_5;
    io_A_Valid_5_delay_49_3 <= io_A_Valid_5_delay_48_4;
    io_A_Valid_5_delay_50_2 <= io_A_Valid_5_delay_49_3;
    io_A_Valid_5_delay_51_1 <= io_A_Valid_5_delay_50_2;
    io_A_Valid_5_delay_52 <= io_A_Valid_5_delay_51_1;
    io_B_Valid_52_delay_1_4 <= io_B_Valid_52;
    io_B_Valid_52_delay_2_3 <= io_B_Valid_52_delay_1_4;
    io_B_Valid_52_delay_3_2 <= io_B_Valid_52_delay_2_3;
    io_B_Valid_52_delay_4_1 <= io_B_Valid_52_delay_3_2;
    io_B_Valid_52_delay_5 <= io_B_Valid_52_delay_4_1;
    io_A_Valid_5_delay_1_52 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_51 <= io_A_Valid_5_delay_1_52;
    io_A_Valid_5_delay_3_50 <= io_A_Valid_5_delay_2_51;
    io_A_Valid_5_delay_4_49 <= io_A_Valid_5_delay_3_50;
    io_A_Valid_5_delay_5_48 <= io_A_Valid_5_delay_4_49;
    io_A_Valid_5_delay_6_47 <= io_A_Valid_5_delay_5_48;
    io_A_Valid_5_delay_7_46 <= io_A_Valid_5_delay_6_47;
    io_A_Valid_5_delay_8_45 <= io_A_Valid_5_delay_7_46;
    io_A_Valid_5_delay_9_44 <= io_A_Valid_5_delay_8_45;
    io_A_Valid_5_delay_10_43 <= io_A_Valid_5_delay_9_44;
    io_A_Valid_5_delay_11_42 <= io_A_Valid_5_delay_10_43;
    io_A_Valid_5_delay_12_41 <= io_A_Valid_5_delay_11_42;
    io_A_Valid_5_delay_13_40 <= io_A_Valid_5_delay_12_41;
    io_A_Valid_5_delay_14_39 <= io_A_Valid_5_delay_13_40;
    io_A_Valid_5_delay_15_38 <= io_A_Valid_5_delay_14_39;
    io_A_Valid_5_delay_16_37 <= io_A_Valid_5_delay_15_38;
    io_A_Valid_5_delay_17_36 <= io_A_Valid_5_delay_16_37;
    io_A_Valid_5_delay_18_35 <= io_A_Valid_5_delay_17_36;
    io_A_Valid_5_delay_19_34 <= io_A_Valid_5_delay_18_35;
    io_A_Valid_5_delay_20_33 <= io_A_Valid_5_delay_19_34;
    io_A_Valid_5_delay_21_32 <= io_A_Valid_5_delay_20_33;
    io_A_Valid_5_delay_22_31 <= io_A_Valid_5_delay_21_32;
    io_A_Valid_5_delay_23_30 <= io_A_Valid_5_delay_22_31;
    io_A_Valid_5_delay_24_29 <= io_A_Valid_5_delay_23_30;
    io_A_Valid_5_delay_25_28 <= io_A_Valid_5_delay_24_29;
    io_A_Valid_5_delay_26_27 <= io_A_Valid_5_delay_25_28;
    io_A_Valid_5_delay_27_26 <= io_A_Valid_5_delay_26_27;
    io_A_Valid_5_delay_28_25 <= io_A_Valid_5_delay_27_26;
    io_A_Valid_5_delay_29_24 <= io_A_Valid_5_delay_28_25;
    io_A_Valid_5_delay_30_23 <= io_A_Valid_5_delay_29_24;
    io_A_Valid_5_delay_31_22 <= io_A_Valid_5_delay_30_23;
    io_A_Valid_5_delay_32_21 <= io_A_Valid_5_delay_31_22;
    io_A_Valid_5_delay_33_20 <= io_A_Valid_5_delay_32_21;
    io_A_Valid_5_delay_34_19 <= io_A_Valid_5_delay_33_20;
    io_A_Valid_5_delay_35_18 <= io_A_Valid_5_delay_34_19;
    io_A_Valid_5_delay_36_17 <= io_A_Valid_5_delay_35_18;
    io_A_Valid_5_delay_37_16 <= io_A_Valid_5_delay_36_17;
    io_A_Valid_5_delay_38_15 <= io_A_Valid_5_delay_37_16;
    io_A_Valid_5_delay_39_14 <= io_A_Valid_5_delay_38_15;
    io_A_Valid_5_delay_40_13 <= io_A_Valid_5_delay_39_14;
    io_A_Valid_5_delay_41_12 <= io_A_Valid_5_delay_40_13;
    io_A_Valid_5_delay_42_11 <= io_A_Valid_5_delay_41_12;
    io_A_Valid_5_delay_43_10 <= io_A_Valid_5_delay_42_11;
    io_A_Valid_5_delay_44_9 <= io_A_Valid_5_delay_43_10;
    io_A_Valid_5_delay_45_8 <= io_A_Valid_5_delay_44_9;
    io_A_Valid_5_delay_46_7 <= io_A_Valid_5_delay_45_8;
    io_A_Valid_5_delay_47_6 <= io_A_Valid_5_delay_46_7;
    io_A_Valid_5_delay_48_5 <= io_A_Valid_5_delay_47_6;
    io_A_Valid_5_delay_49_4 <= io_A_Valid_5_delay_48_5;
    io_A_Valid_5_delay_50_3 <= io_A_Valid_5_delay_49_4;
    io_A_Valid_5_delay_51_2 <= io_A_Valid_5_delay_50_3;
    io_A_Valid_5_delay_52_1 <= io_A_Valid_5_delay_51_2;
    io_A_Valid_5_delay_53 <= io_A_Valid_5_delay_52_1;
    io_B_Valid_53_delay_1_4 <= io_B_Valid_53;
    io_B_Valid_53_delay_2_3 <= io_B_Valid_53_delay_1_4;
    io_B_Valid_53_delay_3_2 <= io_B_Valid_53_delay_2_3;
    io_B_Valid_53_delay_4_1 <= io_B_Valid_53_delay_3_2;
    io_B_Valid_53_delay_5 <= io_B_Valid_53_delay_4_1;
    io_A_Valid_5_delay_1_53 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_52 <= io_A_Valid_5_delay_1_53;
    io_A_Valid_5_delay_3_51 <= io_A_Valid_5_delay_2_52;
    io_A_Valid_5_delay_4_50 <= io_A_Valid_5_delay_3_51;
    io_A_Valid_5_delay_5_49 <= io_A_Valid_5_delay_4_50;
    io_A_Valid_5_delay_6_48 <= io_A_Valid_5_delay_5_49;
    io_A_Valid_5_delay_7_47 <= io_A_Valid_5_delay_6_48;
    io_A_Valid_5_delay_8_46 <= io_A_Valid_5_delay_7_47;
    io_A_Valid_5_delay_9_45 <= io_A_Valid_5_delay_8_46;
    io_A_Valid_5_delay_10_44 <= io_A_Valid_5_delay_9_45;
    io_A_Valid_5_delay_11_43 <= io_A_Valid_5_delay_10_44;
    io_A_Valid_5_delay_12_42 <= io_A_Valid_5_delay_11_43;
    io_A_Valid_5_delay_13_41 <= io_A_Valid_5_delay_12_42;
    io_A_Valid_5_delay_14_40 <= io_A_Valid_5_delay_13_41;
    io_A_Valid_5_delay_15_39 <= io_A_Valid_5_delay_14_40;
    io_A_Valid_5_delay_16_38 <= io_A_Valid_5_delay_15_39;
    io_A_Valid_5_delay_17_37 <= io_A_Valid_5_delay_16_38;
    io_A_Valid_5_delay_18_36 <= io_A_Valid_5_delay_17_37;
    io_A_Valid_5_delay_19_35 <= io_A_Valid_5_delay_18_36;
    io_A_Valid_5_delay_20_34 <= io_A_Valid_5_delay_19_35;
    io_A_Valid_5_delay_21_33 <= io_A_Valid_5_delay_20_34;
    io_A_Valid_5_delay_22_32 <= io_A_Valid_5_delay_21_33;
    io_A_Valid_5_delay_23_31 <= io_A_Valid_5_delay_22_32;
    io_A_Valid_5_delay_24_30 <= io_A_Valid_5_delay_23_31;
    io_A_Valid_5_delay_25_29 <= io_A_Valid_5_delay_24_30;
    io_A_Valid_5_delay_26_28 <= io_A_Valid_5_delay_25_29;
    io_A_Valid_5_delay_27_27 <= io_A_Valid_5_delay_26_28;
    io_A_Valid_5_delay_28_26 <= io_A_Valid_5_delay_27_27;
    io_A_Valid_5_delay_29_25 <= io_A_Valid_5_delay_28_26;
    io_A_Valid_5_delay_30_24 <= io_A_Valid_5_delay_29_25;
    io_A_Valid_5_delay_31_23 <= io_A_Valid_5_delay_30_24;
    io_A_Valid_5_delay_32_22 <= io_A_Valid_5_delay_31_23;
    io_A_Valid_5_delay_33_21 <= io_A_Valid_5_delay_32_22;
    io_A_Valid_5_delay_34_20 <= io_A_Valid_5_delay_33_21;
    io_A_Valid_5_delay_35_19 <= io_A_Valid_5_delay_34_20;
    io_A_Valid_5_delay_36_18 <= io_A_Valid_5_delay_35_19;
    io_A_Valid_5_delay_37_17 <= io_A_Valid_5_delay_36_18;
    io_A_Valid_5_delay_38_16 <= io_A_Valid_5_delay_37_17;
    io_A_Valid_5_delay_39_15 <= io_A_Valid_5_delay_38_16;
    io_A_Valid_5_delay_40_14 <= io_A_Valid_5_delay_39_15;
    io_A_Valid_5_delay_41_13 <= io_A_Valid_5_delay_40_14;
    io_A_Valid_5_delay_42_12 <= io_A_Valid_5_delay_41_13;
    io_A_Valid_5_delay_43_11 <= io_A_Valid_5_delay_42_12;
    io_A_Valid_5_delay_44_10 <= io_A_Valid_5_delay_43_11;
    io_A_Valid_5_delay_45_9 <= io_A_Valid_5_delay_44_10;
    io_A_Valid_5_delay_46_8 <= io_A_Valid_5_delay_45_9;
    io_A_Valid_5_delay_47_7 <= io_A_Valid_5_delay_46_8;
    io_A_Valid_5_delay_48_6 <= io_A_Valid_5_delay_47_7;
    io_A_Valid_5_delay_49_5 <= io_A_Valid_5_delay_48_6;
    io_A_Valid_5_delay_50_4 <= io_A_Valid_5_delay_49_5;
    io_A_Valid_5_delay_51_3 <= io_A_Valid_5_delay_50_4;
    io_A_Valid_5_delay_52_2 <= io_A_Valid_5_delay_51_3;
    io_A_Valid_5_delay_53_1 <= io_A_Valid_5_delay_52_2;
    io_A_Valid_5_delay_54 <= io_A_Valid_5_delay_53_1;
    io_B_Valid_54_delay_1_4 <= io_B_Valid_54;
    io_B_Valid_54_delay_2_3 <= io_B_Valid_54_delay_1_4;
    io_B_Valid_54_delay_3_2 <= io_B_Valid_54_delay_2_3;
    io_B_Valid_54_delay_4_1 <= io_B_Valid_54_delay_3_2;
    io_B_Valid_54_delay_5 <= io_B_Valid_54_delay_4_1;
    io_A_Valid_5_delay_1_54 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_53 <= io_A_Valid_5_delay_1_54;
    io_A_Valid_5_delay_3_52 <= io_A_Valid_5_delay_2_53;
    io_A_Valid_5_delay_4_51 <= io_A_Valid_5_delay_3_52;
    io_A_Valid_5_delay_5_50 <= io_A_Valid_5_delay_4_51;
    io_A_Valid_5_delay_6_49 <= io_A_Valid_5_delay_5_50;
    io_A_Valid_5_delay_7_48 <= io_A_Valid_5_delay_6_49;
    io_A_Valid_5_delay_8_47 <= io_A_Valid_5_delay_7_48;
    io_A_Valid_5_delay_9_46 <= io_A_Valid_5_delay_8_47;
    io_A_Valid_5_delay_10_45 <= io_A_Valid_5_delay_9_46;
    io_A_Valid_5_delay_11_44 <= io_A_Valid_5_delay_10_45;
    io_A_Valid_5_delay_12_43 <= io_A_Valid_5_delay_11_44;
    io_A_Valid_5_delay_13_42 <= io_A_Valid_5_delay_12_43;
    io_A_Valid_5_delay_14_41 <= io_A_Valid_5_delay_13_42;
    io_A_Valid_5_delay_15_40 <= io_A_Valid_5_delay_14_41;
    io_A_Valid_5_delay_16_39 <= io_A_Valid_5_delay_15_40;
    io_A_Valid_5_delay_17_38 <= io_A_Valid_5_delay_16_39;
    io_A_Valid_5_delay_18_37 <= io_A_Valid_5_delay_17_38;
    io_A_Valid_5_delay_19_36 <= io_A_Valid_5_delay_18_37;
    io_A_Valid_5_delay_20_35 <= io_A_Valid_5_delay_19_36;
    io_A_Valid_5_delay_21_34 <= io_A_Valid_5_delay_20_35;
    io_A_Valid_5_delay_22_33 <= io_A_Valid_5_delay_21_34;
    io_A_Valid_5_delay_23_32 <= io_A_Valid_5_delay_22_33;
    io_A_Valid_5_delay_24_31 <= io_A_Valid_5_delay_23_32;
    io_A_Valid_5_delay_25_30 <= io_A_Valid_5_delay_24_31;
    io_A_Valid_5_delay_26_29 <= io_A_Valid_5_delay_25_30;
    io_A_Valid_5_delay_27_28 <= io_A_Valid_5_delay_26_29;
    io_A_Valid_5_delay_28_27 <= io_A_Valid_5_delay_27_28;
    io_A_Valid_5_delay_29_26 <= io_A_Valid_5_delay_28_27;
    io_A_Valid_5_delay_30_25 <= io_A_Valid_5_delay_29_26;
    io_A_Valid_5_delay_31_24 <= io_A_Valid_5_delay_30_25;
    io_A_Valid_5_delay_32_23 <= io_A_Valid_5_delay_31_24;
    io_A_Valid_5_delay_33_22 <= io_A_Valid_5_delay_32_23;
    io_A_Valid_5_delay_34_21 <= io_A_Valid_5_delay_33_22;
    io_A_Valid_5_delay_35_20 <= io_A_Valid_5_delay_34_21;
    io_A_Valid_5_delay_36_19 <= io_A_Valid_5_delay_35_20;
    io_A_Valid_5_delay_37_18 <= io_A_Valid_5_delay_36_19;
    io_A_Valid_5_delay_38_17 <= io_A_Valid_5_delay_37_18;
    io_A_Valid_5_delay_39_16 <= io_A_Valid_5_delay_38_17;
    io_A_Valid_5_delay_40_15 <= io_A_Valid_5_delay_39_16;
    io_A_Valid_5_delay_41_14 <= io_A_Valid_5_delay_40_15;
    io_A_Valid_5_delay_42_13 <= io_A_Valid_5_delay_41_14;
    io_A_Valid_5_delay_43_12 <= io_A_Valid_5_delay_42_13;
    io_A_Valid_5_delay_44_11 <= io_A_Valid_5_delay_43_12;
    io_A_Valid_5_delay_45_10 <= io_A_Valid_5_delay_44_11;
    io_A_Valid_5_delay_46_9 <= io_A_Valid_5_delay_45_10;
    io_A_Valid_5_delay_47_8 <= io_A_Valid_5_delay_46_9;
    io_A_Valid_5_delay_48_7 <= io_A_Valid_5_delay_47_8;
    io_A_Valid_5_delay_49_6 <= io_A_Valid_5_delay_48_7;
    io_A_Valid_5_delay_50_5 <= io_A_Valid_5_delay_49_6;
    io_A_Valid_5_delay_51_4 <= io_A_Valid_5_delay_50_5;
    io_A_Valid_5_delay_52_3 <= io_A_Valid_5_delay_51_4;
    io_A_Valid_5_delay_53_2 <= io_A_Valid_5_delay_52_3;
    io_A_Valid_5_delay_54_1 <= io_A_Valid_5_delay_53_2;
    io_A_Valid_5_delay_55 <= io_A_Valid_5_delay_54_1;
    io_B_Valid_55_delay_1_4 <= io_B_Valid_55;
    io_B_Valid_55_delay_2_3 <= io_B_Valid_55_delay_1_4;
    io_B_Valid_55_delay_3_2 <= io_B_Valid_55_delay_2_3;
    io_B_Valid_55_delay_4_1 <= io_B_Valid_55_delay_3_2;
    io_B_Valid_55_delay_5 <= io_B_Valid_55_delay_4_1;
    io_A_Valid_5_delay_1_55 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_54 <= io_A_Valid_5_delay_1_55;
    io_A_Valid_5_delay_3_53 <= io_A_Valid_5_delay_2_54;
    io_A_Valid_5_delay_4_52 <= io_A_Valid_5_delay_3_53;
    io_A_Valid_5_delay_5_51 <= io_A_Valid_5_delay_4_52;
    io_A_Valid_5_delay_6_50 <= io_A_Valid_5_delay_5_51;
    io_A_Valid_5_delay_7_49 <= io_A_Valid_5_delay_6_50;
    io_A_Valid_5_delay_8_48 <= io_A_Valid_5_delay_7_49;
    io_A_Valid_5_delay_9_47 <= io_A_Valid_5_delay_8_48;
    io_A_Valid_5_delay_10_46 <= io_A_Valid_5_delay_9_47;
    io_A_Valid_5_delay_11_45 <= io_A_Valid_5_delay_10_46;
    io_A_Valid_5_delay_12_44 <= io_A_Valid_5_delay_11_45;
    io_A_Valid_5_delay_13_43 <= io_A_Valid_5_delay_12_44;
    io_A_Valid_5_delay_14_42 <= io_A_Valid_5_delay_13_43;
    io_A_Valid_5_delay_15_41 <= io_A_Valid_5_delay_14_42;
    io_A_Valid_5_delay_16_40 <= io_A_Valid_5_delay_15_41;
    io_A_Valid_5_delay_17_39 <= io_A_Valid_5_delay_16_40;
    io_A_Valid_5_delay_18_38 <= io_A_Valid_5_delay_17_39;
    io_A_Valid_5_delay_19_37 <= io_A_Valid_5_delay_18_38;
    io_A_Valid_5_delay_20_36 <= io_A_Valid_5_delay_19_37;
    io_A_Valid_5_delay_21_35 <= io_A_Valid_5_delay_20_36;
    io_A_Valid_5_delay_22_34 <= io_A_Valid_5_delay_21_35;
    io_A_Valid_5_delay_23_33 <= io_A_Valid_5_delay_22_34;
    io_A_Valid_5_delay_24_32 <= io_A_Valid_5_delay_23_33;
    io_A_Valid_5_delay_25_31 <= io_A_Valid_5_delay_24_32;
    io_A_Valid_5_delay_26_30 <= io_A_Valid_5_delay_25_31;
    io_A_Valid_5_delay_27_29 <= io_A_Valid_5_delay_26_30;
    io_A_Valid_5_delay_28_28 <= io_A_Valid_5_delay_27_29;
    io_A_Valid_5_delay_29_27 <= io_A_Valid_5_delay_28_28;
    io_A_Valid_5_delay_30_26 <= io_A_Valid_5_delay_29_27;
    io_A_Valid_5_delay_31_25 <= io_A_Valid_5_delay_30_26;
    io_A_Valid_5_delay_32_24 <= io_A_Valid_5_delay_31_25;
    io_A_Valid_5_delay_33_23 <= io_A_Valid_5_delay_32_24;
    io_A_Valid_5_delay_34_22 <= io_A_Valid_5_delay_33_23;
    io_A_Valid_5_delay_35_21 <= io_A_Valid_5_delay_34_22;
    io_A_Valid_5_delay_36_20 <= io_A_Valid_5_delay_35_21;
    io_A_Valid_5_delay_37_19 <= io_A_Valid_5_delay_36_20;
    io_A_Valid_5_delay_38_18 <= io_A_Valid_5_delay_37_19;
    io_A_Valid_5_delay_39_17 <= io_A_Valid_5_delay_38_18;
    io_A_Valid_5_delay_40_16 <= io_A_Valid_5_delay_39_17;
    io_A_Valid_5_delay_41_15 <= io_A_Valid_5_delay_40_16;
    io_A_Valid_5_delay_42_14 <= io_A_Valid_5_delay_41_15;
    io_A_Valid_5_delay_43_13 <= io_A_Valid_5_delay_42_14;
    io_A_Valid_5_delay_44_12 <= io_A_Valid_5_delay_43_13;
    io_A_Valid_5_delay_45_11 <= io_A_Valid_5_delay_44_12;
    io_A_Valid_5_delay_46_10 <= io_A_Valid_5_delay_45_11;
    io_A_Valid_5_delay_47_9 <= io_A_Valid_5_delay_46_10;
    io_A_Valid_5_delay_48_8 <= io_A_Valid_5_delay_47_9;
    io_A_Valid_5_delay_49_7 <= io_A_Valid_5_delay_48_8;
    io_A_Valid_5_delay_50_6 <= io_A_Valid_5_delay_49_7;
    io_A_Valid_5_delay_51_5 <= io_A_Valid_5_delay_50_6;
    io_A_Valid_5_delay_52_4 <= io_A_Valid_5_delay_51_5;
    io_A_Valid_5_delay_53_3 <= io_A_Valid_5_delay_52_4;
    io_A_Valid_5_delay_54_2 <= io_A_Valid_5_delay_53_3;
    io_A_Valid_5_delay_55_1 <= io_A_Valid_5_delay_54_2;
    io_A_Valid_5_delay_56 <= io_A_Valid_5_delay_55_1;
    io_B_Valid_56_delay_1_4 <= io_B_Valid_56;
    io_B_Valid_56_delay_2_3 <= io_B_Valid_56_delay_1_4;
    io_B_Valid_56_delay_3_2 <= io_B_Valid_56_delay_2_3;
    io_B_Valid_56_delay_4_1 <= io_B_Valid_56_delay_3_2;
    io_B_Valid_56_delay_5 <= io_B_Valid_56_delay_4_1;
    io_A_Valid_5_delay_1_56 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_55 <= io_A_Valid_5_delay_1_56;
    io_A_Valid_5_delay_3_54 <= io_A_Valid_5_delay_2_55;
    io_A_Valid_5_delay_4_53 <= io_A_Valid_5_delay_3_54;
    io_A_Valid_5_delay_5_52 <= io_A_Valid_5_delay_4_53;
    io_A_Valid_5_delay_6_51 <= io_A_Valid_5_delay_5_52;
    io_A_Valid_5_delay_7_50 <= io_A_Valid_5_delay_6_51;
    io_A_Valid_5_delay_8_49 <= io_A_Valid_5_delay_7_50;
    io_A_Valid_5_delay_9_48 <= io_A_Valid_5_delay_8_49;
    io_A_Valid_5_delay_10_47 <= io_A_Valid_5_delay_9_48;
    io_A_Valid_5_delay_11_46 <= io_A_Valid_5_delay_10_47;
    io_A_Valid_5_delay_12_45 <= io_A_Valid_5_delay_11_46;
    io_A_Valid_5_delay_13_44 <= io_A_Valid_5_delay_12_45;
    io_A_Valid_5_delay_14_43 <= io_A_Valid_5_delay_13_44;
    io_A_Valid_5_delay_15_42 <= io_A_Valid_5_delay_14_43;
    io_A_Valid_5_delay_16_41 <= io_A_Valid_5_delay_15_42;
    io_A_Valid_5_delay_17_40 <= io_A_Valid_5_delay_16_41;
    io_A_Valid_5_delay_18_39 <= io_A_Valid_5_delay_17_40;
    io_A_Valid_5_delay_19_38 <= io_A_Valid_5_delay_18_39;
    io_A_Valid_5_delay_20_37 <= io_A_Valid_5_delay_19_38;
    io_A_Valid_5_delay_21_36 <= io_A_Valid_5_delay_20_37;
    io_A_Valid_5_delay_22_35 <= io_A_Valid_5_delay_21_36;
    io_A_Valid_5_delay_23_34 <= io_A_Valid_5_delay_22_35;
    io_A_Valid_5_delay_24_33 <= io_A_Valid_5_delay_23_34;
    io_A_Valid_5_delay_25_32 <= io_A_Valid_5_delay_24_33;
    io_A_Valid_5_delay_26_31 <= io_A_Valid_5_delay_25_32;
    io_A_Valid_5_delay_27_30 <= io_A_Valid_5_delay_26_31;
    io_A_Valid_5_delay_28_29 <= io_A_Valid_5_delay_27_30;
    io_A_Valid_5_delay_29_28 <= io_A_Valid_5_delay_28_29;
    io_A_Valid_5_delay_30_27 <= io_A_Valid_5_delay_29_28;
    io_A_Valid_5_delay_31_26 <= io_A_Valid_5_delay_30_27;
    io_A_Valid_5_delay_32_25 <= io_A_Valid_5_delay_31_26;
    io_A_Valid_5_delay_33_24 <= io_A_Valid_5_delay_32_25;
    io_A_Valid_5_delay_34_23 <= io_A_Valid_5_delay_33_24;
    io_A_Valid_5_delay_35_22 <= io_A_Valid_5_delay_34_23;
    io_A_Valid_5_delay_36_21 <= io_A_Valid_5_delay_35_22;
    io_A_Valid_5_delay_37_20 <= io_A_Valid_5_delay_36_21;
    io_A_Valid_5_delay_38_19 <= io_A_Valid_5_delay_37_20;
    io_A_Valid_5_delay_39_18 <= io_A_Valid_5_delay_38_19;
    io_A_Valid_5_delay_40_17 <= io_A_Valid_5_delay_39_18;
    io_A_Valid_5_delay_41_16 <= io_A_Valid_5_delay_40_17;
    io_A_Valid_5_delay_42_15 <= io_A_Valid_5_delay_41_16;
    io_A_Valid_5_delay_43_14 <= io_A_Valid_5_delay_42_15;
    io_A_Valid_5_delay_44_13 <= io_A_Valid_5_delay_43_14;
    io_A_Valid_5_delay_45_12 <= io_A_Valid_5_delay_44_13;
    io_A_Valid_5_delay_46_11 <= io_A_Valid_5_delay_45_12;
    io_A_Valid_5_delay_47_10 <= io_A_Valid_5_delay_46_11;
    io_A_Valid_5_delay_48_9 <= io_A_Valid_5_delay_47_10;
    io_A_Valid_5_delay_49_8 <= io_A_Valid_5_delay_48_9;
    io_A_Valid_5_delay_50_7 <= io_A_Valid_5_delay_49_8;
    io_A_Valid_5_delay_51_6 <= io_A_Valid_5_delay_50_7;
    io_A_Valid_5_delay_52_5 <= io_A_Valid_5_delay_51_6;
    io_A_Valid_5_delay_53_4 <= io_A_Valid_5_delay_52_5;
    io_A_Valid_5_delay_54_3 <= io_A_Valid_5_delay_53_4;
    io_A_Valid_5_delay_55_2 <= io_A_Valid_5_delay_54_3;
    io_A_Valid_5_delay_56_1 <= io_A_Valid_5_delay_55_2;
    io_A_Valid_5_delay_57 <= io_A_Valid_5_delay_56_1;
    io_B_Valid_57_delay_1_4 <= io_B_Valid_57;
    io_B_Valid_57_delay_2_3 <= io_B_Valid_57_delay_1_4;
    io_B_Valid_57_delay_3_2 <= io_B_Valid_57_delay_2_3;
    io_B_Valid_57_delay_4_1 <= io_B_Valid_57_delay_3_2;
    io_B_Valid_57_delay_5 <= io_B_Valid_57_delay_4_1;
    io_A_Valid_5_delay_1_57 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_56 <= io_A_Valid_5_delay_1_57;
    io_A_Valid_5_delay_3_55 <= io_A_Valid_5_delay_2_56;
    io_A_Valid_5_delay_4_54 <= io_A_Valid_5_delay_3_55;
    io_A_Valid_5_delay_5_53 <= io_A_Valid_5_delay_4_54;
    io_A_Valid_5_delay_6_52 <= io_A_Valid_5_delay_5_53;
    io_A_Valid_5_delay_7_51 <= io_A_Valid_5_delay_6_52;
    io_A_Valid_5_delay_8_50 <= io_A_Valid_5_delay_7_51;
    io_A_Valid_5_delay_9_49 <= io_A_Valid_5_delay_8_50;
    io_A_Valid_5_delay_10_48 <= io_A_Valid_5_delay_9_49;
    io_A_Valid_5_delay_11_47 <= io_A_Valid_5_delay_10_48;
    io_A_Valid_5_delay_12_46 <= io_A_Valid_5_delay_11_47;
    io_A_Valid_5_delay_13_45 <= io_A_Valid_5_delay_12_46;
    io_A_Valid_5_delay_14_44 <= io_A_Valid_5_delay_13_45;
    io_A_Valid_5_delay_15_43 <= io_A_Valid_5_delay_14_44;
    io_A_Valid_5_delay_16_42 <= io_A_Valid_5_delay_15_43;
    io_A_Valid_5_delay_17_41 <= io_A_Valid_5_delay_16_42;
    io_A_Valid_5_delay_18_40 <= io_A_Valid_5_delay_17_41;
    io_A_Valid_5_delay_19_39 <= io_A_Valid_5_delay_18_40;
    io_A_Valid_5_delay_20_38 <= io_A_Valid_5_delay_19_39;
    io_A_Valid_5_delay_21_37 <= io_A_Valid_5_delay_20_38;
    io_A_Valid_5_delay_22_36 <= io_A_Valid_5_delay_21_37;
    io_A_Valid_5_delay_23_35 <= io_A_Valid_5_delay_22_36;
    io_A_Valid_5_delay_24_34 <= io_A_Valid_5_delay_23_35;
    io_A_Valid_5_delay_25_33 <= io_A_Valid_5_delay_24_34;
    io_A_Valid_5_delay_26_32 <= io_A_Valid_5_delay_25_33;
    io_A_Valid_5_delay_27_31 <= io_A_Valid_5_delay_26_32;
    io_A_Valid_5_delay_28_30 <= io_A_Valid_5_delay_27_31;
    io_A_Valid_5_delay_29_29 <= io_A_Valid_5_delay_28_30;
    io_A_Valid_5_delay_30_28 <= io_A_Valid_5_delay_29_29;
    io_A_Valid_5_delay_31_27 <= io_A_Valid_5_delay_30_28;
    io_A_Valid_5_delay_32_26 <= io_A_Valid_5_delay_31_27;
    io_A_Valid_5_delay_33_25 <= io_A_Valid_5_delay_32_26;
    io_A_Valid_5_delay_34_24 <= io_A_Valid_5_delay_33_25;
    io_A_Valid_5_delay_35_23 <= io_A_Valid_5_delay_34_24;
    io_A_Valid_5_delay_36_22 <= io_A_Valid_5_delay_35_23;
    io_A_Valid_5_delay_37_21 <= io_A_Valid_5_delay_36_22;
    io_A_Valid_5_delay_38_20 <= io_A_Valid_5_delay_37_21;
    io_A_Valid_5_delay_39_19 <= io_A_Valid_5_delay_38_20;
    io_A_Valid_5_delay_40_18 <= io_A_Valid_5_delay_39_19;
    io_A_Valid_5_delay_41_17 <= io_A_Valid_5_delay_40_18;
    io_A_Valid_5_delay_42_16 <= io_A_Valid_5_delay_41_17;
    io_A_Valid_5_delay_43_15 <= io_A_Valid_5_delay_42_16;
    io_A_Valid_5_delay_44_14 <= io_A_Valid_5_delay_43_15;
    io_A_Valid_5_delay_45_13 <= io_A_Valid_5_delay_44_14;
    io_A_Valid_5_delay_46_12 <= io_A_Valid_5_delay_45_13;
    io_A_Valid_5_delay_47_11 <= io_A_Valid_5_delay_46_12;
    io_A_Valid_5_delay_48_10 <= io_A_Valid_5_delay_47_11;
    io_A_Valid_5_delay_49_9 <= io_A_Valid_5_delay_48_10;
    io_A_Valid_5_delay_50_8 <= io_A_Valid_5_delay_49_9;
    io_A_Valid_5_delay_51_7 <= io_A_Valid_5_delay_50_8;
    io_A_Valid_5_delay_52_6 <= io_A_Valid_5_delay_51_7;
    io_A_Valid_5_delay_53_5 <= io_A_Valid_5_delay_52_6;
    io_A_Valid_5_delay_54_4 <= io_A_Valid_5_delay_53_5;
    io_A_Valid_5_delay_55_3 <= io_A_Valid_5_delay_54_4;
    io_A_Valid_5_delay_56_2 <= io_A_Valid_5_delay_55_3;
    io_A_Valid_5_delay_57_1 <= io_A_Valid_5_delay_56_2;
    io_A_Valid_5_delay_58 <= io_A_Valid_5_delay_57_1;
    io_B_Valid_58_delay_1_4 <= io_B_Valid_58;
    io_B_Valid_58_delay_2_3 <= io_B_Valid_58_delay_1_4;
    io_B_Valid_58_delay_3_2 <= io_B_Valid_58_delay_2_3;
    io_B_Valid_58_delay_4_1 <= io_B_Valid_58_delay_3_2;
    io_B_Valid_58_delay_5 <= io_B_Valid_58_delay_4_1;
    io_A_Valid_5_delay_1_58 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_57 <= io_A_Valid_5_delay_1_58;
    io_A_Valid_5_delay_3_56 <= io_A_Valid_5_delay_2_57;
    io_A_Valid_5_delay_4_55 <= io_A_Valid_5_delay_3_56;
    io_A_Valid_5_delay_5_54 <= io_A_Valid_5_delay_4_55;
    io_A_Valid_5_delay_6_53 <= io_A_Valid_5_delay_5_54;
    io_A_Valid_5_delay_7_52 <= io_A_Valid_5_delay_6_53;
    io_A_Valid_5_delay_8_51 <= io_A_Valid_5_delay_7_52;
    io_A_Valid_5_delay_9_50 <= io_A_Valid_5_delay_8_51;
    io_A_Valid_5_delay_10_49 <= io_A_Valid_5_delay_9_50;
    io_A_Valid_5_delay_11_48 <= io_A_Valid_5_delay_10_49;
    io_A_Valid_5_delay_12_47 <= io_A_Valid_5_delay_11_48;
    io_A_Valid_5_delay_13_46 <= io_A_Valid_5_delay_12_47;
    io_A_Valid_5_delay_14_45 <= io_A_Valid_5_delay_13_46;
    io_A_Valid_5_delay_15_44 <= io_A_Valid_5_delay_14_45;
    io_A_Valid_5_delay_16_43 <= io_A_Valid_5_delay_15_44;
    io_A_Valid_5_delay_17_42 <= io_A_Valid_5_delay_16_43;
    io_A_Valid_5_delay_18_41 <= io_A_Valid_5_delay_17_42;
    io_A_Valid_5_delay_19_40 <= io_A_Valid_5_delay_18_41;
    io_A_Valid_5_delay_20_39 <= io_A_Valid_5_delay_19_40;
    io_A_Valid_5_delay_21_38 <= io_A_Valid_5_delay_20_39;
    io_A_Valid_5_delay_22_37 <= io_A_Valid_5_delay_21_38;
    io_A_Valid_5_delay_23_36 <= io_A_Valid_5_delay_22_37;
    io_A_Valid_5_delay_24_35 <= io_A_Valid_5_delay_23_36;
    io_A_Valid_5_delay_25_34 <= io_A_Valid_5_delay_24_35;
    io_A_Valid_5_delay_26_33 <= io_A_Valid_5_delay_25_34;
    io_A_Valid_5_delay_27_32 <= io_A_Valid_5_delay_26_33;
    io_A_Valid_5_delay_28_31 <= io_A_Valid_5_delay_27_32;
    io_A_Valid_5_delay_29_30 <= io_A_Valid_5_delay_28_31;
    io_A_Valid_5_delay_30_29 <= io_A_Valid_5_delay_29_30;
    io_A_Valid_5_delay_31_28 <= io_A_Valid_5_delay_30_29;
    io_A_Valid_5_delay_32_27 <= io_A_Valid_5_delay_31_28;
    io_A_Valid_5_delay_33_26 <= io_A_Valid_5_delay_32_27;
    io_A_Valid_5_delay_34_25 <= io_A_Valid_5_delay_33_26;
    io_A_Valid_5_delay_35_24 <= io_A_Valid_5_delay_34_25;
    io_A_Valid_5_delay_36_23 <= io_A_Valid_5_delay_35_24;
    io_A_Valid_5_delay_37_22 <= io_A_Valid_5_delay_36_23;
    io_A_Valid_5_delay_38_21 <= io_A_Valid_5_delay_37_22;
    io_A_Valid_5_delay_39_20 <= io_A_Valid_5_delay_38_21;
    io_A_Valid_5_delay_40_19 <= io_A_Valid_5_delay_39_20;
    io_A_Valid_5_delay_41_18 <= io_A_Valid_5_delay_40_19;
    io_A_Valid_5_delay_42_17 <= io_A_Valid_5_delay_41_18;
    io_A_Valid_5_delay_43_16 <= io_A_Valid_5_delay_42_17;
    io_A_Valid_5_delay_44_15 <= io_A_Valid_5_delay_43_16;
    io_A_Valid_5_delay_45_14 <= io_A_Valid_5_delay_44_15;
    io_A_Valid_5_delay_46_13 <= io_A_Valid_5_delay_45_14;
    io_A_Valid_5_delay_47_12 <= io_A_Valid_5_delay_46_13;
    io_A_Valid_5_delay_48_11 <= io_A_Valid_5_delay_47_12;
    io_A_Valid_5_delay_49_10 <= io_A_Valid_5_delay_48_11;
    io_A_Valid_5_delay_50_9 <= io_A_Valid_5_delay_49_10;
    io_A_Valid_5_delay_51_8 <= io_A_Valid_5_delay_50_9;
    io_A_Valid_5_delay_52_7 <= io_A_Valid_5_delay_51_8;
    io_A_Valid_5_delay_53_6 <= io_A_Valid_5_delay_52_7;
    io_A_Valid_5_delay_54_5 <= io_A_Valid_5_delay_53_6;
    io_A_Valid_5_delay_55_4 <= io_A_Valid_5_delay_54_5;
    io_A_Valid_5_delay_56_3 <= io_A_Valid_5_delay_55_4;
    io_A_Valid_5_delay_57_2 <= io_A_Valid_5_delay_56_3;
    io_A_Valid_5_delay_58_1 <= io_A_Valid_5_delay_57_2;
    io_A_Valid_5_delay_59 <= io_A_Valid_5_delay_58_1;
    io_B_Valid_59_delay_1_4 <= io_B_Valid_59;
    io_B_Valid_59_delay_2_3 <= io_B_Valid_59_delay_1_4;
    io_B_Valid_59_delay_3_2 <= io_B_Valid_59_delay_2_3;
    io_B_Valid_59_delay_4_1 <= io_B_Valid_59_delay_3_2;
    io_B_Valid_59_delay_5 <= io_B_Valid_59_delay_4_1;
    io_A_Valid_5_delay_1_59 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_58 <= io_A_Valid_5_delay_1_59;
    io_A_Valid_5_delay_3_57 <= io_A_Valid_5_delay_2_58;
    io_A_Valid_5_delay_4_56 <= io_A_Valid_5_delay_3_57;
    io_A_Valid_5_delay_5_55 <= io_A_Valid_5_delay_4_56;
    io_A_Valid_5_delay_6_54 <= io_A_Valid_5_delay_5_55;
    io_A_Valid_5_delay_7_53 <= io_A_Valid_5_delay_6_54;
    io_A_Valid_5_delay_8_52 <= io_A_Valid_5_delay_7_53;
    io_A_Valid_5_delay_9_51 <= io_A_Valid_5_delay_8_52;
    io_A_Valid_5_delay_10_50 <= io_A_Valid_5_delay_9_51;
    io_A_Valid_5_delay_11_49 <= io_A_Valid_5_delay_10_50;
    io_A_Valid_5_delay_12_48 <= io_A_Valid_5_delay_11_49;
    io_A_Valid_5_delay_13_47 <= io_A_Valid_5_delay_12_48;
    io_A_Valid_5_delay_14_46 <= io_A_Valid_5_delay_13_47;
    io_A_Valid_5_delay_15_45 <= io_A_Valid_5_delay_14_46;
    io_A_Valid_5_delay_16_44 <= io_A_Valid_5_delay_15_45;
    io_A_Valid_5_delay_17_43 <= io_A_Valid_5_delay_16_44;
    io_A_Valid_5_delay_18_42 <= io_A_Valid_5_delay_17_43;
    io_A_Valid_5_delay_19_41 <= io_A_Valid_5_delay_18_42;
    io_A_Valid_5_delay_20_40 <= io_A_Valid_5_delay_19_41;
    io_A_Valid_5_delay_21_39 <= io_A_Valid_5_delay_20_40;
    io_A_Valid_5_delay_22_38 <= io_A_Valid_5_delay_21_39;
    io_A_Valid_5_delay_23_37 <= io_A_Valid_5_delay_22_38;
    io_A_Valid_5_delay_24_36 <= io_A_Valid_5_delay_23_37;
    io_A_Valid_5_delay_25_35 <= io_A_Valid_5_delay_24_36;
    io_A_Valid_5_delay_26_34 <= io_A_Valid_5_delay_25_35;
    io_A_Valid_5_delay_27_33 <= io_A_Valid_5_delay_26_34;
    io_A_Valid_5_delay_28_32 <= io_A_Valid_5_delay_27_33;
    io_A_Valid_5_delay_29_31 <= io_A_Valid_5_delay_28_32;
    io_A_Valid_5_delay_30_30 <= io_A_Valid_5_delay_29_31;
    io_A_Valid_5_delay_31_29 <= io_A_Valid_5_delay_30_30;
    io_A_Valid_5_delay_32_28 <= io_A_Valid_5_delay_31_29;
    io_A_Valid_5_delay_33_27 <= io_A_Valid_5_delay_32_28;
    io_A_Valid_5_delay_34_26 <= io_A_Valid_5_delay_33_27;
    io_A_Valid_5_delay_35_25 <= io_A_Valid_5_delay_34_26;
    io_A_Valid_5_delay_36_24 <= io_A_Valid_5_delay_35_25;
    io_A_Valid_5_delay_37_23 <= io_A_Valid_5_delay_36_24;
    io_A_Valid_5_delay_38_22 <= io_A_Valid_5_delay_37_23;
    io_A_Valid_5_delay_39_21 <= io_A_Valid_5_delay_38_22;
    io_A_Valid_5_delay_40_20 <= io_A_Valid_5_delay_39_21;
    io_A_Valid_5_delay_41_19 <= io_A_Valid_5_delay_40_20;
    io_A_Valid_5_delay_42_18 <= io_A_Valid_5_delay_41_19;
    io_A_Valid_5_delay_43_17 <= io_A_Valid_5_delay_42_18;
    io_A_Valid_5_delay_44_16 <= io_A_Valid_5_delay_43_17;
    io_A_Valid_5_delay_45_15 <= io_A_Valid_5_delay_44_16;
    io_A_Valid_5_delay_46_14 <= io_A_Valid_5_delay_45_15;
    io_A_Valid_5_delay_47_13 <= io_A_Valid_5_delay_46_14;
    io_A_Valid_5_delay_48_12 <= io_A_Valid_5_delay_47_13;
    io_A_Valid_5_delay_49_11 <= io_A_Valid_5_delay_48_12;
    io_A_Valid_5_delay_50_10 <= io_A_Valid_5_delay_49_11;
    io_A_Valid_5_delay_51_9 <= io_A_Valid_5_delay_50_10;
    io_A_Valid_5_delay_52_8 <= io_A_Valid_5_delay_51_9;
    io_A_Valid_5_delay_53_7 <= io_A_Valid_5_delay_52_8;
    io_A_Valid_5_delay_54_6 <= io_A_Valid_5_delay_53_7;
    io_A_Valid_5_delay_55_5 <= io_A_Valid_5_delay_54_6;
    io_A_Valid_5_delay_56_4 <= io_A_Valid_5_delay_55_5;
    io_A_Valid_5_delay_57_3 <= io_A_Valid_5_delay_56_4;
    io_A_Valid_5_delay_58_2 <= io_A_Valid_5_delay_57_3;
    io_A_Valid_5_delay_59_1 <= io_A_Valid_5_delay_58_2;
    io_A_Valid_5_delay_60 <= io_A_Valid_5_delay_59_1;
    io_B_Valid_60_delay_1_4 <= io_B_Valid_60;
    io_B_Valid_60_delay_2_3 <= io_B_Valid_60_delay_1_4;
    io_B_Valid_60_delay_3_2 <= io_B_Valid_60_delay_2_3;
    io_B_Valid_60_delay_4_1 <= io_B_Valid_60_delay_3_2;
    io_B_Valid_60_delay_5 <= io_B_Valid_60_delay_4_1;
    io_A_Valid_5_delay_1_60 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_59 <= io_A_Valid_5_delay_1_60;
    io_A_Valid_5_delay_3_58 <= io_A_Valid_5_delay_2_59;
    io_A_Valid_5_delay_4_57 <= io_A_Valid_5_delay_3_58;
    io_A_Valid_5_delay_5_56 <= io_A_Valid_5_delay_4_57;
    io_A_Valid_5_delay_6_55 <= io_A_Valid_5_delay_5_56;
    io_A_Valid_5_delay_7_54 <= io_A_Valid_5_delay_6_55;
    io_A_Valid_5_delay_8_53 <= io_A_Valid_5_delay_7_54;
    io_A_Valid_5_delay_9_52 <= io_A_Valid_5_delay_8_53;
    io_A_Valid_5_delay_10_51 <= io_A_Valid_5_delay_9_52;
    io_A_Valid_5_delay_11_50 <= io_A_Valid_5_delay_10_51;
    io_A_Valid_5_delay_12_49 <= io_A_Valid_5_delay_11_50;
    io_A_Valid_5_delay_13_48 <= io_A_Valid_5_delay_12_49;
    io_A_Valid_5_delay_14_47 <= io_A_Valid_5_delay_13_48;
    io_A_Valid_5_delay_15_46 <= io_A_Valid_5_delay_14_47;
    io_A_Valid_5_delay_16_45 <= io_A_Valid_5_delay_15_46;
    io_A_Valid_5_delay_17_44 <= io_A_Valid_5_delay_16_45;
    io_A_Valid_5_delay_18_43 <= io_A_Valid_5_delay_17_44;
    io_A_Valid_5_delay_19_42 <= io_A_Valid_5_delay_18_43;
    io_A_Valid_5_delay_20_41 <= io_A_Valid_5_delay_19_42;
    io_A_Valid_5_delay_21_40 <= io_A_Valid_5_delay_20_41;
    io_A_Valid_5_delay_22_39 <= io_A_Valid_5_delay_21_40;
    io_A_Valid_5_delay_23_38 <= io_A_Valid_5_delay_22_39;
    io_A_Valid_5_delay_24_37 <= io_A_Valid_5_delay_23_38;
    io_A_Valid_5_delay_25_36 <= io_A_Valid_5_delay_24_37;
    io_A_Valid_5_delay_26_35 <= io_A_Valid_5_delay_25_36;
    io_A_Valid_5_delay_27_34 <= io_A_Valid_5_delay_26_35;
    io_A_Valid_5_delay_28_33 <= io_A_Valid_5_delay_27_34;
    io_A_Valid_5_delay_29_32 <= io_A_Valid_5_delay_28_33;
    io_A_Valid_5_delay_30_31 <= io_A_Valid_5_delay_29_32;
    io_A_Valid_5_delay_31_30 <= io_A_Valid_5_delay_30_31;
    io_A_Valid_5_delay_32_29 <= io_A_Valid_5_delay_31_30;
    io_A_Valid_5_delay_33_28 <= io_A_Valid_5_delay_32_29;
    io_A_Valid_5_delay_34_27 <= io_A_Valid_5_delay_33_28;
    io_A_Valid_5_delay_35_26 <= io_A_Valid_5_delay_34_27;
    io_A_Valid_5_delay_36_25 <= io_A_Valid_5_delay_35_26;
    io_A_Valid_5_delay_37_24 <= io_A_Valid_5_delay_36_25;
    io_A_Valid_5_delay_38_23 <= io_A_Valid_5_delay_37_24;
    io_A_Valid_5_delay_39_22 <= io_A_Valid_5_delay_38_23;
    io_A_Valid_5_delay_40_21 <= io_A_Valid_5_delay_39_22;
    io_A_Valid_5_delay_41_20 <= io_A_Valid_5_delay_40_21;
    io_A_Valid_5_delay_42_19 <= io_A_Valid_5_delay_41_20;
    io_A_Valid_5_delay_43_18 <= io_A_Valid_5_delay_42_19;
    io_A_Valid_5_delay_44_17 <= io_A_Valid_5_delay_43_18;
    io_A_Valid_5_delay_45_16 <= io_A_Valid_5_delay_44_17;
    io_A_Valid_5_delay_46_15 <= io_A_Valid_5_delay_45_16;
    io_A_Valid_5_delay_47_14 <= io_A_Valid_5_delay_46_15;
    io_A_Valid_5_delay_48_13 <= io_A_Valid_5_delay_47_14;
    io_A_Valid_5_delay_49_12 <= io_A_Valid_5_delay_48_13;
    io_A_Valid_5_delay_50_11 <= io_A_Valid_5_delay_49_12;
    io_A_Valid_5_delay_51_10 <= io_A_Valid_5_delay_50_11;
    io_A_Valid_5_delay_52_9 <= io_A_Valid_5_delay_51_10;
    io_A_Valid_5_delay_53_8 <= io_A_Valid_5_delay_52_9;
    io_A_Valid_5_delay_54_7 <= io_A_Valid_5_delay_53_8;
    io_A_Valid_5_delay_55_6 <= io_A_Valid_5_delay_54_7;
    io_A_Valid_5_delay_56_5 <= io_A_Valid_5_delay_55_6;
    io_A_Valid_5_delay_57_4 <= io_A_Valid_5_delay_56_5;
    io_A_Valid_5_delay_58_3 <= io_A_Valid_5_delay_57_4;
    io_A_Valid_5_delay_59_2 <= io_A_Valid_5_delay_58_3;
    io_A_Valid_5_delay_60_1 <= io_A_Valid_5_delay_59_2;
    io_A_Valid_5_delay_61 <= io_A_Valid_5_delay_60_1;
    io_B_Valid_61_delay_1_4 <= io_B_Valid_61;
    io_B_Valid_61_delay_2_3 <= io_B_Valid_61_delay_1_4;
    io_B_Valid_61_delay_3_2 <= io_B_Valid_61_delay_2_3;
    io_B_Valid_61_delay_4_1 <= io_B_Valid_61_delay_3_2;
    io_B_Valid_61_delay_5 <= io_B_Valid_61_delay_4_1;
    io_A_Valid_5_delay_1_61 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_60 <= io_A_Valid_5_delay_1_61;
    io_A_Valid_5_delay_3_59 <= io_A_Valid_5_delay_2_60;
    io_A_Valid_5_delay_4_58 <= io_A_Valid_5_delay_3_59;
    io_A_Valid_5_delay_5_57 <= io_A_Valid_5_delay_4_58;
    io_A_Valid_5_delay_6_56 <= io_A_Valid_5_delay_5_57;
    io_A_Valid_5_delay_7_55 <= io_A_Valid_5_delay_6_56;
    io_A_Valid_5_delay_8_54 <= io_A_Valid_5_delay_7_55;
    io_A_Valid_5_delay_9_53 <= io_A_Valid_5_delay_8_54;
    io_A_Valid_5_delay_10_52 <= io_A_Valid_5_delay_9_53;
    io_A_Valid_5_delay_11_51 <= io_A_Valid_5_delay_10_52;
    io_A_Valid_5_delay_12_50 <= io_A_Valid_5_delay_11_51;
    io_A_Valid_5_delay_13_49 <= io_A_Valid_5_delay_12_50;
    io_A_Valid_5_delay_14_48 <= io_A_Valid_5_delay_13_49;
    io_A_Valid_5_delay_15_47 <= io_A_Valid_5_delay_14_48;
    io_A_Valid_5_delay_16_46 <= io_A_Valid_5_delay_15_47;
    io_A_Valid_5_delay_17_45 <= io_A_Valid_5_delay_16_46;
    io_A_Valid_5_delay_18_44 <= io_A_Valid_5_delay_17_45;
    io_A_Valid_5_delay_19_43 <= io_A_Valid_5_delay_18_44;
    io_A_Valid_5_delay_20_42 <= io_A_Valid_5_delay_19_43;
    io_A_Valid_5_delay_21_41 <= io_A_Valid_5_delay_20_42;
    io_A_Valid_5_delay_22_40 <= io_A_Valid_5_delay_21_41;
    io_A_Valid_5_delay_23_39 <= io_A_Valid_5_delay_22_40;
    io_A_Valid_5_delay_24_38 <= io_A_Valid_5_delay_23_39;
    io_A_Valid_5_delay_25_37 <= io_A_Valid_5_delay_24_38;
    io_A_Valid_5_delay_26_36 <= io_A_Valid_5_delay_25_37;
    io_A_Valid_5_delay_27_35 <= io_A_Valid_5_delay_26_36;
    io_A_Valid_5_delay_28_34 <= io_A_Valid_5_delay_27_35;
    io_A_Valid_5_delay_29_33 <= io_A_Valid_5_delay_28_34;
    io_A_Valid_5_delay_30_32 <= io_A_Valid_5_delay_29_33;
    io_A_Valid_5_delay_31_31 <= io_A_Valid_5_delay_30_32;
    io_A_Valid_5_delay_32_30 <= io_A_Valid_5_delay_31_31;
    io_A_Valid_5_delay_33_29 <= io_A_Valid_5_delay_32_30;
    io_A_Valid_5_delay_34_28 <= io_A_Valid_5_delay_33_29;
    io_A_Valid_5_delay_35_27 <= io_A_Valid_5_delay_34_28;
    io_A_Valid_5_delay_36_26 <= io_A_Valid_5_delay_35_27;
    io_A_Valid_5_delay_37_25 <= io_A_Valid_5_delay_36_26;
    io_A_Valid_5_delay_38_24 <= io_A_Valid_5_delay_37_25;
    io_A_Valid_5_delay_39_23 <= io_A_Valid_5_delay_38_24;
    io_A_Valid_5_delay_40_22 <= io_A_Valid_5_delay_39_23;
    io_A_Valid_5_delay_41_21 <= io_A_Valid_5_delay_40_22;
    io_A_Valid_5_delay_42_20 <= io_A_Valid_5_delay_41_21;
    io_A_Valid_5_delay_43_19 <= io_A_Valid_5_delay_42_20;
    io_A_Valid_5_delay_44_18 <= io_A_Valid_5_delay_43_19;
    io_A_Valid_5_delay_45_17 <= io_A_Valid_5_delay_44_18;
    io_A_Valid_5_delay_46_16 <= io_A_Valid_5_delay_45_17;
    io_A_Valid_5_delay_47_15 <= io_A_Valid_5_delay_46_16;
    io_A_Valid_5_delay_48_14 <= io_A_Valid_5_delay_47_15;
    io_A_Valid_5_delay_49_13 <= io_A_Valid_5_delay_48_14;
    io_A_Valid_5_delay_50_12 <= io_A_Valid_5_delay_49_13;
    io_A_Valid_5_delay_51_11 <= io_A_Valid_5_delay_50_12;
    io_A_Valid_5_delay_52_10 <= io_A_Valid_5_delay_51_11;
    io_A_Valid_5_delay_53_9 <= io_A_Valid_5_delay_52_10;
    io_A_Valid_5_delay_54_8 <= io_A_Valid_5_delay_53_9;
    io_A_Valid_5_delay_55_7 <= io_A_Valid_5_delay_54_8;
    io_A_Valid_5_delay_56_6 <= io_A_Valid_5_delay_55_7;
    io_A_Valid_5_delay_57_5 <= io_A_Valid_5_delay_56_6;
    io_A_Valid_5_delay_58_4 <= io_A_Valid_5_delay_57_5;
    io_A_Valid_5_delay_59_3 <= io_A_Valid_5_delay_58_4;
    io_A_Valid_5_delay_60_2 <= io_A_Valid_5_delay_59_3;
    io_A_Valid_5_delay_61_1 <= io_A_Valid_5_delay_60_2;
    io_A_Valid_5_delay_62 <= io_A_Valid_5_delay_61_1;
    io_B_Valid_62_delay_1_4 <= io_B_Valid_62;
    io_B_Valid_62_delay_2_3 <= io_B_Valid_62_delay_1_4;
    io_B_Valid_62_delay_3_2 <= io_B_Valid_62_delay_2_3;
    io_B_Valid_62_delay_4_1 <= io_B_Valid_62_delay_3_2;
    io_B_Valid_62_delay_5 <= io_B_Valid_62_delay_4_1;
    io_A_Valid_5_delay_1_62 <= io_A_Valid_5;
    io_A_Valid_5_delay_2_61 <= io_A_Valid_5_delay_1_62;
    io_A_Valid_5_delay_3_60 <= io_A_Valid_5_delay_2_61;
    io_A_Valid_5_delay_4_59 <= io_A_Valid_5_delay_3_60;
    io_A_Valid_5_delay_5_58 <= io_A_Valid_5_delay_4_59;
    io_A_Valid_5_delay_6_57 <= io_A_Valid_5_delay_5_58;
    io_A_Valid_5_delay_7_56 <= io_A_Valid_5_delay_6_57;
    io_A_Valid_5_delay_8_55 <= io_A_Valid_5_delay_7_56;
    io_A_Valid_5_delay_9_54 <= io_A_Valid_5_delay_8_55;
    io_A_Valid_5_delay_10_53 <= io_A_Valid_5_delay_9_54;
    io_A_Valid_5_delay_11_52 <= io_A_Valid_5_delay_10_53;
    io_A_Valid_5_delay_12_51 <= io_A_Valid_5_delay_11_52;
    io_A_Valid_5_delay_13_50 <= io_A_Valid_5_delay_12_51;
    io_A_Valid_5_delay_14_49 <= io_A_Valid_5_delay_13_50;
    io_A_Valid_5_delay_15_48 <= io_A_Valid_5_delay_14_49;
    io_A_Valid_5_delay_16_47 <= io_A_Valid_5_delay_15_48;
    io_A_Valid_5_delay_17_46 <= io_A_Valid_5_delay_16_47;
    io_A_Valid_5_delay_18_45 <= io_A_Valid_5_delay_17_46;
    io_A_Valid_5_delay_19_44 <= io_A_Valid_5_delay_18_45;
    io_A_Valid_5_delay_20_43 <= io_A_Valid_5_delay_19_44;
    io_A_Valid_5_delay_21_42 <= io_A_Valid_5_delay_20_43;
    io_A_Valid_5_delay_22_41 <= io_A_Valid_5_delay_21_42;
    io_A_Valid_5_delay_23_40 <= io_A_Valid_5_delay_22_41;
    io_A_Valid_5_delay_24_39 <= io_A_Valid_5_delay_23_40;
    io_A_Valid_5_delay_25_38 <= io_A_Valid_5_delay_24_39;
    io_A_Valid_5_delay_26_37 <= io_A_Valid_5_delay_25_38;
    io_A_Valid_5_delay_27_36 <= io_A_Valid_5_delay_26_37;
    io_A_Valid_5_delay_28_35 <= io_A_Valid_5_delay_27_36;
    io_A_Valid_5_delay_29_34 <= io_A_Valid_5_delay_28_35;
    io_A_Valid_5_delay_30_33 <= io_A_Valid_5_delay_29_34;
    io_A_Valid_5_delay_31_32 <= io_A_Valid_5_delay_30_33;
    io_A_Valid_5_delay_32_31 <= io_A_Valid_5_delay_31_32;
    io_A_Valid_5_delay_33_30 <= io_A_Valid_5_delay_32_31;
    io_A_Valid_5_delay_34_29 <= io_A_Valid_5_delay_33_30;
    io_A_Valid_5_delay_35_28 <= io_A_Valid_5_delay_34_29;
    io_A_Valid_5_delay_36_27 <= io_A_Valid_5_delay_35_28;
    io_A_Valid_5_delay_37_26 <= io_A_Valid_5_delay_36_27;
    io_A_Valid_5_delay_38_25 <= io_A_Valid_5_delay_37_26;
    io_A_Valid_5_delay_39_24 <= io_A_Valid_5_delay_38_25;
    io_A_Valid_5_delay_40_23 <= io_A_Valid_5_delay_39_24;
    io_A_Valid_5_delay_41_22 <= io_A_Valid_5_delay_40_23;
    io_A_Valid_5_delay_42_21 <= io_A_Valid_5_delay_41_22;
    io_A_Valid_5_delay_43_20 <= io_A_Valid_5_delay_42_21;
    io_A_Valid_5_delay_44_19 <= io_A_Valid_5_delay_43_20;
    io_A_Valid_5_delay_45_18 <= io_A_Valid_5_delay_44_19;
    io_A_Valid_5_delay_46_17 <= io_A_Valid_5_delay_45_18;
    io_A_Valid_5_delay_47_16 <= io_A_Valid_5_delay_46_17;
    io_A_Valid_5_delay_48_15 <= io_A_Valid_5_delay_47_16;
    io_A_Valid_5_delay_49_14 <= io_A_Valid_5_delay_48_15;
    io_A_Valid_5_delay_50_13 <= io_A_Valid_5_delay_49_14;
    io_A_Valid_5_delay_51_12 <= io_A_Valid_5_delay_50_13;
    io_A_Valid_5_delay_52_11 <= io_A_Valid_5_delay_51_12;
    io_A_Valid_5_delay_53_10 <= io_A_Valid_5_delay_52_11;
    io_A_Valid_5_delay_54_9 <= io_A_Valid_5_delay_53_10;
    io_A_Valid_5_delay_55_8 <= io_A_Valid_5_delay_54_9;
    io_A_Valid_5_delay_56_7 <= io_A_Valid_5_delay_55_8;
    io_A_Valid_5_delay_57_6 <= io_A_Valid_5_delay_56_7;
    io_A_Valid_5_delay_58_5 <= io_A_Valid_5_delay_57_6;
    io_A_Valid_5_delay_59_4 <= io_A_Valid_5_delay_58_5;
    io_A_Valid_5_delay_60_3 <= io_A_Valid_5_delay_59_4;
    io_A_Valid_5_delay_61_2 <= io_A_Valid_5_delay_60_3;
    io_A_Valid_5_delay_62_1 <= io_A_Valid_5_delay_61_2;
    io_A_Valid_5_delay_63 <= io_A_Valid_5_delay_62_1;
    io_B_Valid_63_delay_1_4 <= io_B_Valid_63;
    io_B_Valid_63_delay_2_3 <= io_B_Valid_63_delay_1_4;
    io_B_Valid_63_delay_3_2 <= io_B_Valid_63_delay_2_3;
    io_B_Valid_63_delay_4_1 <= io_B_Valid_63_delay_3_2;
    io_B_Valid_63_delay_5 <= io_B_Valid_63_delay_4_1;
    io_B_Valid_0_delay_1_5 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_4 <= io_B_Valid_0_delay_1_5;
    io_B_Valid_0_delay_3_3 <= io_B_Valid_0_delay_2_4;
    io_B_Valid_0_delay_4_2 <= io_B_Valid_0_delay_3_3;
    io_B_Valid_0_delay_5_1 <= io_B_Valid_0_delay_4_2;
    io_B_Valid_0_delay_6 <= io_B_Valid_0_delay_5_1;
    io_A_Valid_6_delay_1 <= io_A_Valid_6;
    io_B_Valid_1_delay_1_5 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_4 <= io_B_Valid_1_delay_1_5;
    io_B_Valid_1_delay_3_3 <= io_B_Valid_1_delay_2_4;
    io_B_Valid_1_delay_4_2 <= io_B_Valid_1_delay_3_3;
    io_B_Valid_1_delay_5_1 <= io_B_Valid_1_delay_4_2;
    io_B_Valid_1_delay_6 <= io_B_Valid_1_delay_5_1;
    io_A_Valid_6_delay_1_1 <= io_A_Valid_6;
    io_A_Valid_6_delay_2 <= io_A_Valid_6_delay_1_1;
    io_B_Valid_2_delay_1_5 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_4 <= io_B_Valid_2_delay_1_5;
    io_B_Valid_2_delay_3_3 <= io_B_Valid_2_delay_2_4;
    io_B_Valid_2_delay_4_2 <= io_B_Valid_2_delay_3_3;
    io_B_Valid_2_delay_5_1 <= io_B_Valid_2_delay_4_2;
    io_B_Valid_2_delay_6 <= io_B_Valid_2_delay_5_1;
    io_A_Valid_6_delay_1_2 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_1 <= io_A_Valid_6_delay_1_2;
    io_A_Valid_6_delay_3 <= io_A_Valid_6_delay_2_1;
    io_B_Valid_3_delay_1_5 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_4 <= io_B_Valid_3_delay_1_5;
    io_B_Valid_3_delay_3_3 <= io_B_Valid_3_delay_2_4;
    io_B_Valid_3_delay_4_2 <= io_B_Valid_3_delay_3_3;
    io_B_Valid_3_delay_5_1 <= io_B_Valid_3_delay_4_2;
    io_B_Valid_3_delay_6 <= io_B_Valid_3_delay_5_1;
    io_A_Valid_6_delay_1_3 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_2 <= io_A_Valid_6_delay_1_3;
    io_A_Valid_6_delay_3_1 <= io_A_Valid_6_delay_2_2;
    io_A_Valid_6_delay_4 <= io_A_Valid_6_delay_3_1;
    io_B_Valid_4_delay_1_5 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_4 <= io_B_Valid_4_delay_1_5;
    io_B_Valid_4_delay_3_3 <= io_B_Valid_4_delay_2_4;
    io_B_Valid_4_delay_4_2 <= io_B_Valid_4_delay_3_3;
    io_B_Valid_4_delay_5_1 <= io_B_Valid_4_delay_4_2;
    io_B_Valid_4_delay_6 <= io_B_Valid_4_delay_5_1;
    io_A_Valid_6_delay_1_4 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_3 <= io_A_Valid_6_delay_1_4;
    io_A_Valid_6_delay_3_2 <= io_A_Valid_6_delay_2_3;
    io_A_Valid_6_delay_4_1 <= io_A_Valid_6_delay_3_2;
    io_A_Valid_6_delay_5 <= io_A_Valid_6_delay_4_1;
    io_B_Valid_5_delay_1_5 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_4 <= io_B_Valid_5_delay_1_5;
    io_B_Valid_5_delay_3_3 <= io_B_Valid_5_delay_2_4;
    io_B_Valid_5_delay_4_2 <= io_B_Valid_5_delay_3_3;
    io_B_Valid_5_delay_5_1 <= io_B_Valid_5_delay_4_2;
    io_B_Valid_5_delay_6 <= io_B_Valid_5_delay_5_1;
    io_A_Valid_6_delay_1_5 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_4 <= io_A_Valid_6_delay_1_5;
    io_A_Valid_6_delay_3_3 <= io_A_Valid_6_delay_2_4;
    io_A_Valid_6_delay_4_2 <= io_A_Valid_6_delay_3_3;
    io_A_Valid_6_delay_5_1 <= io_A_Valid_6_delay_4_2;
    io_A_Valid_6_delay_6 <= io_A_Valid_6_delay_5_1;
    io_B_Valid_6_delay_1_5 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_4 <= io_B_Valid_6_delay_1_5;
    io_B_Valid_6_delay_3_3 <= io_B_Valid_6_delay_2_4;
    io_B_Valid_6_delay_4_2 <= io_B_Valid_6_delay_3_3;
    io_B_Valid_6_delay_5_1 <= io_B_Valid_6_delay_4_2;
    io_B_Valid_6_delay_6 <= io_B_Valid_6_delay_5_1;
    io_A_Valid_6_delay_1_6 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_5 <= io_A_Valid_6_delay_1_6;
    io_A_Valid_6_delay_3_4 <= io_A_Valid_6_delay_2_5;
    io_A_Valid_6_delay_4_3 <= io_A_Valid_6_delay_3_4;
    io_A_Valid_6_delay_5_2 <= io_A_Valid_6_delay_4_3;
    io_A_Valid_6_delay_6_1 <= io_A_Valid_6_delay_5_2;
    io_A_Valid_6_delay_7 <= io_A_Valid_6_delay_6_1;
    io_B_Valid_7_delay_1_5 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_4 <= io_B_Valid_7_delay_1_5;
    io_B_Valid_7_delay_3_3 <= io_B_Valid_7_delay_2_4;
    io_B_Valid_7_delay_4_2 <= io_B_Valid_7_delay_3_3;
    io_B_Valid_7_delay_5_1 <= io_B_Valid_7_delay_4_2;
    io_B_Valid_7_delay_6 <= io_B_Valid_7_delay_5_1;
    io_A_Valid_6_delay_1_7 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_6 <= io_A_Valid_6_delay_1_7;
    io_A_Valid_6_delay_3_5 <= io_A_Valid_6_delay_2_6;
    io_A_Valid_6_delay_4_4 <= io_A_Valid_6_delay_3_5;
    io_A_Valid_6_delay_5_3 <= io_A_Valid_6_delay_4_4;
    io_A_Valid_6_delay_6_2 <= io_A_Valid_6_delay_5_3;
    io_A_Valid_6_delay_7_1 <= io_A_Valid_6_delay_6_2;
    io_A_Valid_6_delay_8 <= io_A_Valid_6_delay_7_1;
    io_B_Valid_8_delay_1_5 <= io_B_Valid_8;
    io_B_Valid_8_delay_2_4 <= io_B_Valid_8_delay_1_5;
    io_B_Valid_8_delay_3_3 <= io_B_Valid_8_delay_2_4;
    io_B_Valid_8_delay_4_2 <= io_B_Valid_8_delay_3_3;
    io_B_Valid_8_delay_5_1 <= io_B_Valid_8_delay_4_2;
    io_B_Valid_8_delay_6 <= io_B_Valid_8_delay_5_1;
    io_A_Valid_6_delay_1_8 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_7 <= io_A_Valid_6_delay_1_8;
    io_A_Valid_6_delay_3_6 <= io_A_Valid_6_delay_2_7;
    io_A_Valid_6_delay_4_5 <= io_A_Valid_6_delay_3_6;
    io_A_Valid_6_delay_5_4 <= io_A_Valid_6_delay_4_5;
    io_A_Valid_6_delay_6_3 <= io_A_Valid_6_delay_5_4;
    io_A_Valid_6_delay_7_2 <= io_A_Valid_6_delay_6_3;
    io_A_Valid_6_delay_8_1 <= io_A_Valid_6_delay_7_2;
    io_A_Valid_6_delay_9 <= io_A_Valid_6_delay_8_1;
    io_B_Valid_9_delay_1_5 <= io_B_Valid_9;
    io_B_Valid_9_delay_2_4 <= io_B_Valid_9_delay_1_5;
    io_B_Valid_9_delay_3_3 <= io_B_Valid_9_delay_2_4;
    io_B_Valid_9_delay_4_2 <= io_B_Valid_9_delay_3_3;
    io_B_Valid_9_delay_5_1 <= io_B_Valid_9_delay_4_2;
    io_B_Valid_9_delay_6 <= io_B_Valid_9_delay_5_1;
    io_A_Valid_6_delay_1_9 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_8 <= io_A_Valid_6_delay_1_9;
    io_A_Valid_6_delay_3_7 <= io_A_Valid_6_delay_2_8;
    io_A_Valid_6_delay_4_6 <= io_A_Valid_6_delay_3_7;
    io_A_Valid_6_delay_5_5 <= io_A_Valid_6_delay_4_6;
    io_A_Valid_6_delay_6_4 <= io_A_Valid_6_delay_5_5;
    io_A_Valid_6_delay_7_3 <= io_A_Valid_6_delay_6_4;
    io_A_Valid_6_delay_8_2 <= io_A_Valid_6_delay_7_3;
    io_A_Valid_6_delay_9_1 <= io_A_Valid_6_delay_8_2;
    io_A_Valid_6_delay_10 <= io_A_Valid_6_delay_9_1;
    io_B_Valid_10_delay_1_5 <= io_B_Valid_10;
    io_B_Valid_10_delay_2_4 <= io_B_Valid_10_delay_1_5;
    io_B_Valid_10_delay_3_3 <= io_B_Valid_10_delay_2_4;
    io_B_Valid_10_delay_4_2 <= io_B_Valid_10_delay_3_3;
    io_B_Valid_10_delay_5_1 <= io_B_Valid_10_delay_4_2;
    io_B_Valid_10_delay_6 <= io_B_Valid_10_delay_5_1;
    io_A_Valid_6_delay_1_10 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_9 <= io_A_Valid_6_delay_1_10;
    io_A_Valid_6_delay_3_8 <= io_A_Valid_6_delay_2_9;
    io_A_Valid_6_delay_4_7 <= io_A_Valid_6_delay_3_8;
    io_A_Valid_6_delay_5_6 <= io_A_Valid_6_delay_4_7;
    io_A_Valid_6_delay_6_5 <= io_A_Valid_6_delay_5_6;
    io_A_Valid_6_delay_7_4 <= io_A_Valid_6_delay_6_5;
    io_A_Valid_6_delay_8_3 <= io_A_Valid_6_delay_7_4;
    io_A_Valid_6_delay_9_2 <= io_A_Valid_6_delay_8_3;
    io_A_Valid_6_delay_10_1 <= io_A_Valid_6_delay_9_2;
    io_A_Valid_6_delay_11 <= io_A_Valid_6_delay_10_1;
    io_B_Valid_11_delay_1_5 <= io_B_Valid_11;
    io_B_Valid_11_delay_2_4 <= io_B_Valid_11_delay_1_5;
    io_B_Valid_11_delay_3_3 <= io_B_Valid_11_delay_2_4;
    io_B_Valid_11_delay_4_2 <= io_B_Valid_11_delay_3_3;
    io_B_Valid_11_delay_5_1 <= io_B_Valid_11_delay_4_2;
    io_B_Valid_11_delay_6 <= io_B_Valid_11_delay_5_1;
    io_A_Valid_6_delay_1_11 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_10 <= io_A_Valid_6_delay_1_11;
    io_A_Valid_6_delay_3_9 <= io_A_Valid_6_delay_2_10;
    io_A_Valid_6_delay_4_8 <= io_A_Valid_6_delay_3_9;
    io_A_Valid_6_delay_5_7 <= io_A_Valid_6_delay_4_8;
    io_A_Valid_6_delay_6_6 <= io_A_Valid_6_delay_5_7;
    io_A_Valid_6_delay_7_5 <= io_A_Valid_6_delay_6_6;
    io_A_Valid_6_delay_8_4 <= io_A_Valid_6_delay_7_5;
    io_A_Valid_6_delay_9_3 <= io_A_Valid_6_delay_8_4;
    io_A_Valid_6_delay_10_2 <= io_A_Valid_6_delay_9_3;
    io_A_Valid_6_delay_11_1 <= io_A_Valid_6_delay_10_2;
    io_A_Valid_6_delay_12 <= io_A_Valid_6_delay_11_1;
    io_B_Valid_12_delay_1_5 <= io_B_Valid_12;
    io_B_Valid_12_delay_2_4 <= io_B_Valid_12_delay_1_5;
    io_B_Valid_12_delay_3_3 <= io_B_Valid_12_delay_2_4;
    io_B_Valid_12_delay_4_2 <= io_B_Valid_12_delay_3_3;
    io_B_Valid_12_delay_5_1 <= io_B_Valid_12_delay_4_2;
    io_B_Valid_12_delay_6 <= io_B_Valid_12_delay_5_1;
    io_A_Valid_6_delay_1_12 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_11 <= io_A_Valid_6_delay_1_12;
    io_A_Valid_6_delay_3_10 <= io_A_Valid_6_delay_2_11;
    io_A_Valid_6_delay_4_9 <= io_A_Valid_6_delay_3_10;
    io_A_Valid_6_delay_5_8 <= io_A_Valid_6_delay_4_9;
    io_A_Valid_6_delay_6_7 <= io_A_Valid_6_delay_5_8;
    io_A_Valid_6_delay_7_6 <= io_A_Valid_6_delay_6_7;
    io_A_Valid_6_delay_8_5 <= io_A_Valid_6_delay_7_6;
    io_A_Valid_6_delay_9_4 <= io_A_Valid_6_delay_8_5;
    io_A_Valid_6_delay_10_3 <= io_A_Valid_6_delay_9_4;
    io_A_Valid_6_delay_11_2 <= io_A_Valid_6_delay_10_3;
    io_A_Valid_6_delay_12_1 <= io_A_Valid_6_delay_11_2;
    io_A_Valid_6_delay_13 <= io_A_Valid_6_delay_12_1;
    io_B_Valid_13_delay_1_5 <= io_B_Valid_13;
    io_B_Valid_13_delay_2_4 <= io_B_Valid_13_delay_1_5;
    io_B_Valid_13_delay_3_3 <= io_B_Valid_13_delay_2_4;
    io_B_Valid_13_delay_4_2 <= io_B_Valid_13_delay_3_3;
    io_B_Valid_13_delay_5_1 <= io_B_Valid_13_delay_4_2;
    io_B_Valid_13_delay_6 <= io_B_Valid_13_delay_5_1;
    io_A_Valid_6_delay_1_13 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_12 <= io_A_Valid_6_delay_1_13;
    io_A_Valid_6_delay_3_11 <= io_A_Valid_6_delay_2_12;
    io_A_Valid_6_delay_4_10 <= io_A_Valid_6_delay_3_11;
    io_A_Valid_6_delay_5_9 <= io_A_Valid_6_delay_4_10;
    io_A_Valid_6_delay_6_8 <= io_A_Valid_6_delay_5_9;
    io_A_Valid_6_delay_7_7 <= io_A_Valid_6_delay_6_8;
    io_A_Valid_6_delay_8_6 <= io_A_Valid_6_delay_7_7;
    io_A_Valid_6_delay_9_5 <= io_A_Valid_6_delay_8_6;
    io_A_Valid_6_delay_10_4 <= io_A_Valid_6_delay_9_5;
    io_A_Valid_6_delay_11_3 <= io_A_Valid_6_delay_10_4;
    io_A_Valid_6_delay_12_2 <= io_A_Valid_6_delay_11_3;
    io_A_Valid_6_delay_13_1 <= io_A_Valid_6_delay_12_2;
    io_A_Valid_6_delay_14 <= io_A_Valid_6_delay_13_1;
    io_B_Valid_14_delay_1_5 <= io_B_Valid_14;
    io_B_Valid_14_delay_2_4 <= io_B_Valid_14_delay_1_5;
    io_B_Valid_14_delay_3_3 <= io_B_Valid_14_delay_2_4;
    io_B_Valid_14_delay_4_2 <= io_B_Valid_14_delay_3_3;
    io_B_Valid_14_delay_5_1 <= io_B_Valid_14_delay_4_2;
    io_B_Valid_14_delay_6 <= io_B_Valid_14_delay_5_1;
    io_A_Valid_6_delay_1_14 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_13 <= io_A_Valid_6_delay_1_14;
    io_A_Valid_6_delay_3_12 <= io_A_Valid_6_delay_2_13;
    io_A_Valid_6_delay_4_11 <= io_A_Valid_6_delay_3_12;
    io_A_Valid_6_delay_5_10 <= io_A_Valid_6_delay_4_11;
    io_A_Valid_6_delay_6_9 <= io_A_Valid_6_delay_5_10;
    io_A_Valid_6_delay_7_8 <= io_A_Valid_6_delay_6_9;
    io_A_Valid_6_delay_8_7 <= io_A_Valid_6_delay_7_8;
    io_A_Valid_6_delay_9_6 <= io_A_Valid_6_delay_8_7;
    io_A_Valid_6_delay_10_5 <= io_A_Valid_6_delay_9_6;
    io_A_Valid_6_delay_11_4 <= io_A_Valid_6_delay_10_5;
    io_A_Valid_6_delay_12_3 <= io_A_Valid_6_delay_11_4;
    io_A_Valid_6_delay_13_2 <= io_A_Valid_6_delay_12_3;
    io_A_Valid_6_delay_14_1 <= io_A_Valid_6_delay_13_2;
    io_A_Valid_6_delay_15 <= io_A_Valid_6_delay_14_1;
    io_B_Valid_15_delay_1_5 <= io_B_Valid_15;
    io_B_Valid_15_delay_2_4 <= io_B_Valid_15_delay_1_5;
    io_B_Valid_15_delay_3_3 <= io_B_Valid_15_delay_2_4;
    io_B_Valid_15_delay_4_2 <= io_B_Valid_15_delay_3_3;
    io_B_Valid_15_delay_5_1 <= io_B_Valid_15_delay_4_2;
    io_B_Valid_15_delay_6 <= io_B_Valid_15_delay_5_1;
    io_A_Valid_6_delay_1_15 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_14 <= io_A_Valid_6_delay_1_15;
    io_A_Valid_6_delay_3_13 <= io_A_Valid_6_delay_2_14;
    io_A_Valid_6_delay_4_12 <= io_A_Valid_6_delay_3_13;
    io_A_Valid_6_delay_5_11 <= io_A_Valid_6_delay_4_12;
    io_A_Valid_6_delay_6_10 <= io_A_Valid_6_delay_5_11;
    io_A_Valid_6_delay_7_9 <= io_A_Valid_6_delay_6_10;
    io_A_Valid_6_delay_8_8 <= io_A_Valid_6_delay_7_9;
    io_A_Valid_6_delay_9_7 <= io_A_Valid_6_delay_8_8;
    io_A_Valid_6_delay_10_6 <= io_A_Valid_6_delay_9_7;
    io_A_Valid_6_delay_11_5 <= io_A_Valid_6_delay_10_6;
    io_A_Valid_6_delay_12_4 <= io_A_Valid_6_delay_11_5;
    io_A_Valid_6_delay_13_3 <= io_A_Valid_6_delay_12_4;
    io_A_Valid_6_delay_14_2 <= io_A_Valid_6_delay_13_3;
    io_A_Valid_6_delay_15_1 <= io_A_Valid_6_delay_14_2;
    io_A_Valid_6_delay_16 <= io_A_Valid_6_delay_15_1;
    io_B_Valid_16_delay_1_5 <= io_B_Valid_16;
    io_B_Valid_16_delay_2_4 <= io_B_Valid_16_delay_1_5;
    io_B_Valid_16_delay_3_3 <= io_B_Valid_16_delay_2_4;
    io_B_Valid_16_delay_4_2 <= io_B_Valid_16_delay_3_3;
    io_B_Valid_16_delay_5_1 <= io_B_Valid_16_delay_4_2;
    io_B_Valid_16_delay_6 <= io_B_Valid_16_delay_5_1;
    io_A_Valid_6_delay_1_16 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_15 <= io_A_Valid_6_delay_1_16;
    io_A_Valid_6_delay_3_14 <= io_A_Valid_6_delay_2_15;
    io_A_Valid_6_delay_4_13 <= io_A_Valid_6_delay_3_14;
    io_A_Valid_6_delay_5_12 <= io_A_Valid_6_delay_4_13;
    io_A_Valid_6_delay_6_11 <= io_A_Valid_6_delay_5_12;
    io_A_Valid_6_delay_7_10 <= io_A_Valid_6_delay_6_11;
    io_A_Valid_6_delay_8_9 <= io_A_Valid_6_delay_7_10;
    io_A_Valid_6_delay_9_8 <= io_A_Valid_6_delay_8_9;
    io_A_Valid_6_delay_10_7 <= io_A_Valid_6_delay_9_8;
    io_A_Valid_6_delay_11_6 <= io_A_Valid_6_delay_10_7;
    io_A_Valid_6_delay_12_5 <= io_A_Valid_6_delay_11_6;
    io_A_Valid_6_delay_13_4 <= io_A_Valid_6_delay_12_5;
    io_A_Valid_6_delay_14_3 <= io_A_Valid_6_delay_13_4;
    io_A_Valid_6_delay_15_2 <= io_A_Valid_6_delay_14_3;
    io_A_Valid_6_delay_16_1 <= io_A_Valid_6_delay_15_2;
    io_A_Valid_6_delay_17 <= io_A_Valid_6_delay_16_1;
    io_B_Valid_17_delay_1_5 <= io_B_Valid_17;
    io_B_Valid_17_delay_2_4 <= io_B_Valid_17_delay_1_5;
    io_B_Valid_17_delay_3_3 <= io_B_Valid_17_delay_2_4;
    io_B_Valid_17_delay_4_2 <= io_B_Valid_17_delay_3_3;
    io_B_Valid_17_delay_5_1 <= io_B_Valid_17_delay_4_2;
    io_B_Valid_17_delay_6 <= io_B_Valid_17_delay_5_1;
    io_A_Valid_6_delay_1_17 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_16 <= io_A_Valid_6_delay_1_17;
    io_A_Valid_6_delay_3_15 <= io_A_Valid_6_delay_2_16;
    io_A_Valid_6_delay_4_14 <= io_A_Valid_6_delay_3_15;
    io_A_Valid_6_delay_5_13 <= io_A_Valid_6_delay_4_14;
    io_A_Valid_6_delay_6_12 <= io_A_Valid_6_delay_5_13;
    io_A_Valid_6_delay_7_11 <= io_A_Valid_6_delay_6_12;
    io_A_Valid_6_delay_8_10 <= io_A_Valid_6_delay_7_11;
    io_A_Valid_6_delay_9_9 <= io_A_Valid_6_delay_8_10;
    io_A_Valid_6_delay_10_8 <= io_A_Valid_6_delay_9_9;
    io_A_Valid_6_delay_11_7 <= io_A_Valid_6_delay_10_8;
    io_A_Valid_6_delay_12_6 <= io_A_Valid_6_delay_11_7;
    io_A_Valid_6_delay_13_5 <= io_A_Valid_6_delay_12_6;
    io_A_Valid_6_delay_14_4 <= io_A_Valid_6_delay_13_5;
    io_A_Valid_6_delay_15_3 <= io_A_Valid_6_delay_14_4;
    io_A_Valid_6_delay_16_2 <= io_A_Valid_6_delay_15_3;
    io_A_Valid_6_delay_17_1 <= io_A_Valid_6_delay_16_2;
    io_A_Valid_6_delay_18 <= io_A_Valid_6_delay_17_1;
    io_B_Valid_18_delay_1_5 <= io_B_Valid_18;
    io_B_Valid_18_delay_2_4 <= io_B_Valid_18_delay_1_5;
    io_B_Valid_18_delay_3_3 <= io_B_Valid_18_delay_2_4;
    io_B_Valid_18_delay_4_2 <= io_B_Valid_18_delay_3_3;
    io_B_Valid_18_delay_5_1 <= io_B_Valid_18_delay_4_2;
    io_B_Valid_18_delay_6 <= io_B_Valid_18_delay_5_1;
    io_A_Valid_6_delay_1_18 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_17 <= io_A_Valid_6_delay_1_18;
    io_A_Valid_6_delay_3_16 <= io_A_Valid_6_delay_2_17;
    io_A_Valid_6_delay_4_15 <= io_A_Valid_6_delay_3_16;
    io_A_Valid_6_delay_5_14 <= io_A_Valid_6_delay_4_15;
    io_A_Valid_6_delay_6_13 <= io_A_Valid_6_delay_5_14;
    io_A_Valid_6_delay_7_12 <= io_A_Valid_6_delay_6_13;
    io_A_Valid_6_delay_8_11 <= io_A_Valid_6_delay_7_12;
    io_A_Valid_6_delay_9_10 <= io_A_Valid_6_delay_8_11;
    io_A_Valid_6_delay_10_9 <= io_A_Valid_6_delay_9_10;
    io_A_Valid_6_delay_11_8 <= io_A_Valid_6_delay_10_9;
    io_A_Valid_6_delay_12_7 <= io_A_Valid_6_delay_11_8;
    io_A_Valid_6_delay_13_6 <= io_A_Valid_6_delay_12_7;
    io_A_Valid_6_delay_14_5 <= io_A_Valid_6_delay_13_6;
    io_A_Valid_6_delay_15_4 <= io_A_Valid_6_delay_14_5;
    io_A_Valid_6_delay_16_3 <= io_A_Valid_6_delay_15_4;
    io_A_Valid_6_delay_17_2 <= io_A_Valid_6_delay_16_3;
    io_A_Valid_6_delay_18_1 <= io_A_Valid_6_delay_17_2;
    io_A_Valid_6_delay_19 <= io_A_Valid_6_delay_18_1;
    io_B_Valid_19_delay_1_5 <= io_B_Valid_19;
    io_B_Valid_19_delay_2_4 <= io_B_Valid_19_delay_1_5;
    io_B_Valid_19_delay_3_3 <= io_B_Valid_19_delay_2_4;
    io_B_Valid_19_delay_4_2 <= io_B_Valid_19_delay_3_3;
    io_B_Valid_19_delay_5_1 <= io_B_Valid_19_delay_4_2;
    io_B_Valid_19_delay_6 <= io_B_Valid_19_delay_5_1;
    io_A_Valid_6_delay_1_19 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_18 <= io_A_Valid_6_delay_1_19;
    io_A_Valid_6_delay_3_17 <= io_A_Valid_6_delay_2_18;
    io_A_Valid_6_delay_4_16 <= io_A_Valid_6_delay_3_17;
    io_A_Valid_6_delay_5_15 <= io_A_Valid_6_delay_4_16;
    io_A_Valid_6_delay_6_14 <= io_A_Valid_6_delay_5_15;
    io_A_Valid_6_delay_7_13 <= io_A_Valid_6_delay_6_14;
    io_A_Valid_6_delay_8_12 <= io_A_Valid_6_delay_7_13;
    io_A_Valid_6_delay_9_11 <= io_A_Valid_6_delay_8_12;
    io_A_Valid_6_delay_10_10 <= io_A_Valid_6_delay_9_11;
    io_A_Valid_6_delay_11_9 <= io_A_Valid_6_delay_10_10;
    io_A_Valid_6_delay_12_8 <= io_A_Valid_6_delay_11_9;
    io_A_Valid_6_delay_13_7 <= io_A_Valid_6_delay_12_8;
    io_A_Valid_6_delay_14_6 <= io_A_Valid_6_delay_13_7;
    io_A_Valid_6_delay_15_5 <= io_A_Valid_6_delay_14_6;
    io_A_Valid_6_delay_16_4 <= io_A_Valid_6_delay_15_5;
    io_A_Valid_6_delay_17_3 <= io_A_Valid_6_delay_16_4;
    io_A_Valid_6_delay_18_2 <= io_A_Valid_6_delay_17_3;
    io_A_Valid_6_delay_19_1 <= io_A_Valid_6_delay_18_2;
    io_A_Valid_6_delay_20 <= io_A_Valid_6_delay_19_1;
    io_B_Valid_20_delay_1_5 <= io_B_Valid_20;
    io_B_Valid_20_delay_2_4 <= io_B_Valid_20_delay_1_5;
    io_B_Valid_20_delay_3_3 <= io_B_Valid_20_delay_2_4;
    io_B_Valid_20_delay_4_2 <= io_B_Valid_20_delay_3_3;
    io_B_Valid_20_delay_5_1 <= io_B_Valid_20_delay_4_2;
    io_B_Valid_20_delay_6 <= io_B_Valid_20_delay_5_1;
    io_A_Valid_6_delay_1_20 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_19 <= io_A_Valid_6_delay_1_20;
    io_A_Valid_6_delay_3_18 <= io_A_Valid_6_delay_2_19;
    io_A_Valid_6_delay_4_17 <= io_A_Valid_6_delay_3_18;
    io_A_Valid_6_delay_5_16 <= io_A_Valid_6_delay_4_17;
    io_A_Valid_6_delay_6_15 <= io_A_Valid_6_delay_5_16;
    io_A_Valid_6_delay_7_14 <= io_A_Valid_6_delay_6_15;
    io_A_Valid_6_delay_8_13 <= io_A_Valid_6_delay_7_14;
    io_A_Valid_6_delay_9_12 <= io_A_Valid_6_delay_8_13;
    io_A_Valid_6_delay_10_11 <= io_A_Valid_6_delay_9_12;
    io_A_Valid_6_delay_11_10 <= io_A_Valid_6_delay_10_11;
    io_A_Valid_6_delay_12_9 <= io_A_Valid_6_delay_11_10;
    io_A_Valid_6_delay_13_8 <= io_A_Valid_6_delay_12_9;
    io_A_Valid_6_delay_14_7 <= io_A_Valid_6_delay_13_8;
    io_A_Valid_6_delay_15_6 <= io_A_Valid_6_delay_14_7;
    io_A_Valid_6_delay_16_5 <= io_A_Valid_6_delay_15_6;
    io_A_Valid_6_delay_17_4 <= io_A_Valid_6_delay_16_5;
    io_A_Valid_6_delay_18_3 <= io_A_Valid_6_delay_17_4;
    io_A_Valid_6_delay_19_2 <= io_A_Valid_6_delay_18_3;
    io_A_Valid_6_delay_20_1 <= io_A_Valid_6_delay_19_2;
    io_A_Valid_6_delay_21 <= io_A_Valid_6_delay_20_1;
    io_B_Valid_21_delay_1_5 <= io_B_Valid_21;
    io_B_Valid_21_delay_2_4 <= io_B_Valid_21_delay_1_5;
    io_B_Valid_21_delay_3_3 <= io_B_Valid_21_delay_2_4;
    io_B_Valid_21_delay_4_2 <= io_B_Valid_21_delay_3_3;
    io_B_Valid_21_delay_5_1 <= io_B_Valid_21_delay_4_2;
    io_B_Valid_21_delay_6 <= io_B_Valid_21_delay_5_1;
    io_A_Valid_6_delay_1_21 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_20 <= io_A_Valid_6_delay_1_21;
    io_A_Valid_6_delay_3_19 <= io_A_Valid_6_delay_2_20;
    io_A_Valid_6_delay_4_18 <= io_A_Valid_6_delay_3_19;
    io_A_Valid_6_delay_5_17 <= io_A_Valid_6_delay_4_18;
    io_A_Valid_6_delay_6_16 <= io_A_Valid_6_delay_5_17;
    io_A_Valid_6_delay_7_15 <= io_A_Valid_6_delay_6_16;
    io_A_Valid_6_delay_8_14 <= io_A_Valid_6_delay_7_15;
    io_A_Valid_6_delay_9_13 <= io_A_Valid_6_delay_8_14;
    io_A_Valid_6_delay_10_12 <= io_A_Valid_6_delay_9_13;
    io_A_Valid_6_delay_11_11 <= io_A_Valid_6_delay_10_12;
    io_A_Valid_6_delay_12_10 <= io_A_Valid_6_delay_11_11;
    io_A_Valid_6_delay_13_9 <= io_A_Valid_6_delay_12_10;
    io_A_Valid_6_delay_14_8 <= io_A_Valid_6_delay_13_9;
    io_A_Valid_6_delay_15_7 <= io_A_Valid_6_delay_14_8;
    io_A_Valid_6_delay_16_6 <= io_A_Valid_6_delay_15_7;
    io_A_Valid_6_delay_17_5 <= io_A_Valid_6_delay_16_6;
    io_A_Valid_6_delay_18_4 <= io_A_Valid_6_delay_17_5;
    io_A_Valid_6_delay_19_3 <= io_A_Valid_6_delay_18_4;
    io_A_Valid_6_delay_20_2 <= io_A_Valid_6_delay_19_3;
    io_A_Valid_6_delay_21_1 <= io_A_Valid_6_delay_20_2;
    io_A_Valid_6_delay_22 <= io_A_Valid_6_delay_21_1;
    io_B_Valid_22_delay_1_5 <= io_B_Valid_22;
    io_B_Valid_22_delay_2_4 <= io_B_Valid_22_delay_1_5;
    io_B_Valid_22_delay_3_3 <= io_B_Valid_22_delay_2_4;
    io_B_Valid_22_delay_4_2 <= io_B_Valid_22_delay_3_3;
    io_B_Valid_22_delay_5_1 <= io_B_Valid_22_delay_4_2;
    io_B_Valid_22_delay_6 <= io_B_Valid_22_delay_5_1;
    io_A_Valid_6_delay_1_22 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_21 <= io_A_Valid_6_delay_1_22;
    io_A_Valid_6_delay_3_20 <= io_A_Valid_6_delay_2_21;
    io_A_Valid_6_delay_4_19 <= io_A_Valid_6_delay_3_20;
    io_A_Valid_6_delay_5_18 <= io_A_Valid_6_delay_4_19;
    io_A_Valid_6_delay_6_17 <= io_A_Valid_6_delay_5_18;
    io_A_Valid_6_delay_7_16 <= io_A_Valid_6_delay_6_17;
    io_A_Valid_6_delay_8_15 <= io_A_Valid_6_delay_7_16;
    io_A_Valid_6_delay_9_14 <= io_A_Valid_6_delay_8_15;
    io_A_Valid_6_delay_10_13 <= io_A_Valid_6_delay_9_14;
    io_A_Valid_6_delay_11_12 <= io_A_Valid_6_delay_10_13;
    io_A_Valid_6_delay_12_11 <= io_A_Valid_6_delay_11_12;
    io_A_Valid_6_delay_13_10 <= io_A_Valid_6_delay_12_11;
    io_A_Valid_6_delay_14_9 <= io_A_Valid_6_delay_13_10;
    io_A_Valid_6_delay_15_8 <= io_A_Valid_6_delay_14_9;
    io_A_Valid_6_delay_16_7 <= io_A_Valid_6_delay_15_8;
    io_A_Valid_6_delay_17_6 <= io_A_Valid_6_delay_16_7;
    io_A_Valid_6_delay_18_5 <= io_A_Valid_6_delay_17_6;
    io_A_Valid_6_delay_19_4 <= io_A_Valid_6_delay_18_5;
    io_A_Valid_6_delay_20_3 <= io_A_Valid_6_delay_19_4;
    io_A_Valid_6_delay_21_2 <= io_A_Valid_6_delay_20_3;
    io_A_Valid_6_delay_22_1 <= io_A_Valid_6_delay_21_2;
    io_A_Valid_6_delay_23 <= io_A_Valid_6_delay_22_1;
    io_B_Valid_23_delay_1_5 <= io_B_Valid_23;
    io_B_Valid_23_delay_2_4 <= io_B_Valid_23_delay_1_5;
    io_B_Valid_23_delay_3_3 <= io_B_Valid_23_delay_2_4;
    io_B_Valid_23_delay_4_2 <= io_B_Valid_23_delay_3_3;
    io_B_Valid_23_delay_5_1 <= io_B_Valid_23_delay_4_2;
    io_B_Valid_23_delay_6 <= io_B_Valid_23_delay_5_1;
    io_A_Valid_6_delay_1_23 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_22 <= io_A_Valid_6_delay_1_23;
    io_A_Valid_6_delay_3_21 <= io_A_Valid_6_delay_2_22;
    io_A_Valid_6_delay_4_20 <= io_A_Valid_6_delay_3_21;
    io_A_Valid_6_delay_5_19 <= io_A_Valid_6_delay_4_20;
    io_A_Valid_6_delay_6_18 <= io_A_Valid_6_delay_5_19;
    io_A_Valid_6_delay_7_17 <= io_A_Valid_6_delay_6_18;
    io_A_Valid_6_delay_8_16 <= io_A_Valid_6_delay_7_17;
    io_A_Valid_6_delay_9_15 <= io_A_Valid_6_delay_8_16;
    io_A_Valid_6_delay_10_14 <= io_A_Valid_6_delay_9_15;
    io_A_Valid_6_delay_11_13 <= io_A_Valid_6_delay_10_14;
    io_A_Valid_6_delay_12_12 <= io_A_Valid_6_delay_11_13;
    io_A_Valid_6_delay_13_11 <= io_A_Valid_6_delay_12_12;
    io_A_Valid_6_delay_14_10 <= io_A_Valid_6_delay_13_11;
    io_A_Valid_6_delay_15_9 <= io_A_Valid_6_delay_14_10;
    io_A_Valid_6_delay_16_8 <= io_A_Valid_6_delay_15_9;
    io_A_Valid_6_delay_17_7 <= io_A_Valid_6_delay_16_8;
    io_A_Valid_6_delay_18_6 <= io_A_Valid_6_delay_17_7;
    io_A_Valid_6_delay_19_5 <= io_A_Valid_6_delay_18_6;
    io_A_Valid_6_delay_20_4 <= io_A_Valid_6_delay_19_5;
    io_A_Valid_6_delay_21_3 <= io_A_Valid_6_delay_20_4;
    io_A_Valid_6_delay_22_2 <= io_A_Valid_6_delay_21_3;
    io_A_Valid_6_delay_23_1 <= io_A_Valid_6_delay_22_2;
    io_A_Valid_6_delay_24 <= io_A_Valid_6_delay_23_1;
    io_B_Valid_24_delay_1_5 <= io_B_Valid_24;
    io_B_Valid_24_delay_2_4 <= io_B_Valid_24_delay_1_5;
    io_B_Valid_24_delay_3_3 <= io_B_Valid_24_delay_2_4;
    io_B_Valid_24_delay_4_2 <= io_B_Valid_24_delay_3_3;
    io_B_Valid_24_delay_5_1 <= io_B_Valid_24_delay_4_2;
    io_B_Valid_24_delay_6 <= io_B_Valid_24_delay_5_1;
    io_A_Valid_6_delay_1_24 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_23 <= io_A_Valid_6_delay_1_24;
    io_A_Valid_6_delay_3_22 <= io_A_Valid_6_delay_2_23;
    io_A_Valid_6_delay_4_21 <= io_A_Valid_6_delay_3_22;
    io_A_Valid_6_delay_5_20 <= io_A_Valid_6_delay_4_21;
    io_A_Valid_6_delay_6_19 <= io_A_Valid_6_delay_5_20;
    io_A_Valid_6_delay_7_18 <= io_A_Valid_6_delay_6_19;
    io_A_Valid_6_delay_8_17 <= io_A_Valid_6_delay_7_18;
    io_A_Valid_6_delay_9_16 <= io_A_Valid_6_delay_8_17;
    io_A_Valid_6_delay_10_15 <= io_A_Valid_6_delay_9_16;
    io_A_Valid_6_delay_11_14 <= io_A_Valid_6_delay_10_15;
    io_A_Valid_6_delay_12_13 <= io_A_Valid_6_delay_11_14;
    io_A_Valid_6_delay_13_12 <= io_A_Valid_6_delay_12_13;
    io_A_Valid_6_delay_14_11 <= io_A_Valid_6_delay_13_12;
    io_A_Valid_6_delay_15_10 <= io_A_Valid_6_delay_14_11;
    io_A_Valid_6_delay_16_9 <= io_A_Valid_6_delay_15_10;
    io_A_Valid_6_delay_17_8 <= io_A_Valid_6_delay_16_9;
    io_A_Valid_6_delay_18_7 <= io_A_Valid_6_delay_17_8;
    io_A_Valid_6_delay_19_6 <= io_A_Valid_6_delay_18_7;
    io_A_Valid_6_delay_20_5 <= io_A_Valid_6_delay_19_6;
    io_A_Valid_6_delay_21_4 <= io_A_Valid_6_delay_20_5;
    io_A_Valid_6_delay_22_3 <= io_A_Valid_6_delay_21_4;
    io_A_Valid_6_delay_23_2 <= io_A_Valid_6_delay_22_3;
    io_A_Valid_6_delay_24_1 <= io_A_Valid_6_delay_23_2;
    io_A_Valid_6_delay_25 <= io_A_Valid_6_delay_24_1;
    io_B_Valid_25_delay_1_5 <= io_B_Valid_25;
    io_B_Valid_25_delay_2_4 <= io_B_Valid_25_delay_1_5;
    io_B_Valid_25_delay_3_3 <= io_B_Valid_25_delay_2_4;
    io_B_Valid_25_delay_4_2 <= io_B_Valid_25_delay_3_3;
    io_B_Valid_25_delay_5_1 <= io_B_Valid_25_delay_4_2;
    io_B_Valid_25_delay_6 <= io_B_Valid_25_delay_5_1;
    io_A_Valid_6_delay_1_25 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_24 <= io_A_Valid_6_delay_1_25;
    io_A_Valid_6_delay_3_23 <= io_A_Valid_6_delay_2_24;
    io_A_Valid_6_delay_4_22 <= io_A_Valid_6_delay_3_23;
    io_A_Valid_6_delay_5_21 <= io_A_Valid_6_delay_4_22;
    io_A_Valid_6_delay_6_20 <= io_A_Valid_6_delay_5_21;
    io_A_Valid_6_delay_7_19 <= io_A_Valid_6_delay_6_20;
    io_A_Valid_6_delay_8_18 <= io_A_Valid_6_delay_7_19;
    io_A_Valid_6_delay_9_17 <= io_A_Valid_6_delay_8_18;
    io_A_Valid_6_delay_10_16 <= io_A_Valid_6_delay_9_17;
    io_A_Valid_6_delay_11_15 <= io_A_Valid_6_delay_10_16;
    io_A_Valid_6_delay_12_14 <= io_A_Valid_6_delay_11_15;
    io_A_Valid_6_delay_13_13 <= io_A_Valid_6_delay_12_14;
    io_A_Valid_6_delay_14_12 <= io_A_Valid_6_delay_13_13;
    io_A_Valid_6_delay_15_11 <= io_A_Valid_6_delay_14_12;
    io_A_Valid_6_delay_16_10 <= io_A_Valid_6_delay_15_11;
    io_A_Valid_6_delay_17_9 <= io_A_Valid_6_delay_16_10;
    io_A_Valid_6_delay_18_8 <= io_A_Valid_6_delay_17_9;
    io_A_Valid_6_delay_19_7 <= io_A_Valid_6_delay_18_8;
    io_A_Valid_6_delay_20_6 <= io_A_Valid_6_delay_19_7;
    io_A_Valid_6_delay_21_5 <= io_A_Valid_6_delay_20_6;
    io_A_Valid_6_delay_22_4 <= io_A_Valid_6_delay_21_5;
    io_A_Valid_6_delay_23_3 <= io_A_Valid_6_delay_22_4;
    io_A_Valid_6_delay_24_2 <= io_A_Valid_6_delay_23_3;
    io_A_Valid_6_delay_25_1 <= io_A_Valid_6_delay_24_2;
    io_A_Valid_6_delay_26 <= io_A_Valid_6_delay_25_1;
    io_B_Valid_26_delay_1_5 <= io_B_Valid_26;
    io_B_Valid_26_delay_2_4 <= io_B_Valid_26_delay_1_5;
    io_B_Valid_26_delay_3_3 <= io_B_Valid_26_delay_2_4;
    io_B_Valid_26_delay_4_2 <= io_B_Valid_26_delay_3_3;
    io_B_Valid_26_delay_5_1 <= io_B_Valid_26_delay_4_2;
    io_B_Valid_26_delay_6 <= io_B_Valid_26_delay_5_1;
    io_A_Valid_6_delay_1_26 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_25 <= io_A_Valid_6_delay_1_26;
    io_A_Valid_6_delay_3_24 <= io_A_Valid_6_delay_2_25;
    io_A_Valid_6_delay_4_23 <= io_A_Valid_6_delay_3_24;
    io_A_Valid_6_delay_5_22 <= io_A_Valid_6_delay_4_23;
    io_A_Valid_6_delay_6_21 <= io_A_Valid_6_delay_5_22;
    io_A_Valid_6_delay_7_20 <= io_A_Valid_6_delay_6_21;
    io_A_Valid_6_delay_8_19 <= io_A_Valid_6_delay_7_20;
    io_A_Valid_6_delay_9_18 <= io_A_Valid_6_delay_8_19;
    io_A_Valid_6_delay_10_17 <= io_A_Valid_6_delay_9_18;
    io_A_Valid_6_delay_11_16 <= io_A_Valid_6_delay_10_17;
    io_A_Valid_6_delay_12_15 <= io_A_Valid_6_delay_11_16;
    io_A_Valid_6_delay_13_14 <= io_A_Valid_6_delay_12_15;
    io_A_Valid_6_delay_14_13 <= io_A_Valid_6_delay_13_14;
    io_A_Valid_6_delay_15_12 <= io_A_Valid_6_delay_14_13;
    io_A_Valid_6_delay_16_11 <= io_A_Valid_6_delay_15_12;
    io_A_Valid_6_delay_17_10 <= io_A_Valid_6_delay_16_11;
    io_A_Valid_6_delay_18_9 <= io_A_Valid_6_delay_17_10;
    io_A_Valid_6_delay_19_8 <= io_A_Valid_6_delay_18_9;
    io_A_Valid_6_delay_20_7 <= io_A_Valid_6_delay_19_8;
    io_A_Valid_6_delay_21_6 <= io_A_Valid_6_delay_20_7;
    io_A_Valid_6_delay_22_5 <= io_A_Valid_6_delay_21_6;
    io_A_Valid_6_delay_23_4 <= io_A_Valid_6_delay_22_5;
    io_A_Valid_6_delay_24_3 <= io_A_Valid_6_delay_23_4;
    io_A_Valid_6_delay_25_2 <= io_A_Valid_6_delay_24_3;
    io_A_Valid_6_delay_26_1 <= io_A_Valid_6_delay_25_2;
    io_A_Valid_6_delay_27 <= io_A_Valid_6_delay_26_1;
    io_B_Valid_27_delay_1_5 <= io_B_Valid_27;
    io_B_Valid_27_delay_2_4 <= io_B_Valid_27_delay_1_5;
    io_B_Valid_27_delay_3_3 <= io_B_Valid_27_delay_2_4;
    io_B_Valid_27_delay_4_2 <= io_B_Valid_27_delay_3_3;
    io_B_Valid_27_delay_5_1 <= io_B_Valid_27_delay_4_2;
    io_B_Valid_27_delay_6 <= io_B_Valid_27_delay_5_1;
    io_A_Valid_6_delay_1_27 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_26 <= io_A_Valid_6_delay_1_27;
    io_A_Valid_6_delay_3_25 <= io_A_Valid_6_delay_2_26;
    io_A_Valid_6_delay_4_24 <= io_A_Valid_6_delay_3_25;
    io_A_Valid_6_delay_5_23 <= io_A_Valid_6_delay_4_24;
    io_A_Valid_6_delay_6_22 <= io_A_Valid_6_delay_5_23;
    io_A_Valid_6_delay_7_21 <= io_A_Valid_6_delay_6_22;
    io_A_Valid_6_delay_8_20 <= io_A_Valid_6_delay_7_21;
    io_A_Valid_6_delay_9_19 <= io_A_Valid_6_delay_8_20;
    io_A_Valid_6_delay_10_18 <= io_A_Valid_6_delay_9_19;
    io_A_Valid_6_delay_11_17 <= io_A_Valid_6_delay_10_18;
    io_A_Valid_6_delay_12_16 <= io_A_Valid_6_delay_11_17;
    io_A_Valid_6_delay_13_15 <= io_A_Valid_6_delay_12_16;
    io_A_Valid_6_delay_14_14 <= io_A_Valid_6_delay_13_15;
    io_A_Valid_6_delay_15_13 <= io_A_Valid_6_delay_14_14;
    io_A_Valid_6_delay_16_12 <= io_A_Valid_6_delay_15_13;
    io_A_Valid_6_delay_17_11 <= io_A_Valid_6_delay_16_12;
    io_A_Valid_6_delay_18_10 <= io_A_Valid_6_delay_17_11;
    io_A_Valid_6_delay_19_9 <= io_A_Valid_6_delay_18_10;
    io_A_Valid_6_delay_20_8 <= io_A_Valid_6_delay_19_9;
    io_A_Valid_6_delay_21_7 <= io_A_Valid_6_delay_20_8;
    io_A_Valid_6_delay_22_6 <= io_A_Valid_6_delay_21_7;
    io_A_Valid_6_delay_23_5 <= io_A_Valid_6_delay_22_6;
    io_A_Valid_6_delay_24_4 <= io_A_Valid_6_delay_23_5;
    io_A_Valid_6_delay_25_3 <= io_A_Valid_6_delay_24_4;
    io_A_Valid_6_delay_26_2 <= io_A_Valid_6_delay_25_3;
    io_A_Valid_6_delay_27_1 <= io_A_Valid_6_delay_26_2;
    io_A_Valid_6_delay_28 <= io_A_Valid_6_delay_27_1;
    io_B_Valid_28_delay_1_5 <= io_B_Valid_28;
    io_B_Valid_28_delay_2_4 <= io_B_Valid_28_delay_1_5;
    io_B_Valid_28_delay_3_3 <= io_B_Valid_28_delay_2_4;
    io_B_Valid_28_delay_4_2 <= io_B_Valid_28_delay_3_3;
    io_B_Valid_28_delay_5_1 <= io_B_Valid_28_delay_4_2;
    io_B_Valid_28_delay_6 <= io_B_Valid_28_delay_5_1;
    io_A_Valid_6_delay_1_28 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_27 <= io_A_Valid_6_delay_1_28;
    io_A_Valid_6_delay_3_26 <= io_A_Valid_6_delay_2_27;
    io_A_Valid_6_delay_4_25 <= io_A_Valid_6_delay_3_26;
    io_A_Valid_6_delay_5_24 <= io_A_Valid_6_delay_4_25;
    io_A_Valid_6_delay_6_23 <= io_A_Valid_6_delay_5_24;
    io_A_Valid_6_delay_7_22 <= io_A_Valid_6_delay_6_23;
    io_A_Valid_6_delay_8_21 <= io_A_Valid_6_delay_7_22;
    io_A_Valid_6_delay_9_20 <= io_A_Valid_6_delay_8_21;
    io_A_Valid_6_delay_10_19 <= io_A_Valid_6_delay_9_20;
    io_A_Valid_6_delay_11_18 <= io_A_Valid_6_delay_10_19;
    io_A_Valid_6_delay_12_17 <= io_A_Valid_6_delay_11_18;
    io_A_Valid_6_delay_13_16 <= io_A_Valid_6_delay_12_17;
    io_A_Valid_6_delay_14_15 <= io_A_Valid_6_delay_13_16;
    io_A_Valid_6_delay_15_14 <= io_A_Valid_6_delay_14_15;
    io_A_Valid_6_delay_16_13 <= io_A_Valid_6_delay_15_14;
    io_A_Valid_6_delay_17_12 <= io_A_Valid_6_delay_16_13;
    io_A_Valid_6_delay_18_11 <= io_A_Valid_6_delay_17_12;
    io_A_Valid_6_delay_19_10 <= io_A_Valid_6_delay_18_11;
    io_A_Valid_6_delay_20_9 <= io_A_Valid_6_delay_19_10;
    io_A_Valid_6_delay_21_8 <= io_A_Valid_6_delay_20_9;
    io_A_Valid_6_delay_22_7 <= io_A_Valid_6_delay_21_8;
    io_A_Valid_6_delay_23_6 <= io_A_Valid_6_delay_22_7;
    io_A_Valid_6_delay_24_5 <= io_A_Valid_6_delay_23_6;
    io_A_Valid_6_delay_25_4 <= io_A_Valid_6_delay_24_5;
    io_A_Valid_6_delay_26_3 <= io_A_Valid_6_delay_25_4;
    io_A_Valid_6_delay_27_2 <= io_A_Valid_6_delay_26_3;
    io_A_Valid_6_delay_28_1 <= io_A_Valid_6_delay_27_2;
    io_A_Valid_6_delay_29 <= io_A_Valid_6_delay_28_1;
    io_B_Valid_29_delay_1_5 <= io_B_Valid_29;
    io_B_Valid_29_delay_2_4 <= io_B_Valid_29_delay_1_5;
    io_B_Valid_29_delay_3_3 <= io_B_Valid_29_delay_2_4;
    io_B_Valid_29_delay_4_2 <= io_B_Valid_29_delay_3_3;
    io_B_Valid_29_delay_5_1 <= io_B_Valid_29_delay_4_2;
    io_B_Valid_29_delay_6 <= io_B_Valid_29_delay_5_1;
    io_A_Valid_6_delay_1_29 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_28 <= io_A_Valid_6_delay_1_29;
    io_A_Valid_6_delay_3_27 <= io_A_Valid_6_delay_2_28;
    io_A_Valid_6_delay_4_26 <= io_A_Valid_6_delay_3_27;
    io_A_Valid_6_delay_5_25 <= io_A_Valid_6_delay_4_26;
    io_A_Valid_6_delay_6_24 <= io_A_Valid_6_delay_5_25;
    io_A_Valid_6_delay_7_23 <= io_A_Valid_6_delay_6_24;
    io_A_Valid_6_delay_8_22 <= io_A_Valid_6_delay_7_23;
    io_A_Valid_6_delay_9_21 <= io_A_Valid_6_delay_8_22;
    io_A_Valid_6_delay_10_20 <= io_A_Valid_6_delay_9_21;
    io_A_Valid_6_delay_11_19 <= io_A_Valid_6_delay_10_20;
    io_A_Valid_6_delay_12_18 <= io_A_Valid_6_delay_11_19;
    io_A_Valid_6_delay_13_17 <= io_A_Valid_6_delay_12_18;
    io_A_Valid_6_delay_14_16 <= io_A_Valid_6_delay_13_17;
    io_A_Valid_6_delay_15_15 <= io_A_Valid_6_delay_14_16;
    io_A_Valid_6_delay_16_14 <= io_A_Valid_6_delay_15_15;
    io_A_Valid_6_delay_17_13 <= io_A_Valid_6_delay_16_14;
    io_A_Valid_6_delay_18_12 <= io_A_Valid_6_delay_17_13;
    io_A_Valid_6_delay_19_11 <= io_A_Valid_6_delay_18_12;
    io_A_Valid_6_delay_20_10 <= io_A_Valid_6_delay_19_11;
    io_A_Valid_6_delay_21_9 <= io_A_Valid_6_delay_20_10;
    io_A_Valid_6_delay_22_8 <= io_A_Valid_6_delay_21_9;
    io_A_Valid_6_delay_23_7 <= io_A_Valid_6_delay_22_8;
    io_A_Valid_6_delay_24_6 <= io_A_Valid_6_delay_23_7;
    io_A_Valid_6_delay_25_5 <= io_A_Valid_6_delay_24_6;
    io_A_Valid_6_delay_26_4 <= io_A_Valid_6_delay_25_5;
    io_A_Valid_6_delay_27_3 <= io_A_Valid_6_delay_26_4;
    io_A_Valid_6_delay_28_2 <= io_A_Valid_6_delay_27_3;
    io_A_Valid_6_delay_29_1 <= io_A_Valid_6_delay_28_2;
    io_A_Valid_6_delay_30 <= io_A_Valid_6_delay_29_1;
    io_B_Valid_30_delay_1_5 <= io_B_Valid_30;
    io_B_Valid_30_delay_2_4 <= io_B_Valid_30_delay_1_5;
    io_B_Valid_30_delay_3_3 <= io_B_Valid_30_delay_2_4;
    io_B_Valid_30_delay_4_2 <= io_B_Valid_30_delay_3_3;
    io_B_Valid_30_delay_5_1 <= io_B_Valid_30_delay_4_2;
    io_B_Valid_30_delay_6 <= io_B_Valid_30_delay_5_1;
    io_A_Valid_6_delay_1_30 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_29 <= io_A_Valid_6_delay_1_30;
    io_A_Valid_6_delay_3_28 <= io_A_Valid_6_delay_2_29;
    io_A_Valid_6_delay_4_27 <= io_A_Valid_6_delay_3_28;
    io_A_Valid_6_delay_5_26 <= io_A_Valid_6_delay_4_27;
    io_A_Valid_6_delay_6_25 <= io_A_Valid_6_delay_5_26;
    io_A_Valid_6_delay_7_24 <= io_A_Valid_6_delay_6_25;
    io_A_Valid_6_delay_8_23 <= io_A_Valid_6_delay_7_24;
    io_A_Valid_6_delay_9_22 <= io_A_Valid_6_delay_8_23;
    io_A_Valid_6_delay_10_21 <= io_A_Valid_6_delay_9_22;
    io_A_Valid_6_delay_11_20 <= io_A_Valid_6_delay_10_21;
    io_A_Valid_6_delay_12_19 <= io_A_Valid_6_delay_11_20;
    io_A_Valid_6_delay_13_18 <= io_A_Valid_6_delay_12_19;
    io_A_Valid_6_delay_14_17 <= io_A_Valid_6_delay_13_18;
    io_A_Valid_6_delay_15_16 <= io_A_Valid_6_delay_14_17;
    io_A_Valid_6_delay_16_15 <= io_A_Valid_6_delay_15_16;
    io_A_Valid_6_delay_17_14 <= io_A_Valid_6_delay_16_15;
    io_A_Valid_6_delay_18_13 <= io_A_Valid_6_delay_17_14;
    io_A_Valid_6_delay_19_12 <= io_A_Valid_6_delay_18_13;
    io_A_Valid_6_delay_20_11 <= io_A_Valid_6_delay_19_12;
    io_A_Valid_6_delay_21_10 <= io_A_Valid_6_delay_20_11;
    io_A_Valid_6_delay_22_9 <= io_A_Valid_6_delay_21_10;
    io_A_Valid_6_delay_23_8 <= io_A_Valid_6_delay_22_9;
    io_A_Valid_6_delay_24_7 <= io_A_Valid_6_delay_23_8;
    io_A_Valid_6_delay_25_6 <= io_A_Valid_6_delay_24_7;
    io_A_Valid_6_delay_26_5 <= io_A_Valid_6_delay_25_6;
    io_A_Valid_6_delay_27_4 <= io_A_Valid_6_delay_26_5;
    io_A_Valid_6_delay_28_3 <= io_A_Valid_6_delay_27_4;
    io_A_Valid_6_delay_29_2 <= io_A_Valid_6_delay_28_3;
    io_A_Valid_6_delay_30_1 <= io_A_Valid_6_delay_29_2;
    io_A_Valid_6_delay_31 <= io_A_Valid_6_delay_30_1;
    io_B_Valid_31_delay_1_5 <= io_B_Valid_31;
    io_B_Valid_31_delay_2_4 <= io_B_Valid_31_delay_1_5;
    io_B_Valid_31_delay_3_3 <= io_B_Valid_31_delay_2_4;
    io_B_Valid_31_delay_4_2 <= io_B_Valid_31_delay_3_3;
    io_B_Valid_31_delay_5_1 <= io_B_Valid_31_delay_4_2;
    io_B_Valid_31_delay_6 <= io_B_Valid_31_delay_5_1;
    io_A_Valid_6_delay_1_31 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_30 <= io_A_Valid_6_delay_1_31;
    io_A_Valid_6_delay_3_29 <= io_A_Valid_6_delay_2_30;
    io_A_Valid_6_delay_4_28 <= io_A_Valid_6_delay_3_29;
    io_A_Valid_6_delay_5_27 <= io_A_Valid_6_delay_4_28;
    io_A_Valid_6_delay_6_26 <= io_A_Valid_6_delay_5_27;
    io_A_Valid_6_delay_7_25 <= io_A_Valid_6_delay_6_26;
    io_A_Valid_6_delay_8_24 <= io_A_Valid_6_delay_7_25;
    io_A_Valid_6_delay_9_23 <= io_A_Valid_6_delay_8_24;
    io_A_Valid_6_delay_10_22 <= io_A_Valid_6_delay_9_23;
    io_A_Valid_6_delay_11_21 <= io_A_Valid_6_delay_10_22;
    io_A_Valid_6_delay_12_20 <= io_A_Valid_6_delay_11_21;
    io_A_Valid_6_delay_13_19 <= io_A_Valid_6_delay_12_20;
    io_A_Valid_6_delay_14_18 <= io_A_Valid_6_delay_13_19;
    io_A_Valid_6_delay_15_17 <= io_A_Valid_6_delay_14_18;
    io_A_Valid_6_delay_16_16 <= io_A_Valid_6_delay_15_17;
    io_A_Valid_6_delay_17_15 <= io_A_Valid_6_delay_16_16;
    io_A_Valid_6_delay_18_14 <= io_A_Valid_6_delay_17_15;
    io_A_Valid_6_delay_19_13 <= io_A_Valid_6_delay_18_14;
    io_A_Valid_6_delay_20_12 <= io_A_Valid_6_delay_19_13;
    io_A_Valid_6_delay_21_11 <= io_A_Valid_6_delay_20_12;
    io_A_Valid_6_delay_22_10 <= io_A_Valid_6_delay_21_11;
    io_A_Valid_6_delay_23_9 <= io_A_Valid_6_delay_22_10;
    io_A_Valid_6_delay_24_8 <= io_A_Valid_6_delay_23_9;
    io_A_Valid_6_delay_25_7 <= io_A_Valid_6_delay_24_8;
    io_A_Valid_6_delay_26_6 <= io_A_Valid_6_delay_25_7;
    io_A_Valid_6_delay_27_5 <= io_A_Valid_6_delay_26_6;
    io_A_Valid_6_delay_28_4 <= io_A_Valid_6_delay_27_5;
    io_A_Valid_6_delay_29_3 <= io_A_Valid_6_delay_28_4;
    io_A_Valid_6_delay_30_2 <= io_A_Valid_6_delay_29_3;
    io_A_Valid_6_delay_31_1 <= io_A_Valid_6_delay_30_2;
    io_A_Valid_6_delay_32 <= io_A_Valid_6_delay_31_1;
    io_B_Valid_32_delay_1_5 <= io_B_Valid_32;
    io_B_Valid_32_delay_2_4 <= io_B_Valid_32_delay_1_5;
    io_B_Valid_32_delay_3_3 <= io_B_Valid_32_delay_2_4;
    io_B_Valid_32_delay_4_2 <= io_B_Valid_32_delay_3_3;
    io_B_Valid_32_delay_5_1 <= io_B_Valid_32_delay_4_2;
    io_B_Valid_32_delay_6 <= io_B_Valid_32_delay_5_1;
    io_A_Valid_6_delay_1_32 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_31 <= io_A_Valid_6_delay_1_32;
    io_A_Valid_6_delay_3_30 <= io_A_Valid_6_delay_2_31;
    io_A_Valid_6_delay_4_29 <= io_A_Valid_6_delay_3_30;
    io_A_Valid_6_delay_5_28 <= io_A_Valid_6_delay_4_29;
    io_A_Valid_6_delay_6_27 <= io_A_Valid_6_delay_5_28;
    io_A_Valid_6_delay_7_26 <= io_A_Valid_6_delay_6_27;
    io_A_Valid_6_delay_8_25 <= io_A_Valid_6_delay_7_26;
    io_A_Valid_6_delay_9_24 <= io_A_Valid_6_delay_8_25;
    io_A_Valid_6_delay_10_23 <= io_A_Valid_6_delay_9_24;
    io_A_Valid_6_delay_11_22 <= io_A_Valid_6_delay_10_23;
    io_A_Valid_6_delay_12_21 <= io_A_Valid_6_delay_11_22;
    io_A_Valid_6_delay_13_20 <= io_A_Valid_6_delay_12_21;
    io_A_Valid_6_delay_14_19 <= io_A_Valid_6_delay_13_20;
    io_A_Valid_6_delay_15_18 <= io_A_Valid_6_delay_14_19;
    io_A_Valid_6_delay_16_17 <= io_A_Valid_6_delay_15_18;
    io_A_Valid_6_delay_17_16 <= io_A_Valid_6_delay_16_17;
    io_A_Valid_6_delay_18_15 <= io_A_Valid_6_delay_17_16;
    io_A_Valid_6_delay_19_14 <= io_A_Valid_6_delay_18_15;
    io_A_Valid_6_delay_20_13 <= io_A_Valid_6_delay_19_14;
    io_A_Valid_6_delay_21_12 <= io_A_Valid_6_delay_20_13;
    io_A_Valid_6_delay_22_11 <= io_A_Valid_6_delay_21_12;
    io_A_Valid_6_delay_23_10 <= io_A_Valid_6_delay_22_11;
    io_A_Valid_6_delay_24_9 <= io_A_Valid_6_delay_23_10;
    io_A_Valid_6_delay_25_8 <= io_A_Valid_6_delay_24_9;
    io_A_Valid_6_delay_26_7 <= io_A_Valid_6_delay_25_8;
    io_A_Valid_6_delay_27_6 <= io_A_Valid_6_delay_26_7;
    io_A_Valid_6_delay_28_5 <= io_A_Valid_6_delay_27_6;
    io_A_Valid_6_delay_29_4 <= io_A_Valid_6_delay_28_5;
    io_A_Valid_6_delay_30_3 <= io_A_Valid_6_delay_29_4;
    io_A_Valid_6_delay_31_2 <= io_A_Valid_6_delay_30_3;
    io_A_Valid_6_delay_32_1 <= io_A_Valid_6_delay_31_2;
    io_A_Valid_6_delay_33 <= io_A_Valid_6_delay_32_1;
    io_B_Valid_33_delay_1_5 <= io_B_Valid_33;
    io_B_Valid_33_delay_2_4 <= io_B_Valid_33_delay_1_5;
    io_B_Valid_33_delay_3_3 <= io_B_Valid_33_delay_2_4;
    io_B_Valid_33_delay_4_2 <= io_B_Valid_33_delay_3_3;
    io_B_Valid_33_delay_5_1 <= io_B_Valid_33_delay_4_2;
    io_B_Valid_33_delay_6 <= io_B_Valid_33_delay_5_1;
    io_A_Valid_6_delay_1_33 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_32 <= io_A_Valid_6_delay_1_33;
    io_A_Valid_6_delay_3_31 <= io_A_Valid_6_delay_2_32;
    io_A_Valid_6_delay_4_30 <= io_A_Valid_6_delay_3_31;
    io_A_Valid_6_delay_5_29 <= io_A_Valid_6_delay_4_30;
    io_A_Valid_6_delay_6_28 <= io_A_Valid_6_delay_5_29;
    io_A_Valid_6_delay_7_27 <= io_A_Valid_6_delay_6_28;
    io_A_Valid_6_delay_8_26 <= io_A_Valid_6_delay_7_27;
    io_A_Valid_6_delay_9_25 <= io_A_Valid_6_delay_8_26;
    io_A_Valid_6_delay_10_24 <= io_A_Valid_6_delay_9_25;
    io_A_Valid_6_delay_11_23 <= io_A_Valid_6_delay_10_24;
    io_A_Valid_6_delay_12_22 <= io_A_Valid_6_delay_11_23;
    io_A_Valid_6_delay_13_21 <= io_A_Valid_6_delay_12_22;
    io_A_Valid_6_delay_14_20 <= io_A_Valid_6_delay_13_21;
    io_A_Valid_6_delay_15_19 <= io_A_Valid_6_delay_14_20;
    io_A_Valid_6_delay_16_18 <= io_A_Valid_6_delay_15_19;
    io_A_Valid_6_delay_17_17 <= io_A_Valid_6_delay_16_18;
    io_A_Valid_6_delay_18_16 <= io_A_Valid_6_delay_17_17;
    io_A_Valid_6_delay_19_15 <= io_A_Valid_6_delay_18_16;
    io_A_Valid_6_delay_20_14 <= io_A_Valid_6_delay_19_15;
    io_A_Valid_6_delay_21_13 <= io_A_Valid_6_delay_20_14;
    io_A_Valid_6_delay_22_12 <= io_A_Valid_6_delay_21_13;
    io_A_Valid_6_delay_23_11 <= io_A_Valid_6_delay_22_12;
    io_A_Valid_6_delay_24_10 <= io_A_Valid_6_delay_23_11;
    io_A_Valid_6_delay_25_9 <= io_A_Valid_6_delay_24_10;
    io_A_Valid_6_delay_26_8 <= io_A_Valid_6_delay_25_9;
    io_A_Valid_6_delay_27_7 <= io_A_Valid_6_delay_26_8;
    io_A_Valid_6_delay_28_6 <= io_A_Valid_6_delay_27_7;
    io_A_Valid_6_delay_29_5 <= io_A_Valid_6_delay_28_6;
    io_A_Valid_6_delay_30_4 <= io_A_Valid_6_delay_29_5;
    io_A_Valid_6_delay_31_3 <= io_A_Valid_6_delay_30_4;
    io_A_Valid_6_delay_32_2 <= io_A_Valid_6_delay_31_3;
    io_A_Valid_6_delay_33_1 <= io_A_Valid_6_delay_32_2;
    io_A_Valid_6_delay_34 <= io_A_Valid_6_delay_33_1;
    io_B_Valid_34_delay_1_5 <= io_B_Valid_34;
    io_B_Valid_34_delay_2_4 <= io_B_Valid_34_delay_1_5;
    io_B_Valid_34_delay_3_3 <= io_B_Valid_34_delay_2_4;
    io_B_Valid_34_delay_4_2 <= io_B_Valid_34_delay_3_3;
    io_B_Valid_34_delay_5_1 <= io_B_Valid_34_delay_4_2;
    io_B_Valid_34_delay_6 <= io_B_Valid_34_delay_5_1;
    io_A_Valid_6_delay_1_34 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_33 <= io_A_Valid_6_delay_1_34;
    io_A_Valid_6_delay_3_32 <= io_A_Valid_6_delay_2_33;
    io_A_Valid_6_delay_4_31 <= io_A_Valid_6_delay_3_32;
    io_A_Valid_6_delay_5_30 <= io_A_Valid_6_delay_4_31;
    io_A_Valid_6_delay_6_29 <= io_A_Valid_6_delay_5_30;
    io_A_Valid_6_delay_7_28 <= io_A_Valid_6_delay_6_29;
    io_A_Valid_6_delay_8_27 <= io_A_Valid_6_delay_7_28;
    io_A_Valid_6_delay_9_26 <= io_A_Valid_6_delay_8_27;
    io_A_Valid_6_delay_10_25 <= io_A_Valid_6_delay_9_26;
    io_A_Valid_6_delay_11_24 <= io_A_Valid_6_delay_10_25;
    io_A_Valid_6_delay_12_23 <= io_A_Valid_6_delay_11_24;
    io_A_Valid_6_delay_13_22 <= io_A_Valid_6_delay_12_23;
    io_A_Valid_6_delay_14_21 <= io_A_Valid_6_delay_13_22;
    io_A_Valid_6_delay_15_20 <= io_A_Valid_6_delay_14_21;
    io_A_Valid_6_delay_16_19 <= io_A_Valid_6_delay_15_20;
    io_A_Valid_6_delay_17_18 <= io_A_Valid_6_delay_16_19;
    io_A_Valid_6_delay_18_17 <= io_A_Valid_6_delay_17_18;
    io_A_Valid_6_delay_19_16 <= io_A_Valid_6_delay_18_17;
    io_A_Valid_6_delay_20_15 <= io_A_Valid_6_delay_19_16;
    io_A_Valid_6_delay_21_14 <= io_A_Valid_6_delay_20_15;
    io_A_Valid_6_delay_22_13 <= io_A_Valid_6_delay_21_14;
    io_A_Valid_6_delay_23_12 <= io_A_Valid_6_delay_22_13;
    io_A_Valid_6_delay_24_11 <= io_A_Valid_6_delay_23_12;
    io_A_Valid_6_delay_25_10 <= io_A_Valid_6_delay_24_11;
    io_A_Valid_6_delay_26_9 <= io_A_Valid_6_delay_25_10;
    io_A_Valid_6_delay_27_8 <= io_A_Valid_6_delay_26_9;
    io_A_Valid_6_delay_28_7 <= io_A_Valid_6_delay_27_8;
    io_A_Valid_6_delay_29_6 <= io_A_Valid_6_delay_28_7;
    io_A_Valid_6_delay_30_5 <= io_A_Valid_6_delay_29_6;
    io_A_Valid_6_delay_31_4 <= io_A_Valid_6_delay_30_5;
    io_A_Valid_6_delay_32_3 <= io_A_Valid_6_delay_31_4;
    io_A_Valid_6_delay_33_2 <= io_A_Valid_6_delay_32_3;
    io_A_Valid_6_delay_34_1 <= io_A_Valid_6_delay_33_2;
    io_A_Valid_6_delay_35 <= io_A_Valid_6_delay_34_1;
    io_B_Valid_35_delay_1_5 <= io_B_Valid_35;
    io_B_Valid_35_delay_2_4 <= io_B_Valid_35_delay_1_5;
    io_B_Valid_35_delay_3_3 <= io_B_Valid_35_delay_2_4;
    io_B_Valid_35_delay_4_2 <= io_B_Valid_35_delay_3_3;
    io_B_Valid_35_delay_5_1 <= io_B_Valid_35_delay_4_2;
    io_B_Valid_35_delay_6 <= io_B_Valid_35_delay_5_1;
    io_A_Valid_6_delay_1_35 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_34 <= io_A_Valid_6_delay_1_35;
    io_A_Valid_6_delay_3_33 <= io_A_Valid_6_delay_2_34;
    io_A_Valid_6_delay_4_32 <= io_A_Valid_6_delay_3_33;
    io_A_Valid_6_delay_5_31 <= io_A_Valid_6_delay_4_32;
    io_A_Valid_6_delay_6_30 <= io_A_Valid_6_delay_5_31;
    io_A_Valid_6_delay_7_29 <= io_A_Valid_6_delay_6_30;
    io_A_Valid_6_delay_8_28 <= io_A_Valid_6_delay_7_29;
    io_A_Valid_6_delay_9_27 <= io_A_Valid_6_delay_8_28;
    io_A_Valid_6_delay_10_26 <= io_A_Valid_6_delay_9_27;
    io_A_Valid_6_delay_11_25 <= io_A_Valid_6_delay_10_26;
    io_A_Valid_6_delay_12_24 <= io_A_Valid_6_delay_11_25;
    io_A_Valid_6_delay_13_23 <= io_A_Valid_6_delay_12_24;
    io_A_Valid_6_delay_14_22 <= io_A_Valid_6_delay_13_23;
    io_A_Valid_6_delay_15_21 <= io_A_Valid_6_delay_14_22;
    io_A_Valid_6_delay_16_20 <= io_A_Valid_6_delay_15_21;
    io_A_Valid_6_delay_17_19 <= io_A_Valid_6_delay_16_20;
    io_A_Valid_6_delay_18_18 <= io_A_Valid_6_delay_17_19;
    io_A_Valid_6_delay_19_17 <= io_A_Valid_6_delay_18_18;
    io_A_Valid_6_delay_20_16 <= io_A_Valid_6_delay_19_17;
    io_A_Valid_6_delay_21_15 <= io_A_Valid_6_delay_20_16;
    io_A_Valid_6_delay_22_14 <= io_A_Valid_6_delay_21_15;
    io_A_Valid_6_delay_23_13 <= io_A_Valid_6_delay_22_14;
    io_A_Valid_6_delay_24_12 <= io_A_Valid_6_delay_23_13;
    io_A_Valid_6_delay_25_11 <= io_A_Valid_6_delay_24_12;
    io_A_Valid_6_delay_26_10 <= io_A_Valid_6_delay_25_11;
    io_A_Valid_6_delay_27_9 <= io_A_Valid_6_delay_26_10;
    io_A_Valid_6_delay_28_8 <= io_A_Valid_6_delay_27_9;
    io_A_Valid_6_delay_29_7 <= io_A_Valid_6_delay_28_8;
    io_A_Valid_6_delay_30_6 <= io_A_Valid_6_delay_29_7;
    io_A_Valid_6_delay_31_5 <= io_A_Valid_6_delay_30_6;
    io_A_Valid_6_delay_32_4 <= io_A_Valid_6_delay_31_5;
    io_A_Valid_6_delay_33_3 <= io_A_Valid_6_delay_32_4;
    io_A_Valid_6_delay_34_2 <= io_A_Valid_6_delay_33_3;
    io_A_Valid_6_delay_35_1 <= io_A_Valid_6_delay_34_2;
    io_A_Valid_6_delay_36 <= io_A_Valid_6_delay_35_1;
    io_B_Valid_36_delay_1_5 <= io_B_Valid_36;
    io_B_Valid_36_delay_2_4 <= io_B_Valid_36_delay_1_5;
    io_B_Valid_36_delay_3_3 <= io_B_Valid_36_delay_2_4;
    io_B_Valid_36_delay_4_2 <= io_B_Valid_36_delay_3_3;
    io_B_Valid_36_delay_5_1 <= io_B_Valid_36_delay_4_2;
    io_B_Valid_36_delay_6 <= io_B_Valid_36_delay_5_1;
    io_A_Valid_6_delay_1_36 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_35 <= io_A_Valid_6_delay_1_36;
    io_A_Valid_6_delay_3_34 <= io_A_Valid_6_delay_2_35;
    io_A_Valid_6_delay_4_33 <= io_A_Valid_6_delay_3_34;
    io_A_Valid_6_delay_5_32 <= io_A_Valid_6_delay_4_33;
    io_A_Valid_6_delay_6_31 <= io_A_Valid_6_delay_5_32;
    io_A_Valid_6_delay_7_30 <= io_A_Valid_6_delay_6_31;
    io_A_Valid_6_delay_8_29 <= io_A_Valid_6_delay_7_30;
    io_A_Valid_6_delay_9_28 <= io_A_Valid_6_delay_8_29;
    io_A_Valid_6_delay_10_27 <= io_A_Valid_6_delay_9_28;
    io_A_Valid_6_delay_11_26 <= io_A_Valid_6_delay_10_27;
    io_A_Valid_6_delay_12_25 <= io_A_Valid_6_delay_11_26;
    io_A_Valid_6_delay_13_24 <= io_A_Valid_6_delay_12_25;
    io_A_Valid_6_delay_14_23 <= io_A_Valid_6_delay_13_24;
    io_A_Valid_6_delay_15_22 <= io_A_Valid_6_delay_14_23;
    io_A_Valid_6_delay_16_21 <= io_A_Valid_6_delay_15_22;
    io_A_Valid_6_delay_17_20 <= io_A_Valid_6_delay_16_21;
    io_A_Valid_6_delay_18_19 <= io_A_Valid_6_delay_17_20;
    io_A_Valid_6_delay_19_18 <= io_A_Valid_6_delay_18_19;
    io_A_Valid_6_delay_20_17 <= io_A_Valid_6_delay_19_18;
    io_A_Valid_6_delay_21_16 <= io_A_Valid_6_delay_20_17;
    io_A_Valid_6_delay_22_15 <= io_A_Valid_6_delay_21_16;
    io_A_Valid_6_delay_23_14 <= io_A_Valid_6_delay_22_15;
    io_A_Valid_6_delay_24_13 <= io_A_Valid_6_delay_23_14;
    io_A_Valid_6_delay_25_12 <= io_A_Valid_6_delay_24_13;
    io_A_Valid_6_delay_26_11 <= io_A_Valid_6_delay_25_12;
    io_A_Valid_6_delay_27_10 <= io_A_Valid_6_delay_26_11;
    io_A_Valid_6_delay_28_9 <= io_A_Valid_6_delay_27_10;
    io_A_Valid_6_delay_29_8 <= io_A_Valid_6_delay_28_9;
    io_A_Valid_6_delay_30_7 <= io_A_Valid_6_delay_29_8;
    io_A_Valid_6_delay_31_6 <= io_A_Valid_6_delay_30_7;
    io_A_Valid_6_delay_32_5 <= io_A_Valid_6_delay_31_6;
    io_A_Valid_6_delay_33_4 <= io_A_Valid_6_delay_32_5;
    io_A_Valid_6_delay_34_3 <= io_A_Valid_6_delay_33_4;
    io_A_Valid_6_delay_35_2 <= io_A_Valid_6_delay_34_3;
    io_A_Valid_6_delay_36_1 <= io_A_Valid_6_delay_35_2;
    io_A_Valid_6_delay_37 <= io_A_Valid_6_delay_36_1;
    io_B_Valid_37_delay_1_5 <= io_B_Valid_37;
    io_B_Valid_37_delay_2_4 <= io_B_Valid_37_delay_1_5;
    io_B_Valid_37_delay_3_3 <= io_B_Valid_37_delay_2_4;
    io_B_Valid_37_delay_4_2 <= io_B_Valid_37_delay_3_3;
    io_B_Valid_37_delay_5_1 <= io_B_Valid_37_delay_4_2;
    io_B_Valid_37_delay_6 <= io_B_Valid_37_delay_5_1;
    io_A_Valid_6_delay_1_37 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_36 <= io_A_Valid_6_delay_1_37;
    io_A_Valid_6_delay_3_35 <= io_A_Valid_6_delay_2_36;
    io_A_Valid_6_delay_4_34 <= io_A_Valid_6_delay_3_35;
    io_A_Valid_6_delay_5_33 <= io_A_Valid_6_delay_4_34;
    io_A_Valid_6_delay_6_32 <= io_A_Valid_6_delay_5_33;
    io_A_Valid_6_delay_7_31 <= io_A_Valid_6_delay_6_32;
    io_A_Valid_6_delay_8_30 <= io_A_Valid_6_delay_7_31;
    io_A_Valid_6_delay_9_29 <= io_A_Valid_6_delay_8_30;
    io_A_Valid_6_delay_10_28 <= io_A_Valid_6_delay_9_29;
    io_A_Valid_6_delay_11_27 <= io_A_Valid_6_delay_10_28;
    io_A_Valid_6_delay_12_26 <= io_A_Valid_6_delay_11_27;
    io_A_Valid_6_delay_13_25 <= io_A_Valid_6_delay_12_26;
    io_A_Valid_6_delay_14_24 <= io_A_Valid_6_delay_13_25;
    io_A_Valid_6_delay_15_23 <= io_A_Valid_6_delay_14_24;
    io_A_Valid_6_delay_16_22 <= io_A_Valid_6_delay_15_23;
    io_A_Valid_6_delay_17_21 <= io_A_Valid_6_delay_16_22;
    io_A_Valid_6_delay_18_20 <= io_A_Valid_6_delay_17_21;
    io_A_Valid_6_delay_19_19 <= io_A_Valid_6_delay_18_20;
    io_A_Valid_6_delay_20_18 <= io_A_Valid_6_delay_19_19;
    io_A_Valid_6_delay_21_17 <= io_A_Valid_6_delay_20_18;
    io_A_Valid_6_delay_22_16 <= io_A_Valid_6_delay_21_17;
    io_A_Valid_6_delay_23_15 <= io_A_Valid_6_delay_22_16;
    io_A_Valid_6_delay_24_14 <= io_A_Valid_6_delay_23_15;
    io_A_Valid_6_delay_25_13 <= io_A_Valid_6_delay_24_14;
    io_A_Valid_6_delay_26_12 <= io_A_Valid_6_delay_25_13;
    io_A_Valid_6_delay_27_11 <= io_A_Valid_6_delay_26_12;
    io_A_Valid_6_delay_28_10 <= io_A_Valid_6_delay_27_11;
    io_A_Valid_6_delay_29_9 <= io_A_Valid_6_delay_28_10;
    io_A_Valid_6_delay_30_8 <= io_A_Valid_6_delay_29_9;
    io_A_Valid_6_delay_31_7 <= io_A_Valid_6_delay_30_8;
    io_A_Valid_6_delay_32_6 <= io_A_Valid_6_delay_31_7;
    io_A_Valid_6_delay_33_5 <= io_A_Valid_6_delay_32_6;
    io_A_Valid_6_delay_34_4 <= io_A_Valid_6_delay_33_5;
    io_A_Valid_6_delay_35_3 <= io_A_Valid_6_delay_34_4;
    io_A_Valid_6_delay_36_2 <= io_A_Valid_6_delay_35_3;
    io_A_Valid_6_delay_37_1 <= io_A_Valid_6_delay_36_2;
    io_A_Valid_6_delay_38 <= io_A_Valid_6_delay_37_1;
    io_B_Valid_38_delay_1_5 <= io_B_Valid_38;
    io_B_Valid_38_delay_2_4 <= io_B_Valid_38_delay_1_5;
    io_B_Valid_38_delay_3_3 <= io_B_Valid_38_delay_2_4;
    io_B_Valid_38_delay_4_2 <= io_B_Valid_38_delay_3_3;
    io_B_Valid_38_delay_5_1 <= io_B_Valid_38_delay_4_2;
    io_B_Valid_38_delay_6 <= io_B_Valid_38_delay_5_1;
    io_A_Valid_6_delay_1_38 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_37 <= io_A_Valid_6_delay_1_38;
    io_A_Valid_6_delay_3_36 <= io_A_Valid_6_delay_2_37;
    io_A_Valid_6_delay_4_35 <= io_A_Valid_6_delay_3_36;
    io_A_Valid_6_delay_5_34 <= io_A_Valid_6_delay_4_35;
    io_A_Valid_6_delay_6_33 <= io_A_Valid_6_delay_5_34;
    io_A_Valid_6_delay_7_32 <= io_A_Valid_6_delay_6_33;
    io_A_Valid_6_delay_8_31 <= io_A_Valid_6_delay_7_32;
    io_A_Valid_6_delay_9_30 <= io_A_Valid_6_delay_8_31;
    io_A_Valid_6_delay_10_29 <= io_A_Valid_6_delay_9_30;
    io_A_Valid_6_delay_11_28 <= io_A_Valid_6_delay_10_29;
    io_A_Valid_6_delay_12_27 <= io_A_Valid_6_delay_11_28;
    io_A_Valid_6_delay_13_26 <= io_A_Valid_6_delay_12_27;
    io_A_Valid_6_delay_14_25 <= io_A_Valid_6_delay_13_26;
    io_A_Valid_6_delay_15_24 <= io_A_Valid_6_delay_14_25;
    io_A_Valid_6_delay_16_23 <= io_A_Valid_6_delay_15_24;
    io_A_Valid_6_delay_17_22 <= io_A_Valid_6_delay_16_23;
    io_A_Valid_6_delay_18_21 <= io_A_Valid_6_delay_17_22;
    io_A_Valid_6_delay_19_20 <= io_A_Valid_6_delay_18_21;
    io_A_Valid_6_delay_20_19 <= io_A_Valid_6_delay_19_20;
    io_A_Valid_6_delay_21_18 <= io_A_Valid_6_delay_20_19;
    io_A_Valid_6_delay_22_17 <= io_A_Valid_6_delay_21_18;
    io_A_Valid_6_delay_23_16 <= io_A_Valid_6_delay_22_17;
    io_A_Valid_6_delay_24_15 <= io_A_Valid_6_delay_23_16;
    io_A_Valid_6_delay_25_14 <= io_A_Valid_6_delay_24_15;
    io_A_Valid_6_delay_26_13 <= io_A_Valid_6_delay_25_14;
    io_A_Valid_6_delay_27_12 <= io_A_Valid_6_delay_26_13;
    io_A_Valid_6_delay_28_11 <= io_A_Valid_6_delay_27_12;
    io_A_Valid_6_delay_29_10 <= io_A_Valid_6_delay_28_11;
    io_A_Valid_6_delay_30_9 <= io_A_Valid_6_delay_29_10;
    io_A_Valid_6_delay_31_8 <= io_A_Valid_6_delay_30_9;
    io_A_Valid_6_delay_32_7 <= io_A_Valid_6_delay_31_8;
    io_A_Valid_6_delay_33_6 <= io_A_Valid_6_delay_32_7;
    io_A_Valid_6_delay_34_5 <= io_A_Valid_6_delay_33_6;
    io_A_Valid_6_delay_35_4 <= io_A_Valid_6_delay_34_5;
    io_A_Valid_6_delay_36_3 <= io_A_Valid_6_delay_35_4;
    io_A_Valid_6_delay_37_2 <= io_A_Valid_6_delay_36_3;
    io_A_Valid_6_delay_38_1 <= io_A_Valid_6_delay_37_2;
    io_A_Valid_6_delay_39 <= io_A_Valid_6_delay_38_1;
    io_B_Valid_39_delay_1_5 <= io_B_Valid_39;
    io_B_Valid_39_delay_2_4 <= io_B_Valid_39_delay_1_5;
    io_B_Valid_39_delay_3_3 <= io_B_Valid_39_delay_2_4;
    io_B_Valid_39_delay_4_2 <= io_B_Valid_39_delay_3_3;
    io_B_Valid_39_delay_5_1 <= io_B_Valid_39_delay_4_2;
    io_B_Valid_39_delay_6 <= io_B_Valid_39_delay_5_1;
    io_A_Valid_6_delay_1_39 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_38 <= io_A_Valid_6_delay_1_39;
    io_A_Valid_6_delay_3_37 <= io_A_Valid_6_delay_2_38;
    io_A_Valid_6_delay_4_36 <= io_A_Valid_6_delay_3_37;
    io_A_Valid_6_delay_5_35 <= io_A_Valid_6_delay_4_36;
    io_A_Valid_6_delay_6_34 <= io_A_Valid_6_delay_5_35;
    io_A_Valid_6_delay_7_33 <= io_A_Valid_6_delay_6_34;
    io_A_Valid_6_delay_8_32 <= io_A_Valid_6_delay_7_33;
    io_A_Valid_6_delay_9_31 <= io_A_Valid_6_delay_8_32;
    io_A_Valid_6_delay_10_30 <= io_A_Valid_6_delay_9_31;
    io_A_Valid_6_delay_11_29 <= io_A_Valid_6_delay_10_30;
    io_A_Valid_6_delay_12_28 <= io_A_Valid_6_delay_11_29;
    io_A_Valid_6_delay_13_27 <= io_A_Valid_6_delay_12_28;
    io_A_Valid_6_delay_14_26 <= io_A_Valid_6_delay_13_27;
    io_A_Valid_6_delay_15_25 <= io_A_Valid_6_delay_14_26;
    io_A_Valid_6_delay_16_24 <= io_A_Valid_6_delay_15_25;
    io_A_Valid_6_delay_17_23 <= io_A_Valid_6_delay_16_24;
    io_A_Valid_6_delay_18_22 <= io_A_Valid_6_delay_17_23;
    io_A_Valid_6_delay_19_21 <= io_A_Valid_6_delay_18_22;
    io_A_Valid_6_delay_20_20 <= io_A_Valid_6_delay_19_21;
    io_A_Valid_6_delay_21_19 <= io_A_Valid_6_delay_20_20;
    io_A_Valid_6_delay_22_18 <= io_A_Valid_6_delay_21_19;
    io_A_Valid_6_delay_23_17 <= io_A_Valid_6_delay_22_18;
    io_A_Valid_6_delay_24_16 <= io_A_Valid_6_delay_23_17;
    io_A_Valid_6_delay_25_15 <= io_A_Valid_6_delay_24_16;
    io_A_Valid_6_delay_26_14 <= io_A_Valid_6_delay_25_15;
    io_A_Valid_6_delay_27_13 <= io_A_Valid_6_delay_26_14;
    io_A_Valid_6_delay_28_12 <= io_A_Valid_6_delay_27_13;
    io_A_Valid_6_delay_29_11 <= io_A_Valid_6_delay_28_12;
    io_A_Valid_6_delay_30_10 <= io_A_Valid_6_delay_29_11;
    io_A_Valid_6_delay_31_9 <= io_A_Valid_6_delay_30_10;
    io_A_Valid_6_delay_32_8 <= io_A_Valid_6_delay_31_9;
    io_A_Valid_6_delay_33_7 <= io_A_Valid_6_delay_32_8;
    io_A_Valid_6_delay_34_6 <= io_A_Valid_6_delay_33_7;
    io_A_Valid_6_delay_35_5 <= io_A_Valid_6_delay_34_6;
    io_A_Valid_6_delay_36_4 <= io_A_Valid_6_delay_35_5;
    io_A_Valid_6_delay_37_3 <= io_A_Valid_6_delay_36_4;
    io_A_Valid_6_delay_38_2 <= io_A_Valid_6_delay_37_3;
    io_A_Valid_6_delay_39_1 <= io_A_Valid_6_delay_38_2;
    io_A_Valid_6_delay_40 <= io_A_Valid_6_delay_39_1;
    io_B_Valid_40_delay_1_5 <= io_B_Valid_40;
    io_B_Valid_40_delay_2_4 <= io_B_Valid_40_delay_1_5;
    io_B_Valid_40_delay_3_3 <= io_B_Valid_40_delay_2_4;
    io_B_Valid_40_delay_4_2 <= io_B_Valid_40_delay_3_3;
    io_B_Valid_40_delay_5_1 <= io_B_Valid_40_delay_4_2;
    io_B_Valid_40_delay_6 <= io_B_Valid_40_delay_5_1;
    io_A_Valid_6_delay_1_40 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_39 <= io_A_Valid_6_delay_1_40;
    io_A_Valid_6_delay_3_38 <= io_A_Valid_6_delay_2_39;
    io_A_Valid_6_delay_4_37 <= io_A_Valid_6_delay_3_38;
    io_A_Valid_6_delay_5_36 <= io_A_Valid_6_delay_4_37;
    io_A_Valid_6_delay_6_35 <= io_A_Valid_6_delay_5_36;
    io_A_Valid_6_delay_7_34 <= io_A_Valid_6_delay_6_35;
    io_A_Valid_6_delay_8_33 <= io_A_Valid_6_delay_7_34;
    io_A_Valid_6_delay_9_32 <= io_A_Valid_6_delay_8_33;
    io_A_Valid_6_delay_10_31 <= io_A_Valid_6_delay_9_32;
    io_A_Valid_6_delay_11_30 <= io_A_Valid_6_delay_10_31;
    io_A_Valid_6_delay_12_29 <= io_A_Valid_6_delay_11_30;
    io_A_Valid_6_delay_13_28 <= io_A_Valid_6_delay_12_29;
    io_A_Valid_6_delay_14_27 <= io_A_Valid_6_delay_13_28;
    io_A_Valid_6_delay_15_26 <= io_A_Valid_6_delay_14_27;
    io_A_Valid_6_delay_16_25 <= io_A_Valid_6_delay_15_26;
    io_A_Valid_6_delay_17_24 <= io_A_Valid_6_delay_16_25;
    io_A_Valid_6_delay_18_23 <= io_A_Valid_6_delay_17_24;
    io_A_Valid_6_delay_19_22 <= io_A_Valid_6_delay_18_23;
    io_A_Valid_6_delay_20_21 <= io_A_Valid_6_delay_19_22;
    io_A_Valid_6_delay_21_20 <= io_A_Valid_6_delay_20_21;
    io_A_Valid_6_delay_22_19 <= io_A_Valid_6_delay_21_20;
    io_A_Valid_6_delay_23_18 <= io_A_Valid_6_delay_22_19;
    io_A_Valid_6_delay_24_17 <= io_A_Valid_6_delay_23_18;
    io_A_Valid_6_delay_25_16 <= io_A_Valid_6_delay_24_17;
    io_A_Valid_6_delay_26_15 <= io_A_Valid_6_delay_25_16;
    io_A_Valid_6_delay_27_14 <= io_A_Valid_6_delay_26_15;
    io_A_Valid_6_delay_28_13 <= io_A_Valid_6_delay_27_14;
    io_A_Valid_6_delay_29_12 <= io_A_Valid_6_delay_28_13;
    io_A_Valid_6_delay_30_11 <= io_A_Valid_6_delay_29_12;
    io_A_Valid_6_delay_31_10 <= io_A_Valid_6_delay_30_11;
    io_A_Valid_6_delay_32_9 <= io_A_Valid_6_delay_31_10;
    io_A_Valid_6_delay_33_8 <= io_A_Valid_6_delay_32_9;
    io_A_Valid_6_delay_34_7 <= io_A_Valid_6_delay_33_8;
    io_A_Valid_6_delay_35_6 <= io_A_Valid_6_delay_34_7;
    io_A_Valid_6_delay_36_5 <= io_A_Valid_6_delay_35_6;
    io_A_Valid_6_delay_37_4 <= io_A_Valid_6_delay_36_5;
    io_A_Valid_6_delay_38_3 <= io_A_Valid_6_delay_37_4;
    io_A_Valid_6_delay_39_2 <= io_A_Valid_6_delay_38_3;
    io_A_Valid_6_delay_40_1 <= io_A_Valid_6_delay_39_2;
    io_A_Valid_6_delay_41 <= io_A_Valid_6_delay_40_1;
    io_B_Valid_41_delay_1_5 <= io_B_Valid_41;
    io_B_Valid_41_delay_2_4 <= io_B_Valid_41_delay_1_5;
    io_B_Valid_41_delay_3_3 <= io_B_Valid_41_delay_2_4;
    io_B_Valid_41_delay_4_2 <= io_B_Valid_41_delay_3_3;
    io_B_Valid_41_delay_5_1 <= io_B_Valid_41_delay_4_2;
    io_B_Valid_41_delay_6 <= io_B_Valid_41_delay_5_1;
    io_A_Valid_6_delay_1_41 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_40 <= io_A_Valid_6_delay_1_41;
    io_A_Valid_6_delay_3_39 <= io_A_Valid_6_delay_2_40;
    io_A_Valid_6_delay_4_38 <= io_A_Valid_6_delay_3_39;
    io_A_Valid_6_delay_5_37 <= io_A_Valid_6_delay_4_38;
    io_A_Valid_6_delay_6_36 <= io_A_Valid_6_delay_5_37;
    io_A_Valid_6_delay_7_35 <= io_A_Valid_6_delay_6_36;
    io_A_Valid_6_delay_8_34 <= io_A_Valid_6_delay_7_35;
    io_A_Valid_6_delay_9_33 <= io_A_Valid_6_delay_8_34;
    io_A_Valid_6_delay_10_32 <= io_A_Valid_6_delay_9_33;
    io_A_Valid_6_delay_11_31 <= io_A_Valid_6_delay_10_32;
    io_A_Valid_6_delay_12_30 <= io_A_Valid_6_delay_11_31;
    io_A_Valid_6_delay_13_29 <= io_A_Valid_6_delay_12_30;
    io_A_Valid_6_delay_14_28 <= io_A_Valid_6_delay_13_29;
    io_A_Valid_6_delay_15_27 <= io_A_Valid_6_delay_14_28;
    io_A_Valid_6_delay_16_26 <= io_A_Valid_6_delay_15_27;
    io_A_Valid_6_delay_17_25 <= io_A_Valid_6_delay_16_26;
    io_A_Valid_6_delay_18_24 <= io_A_Valid_6_delay_17_25;
    io_A_Valid_6_delay_19_23 <= io_A_Valid_6_delay_18_24;
    io_A_Valid_6_delay_20_22 <= io_A_Valid_6_delay_19_23;
    io_A_Valid_6_delay_21_21 <= io_A_Valid_6_delay_20_22;
    io_A_Valid_6_delay_22_20 <= io_A_Valid_6_delay_21_21;
    io_A_Valid_6_delay_23_19 <= io_A_Valid_6_delay_22_20;
    io_A_Valid_6_delay_24_18 <= io_A_Valid_6_delay_23_19;
    io_A_Valid_6_delay_25_17 <= io_A_Valid_6_delay_24_18;
    io_A_Valid_6_delay_26_16 <= io_A_Valid_6_delay_25_17;
    io_A_Valid_6_delay_27_15 <= io_A_Valid_6_delay_26_16;
    io_A_Valid_6_delay_28_14 <= io_A_Valid_6_delay_27_15;
    io_A_Valid_6_delay_29_13 <= io_A_Valid_6_delay_28_14;
    io_A_Valid_6_delay_30_12 <= io_A_Valid_6_delay_29_13;
    io_A_Valid_6_delay_31_11 <= io_A_Valid_6_delay_30_12;
    io_A_Valid_6_delay_32_10 <= io_A_Valid_6_delay_31_11;
    io_A_Valid_6_delay_33_9 <= io_A_Valid_6_delay_32_10;
    io_A_Valid_6_delay_34_8 <= io_A_Valid_6_delay_33_9;
    io_A_Valid_6_delay_35_7 <= io_A_Valid_6_delay_34_8;
    io_A_Valid_6_delay_36_6 <= io_A_Valid_6_delay_35_7;
    io_A_Valid_6_delay_37_5 <= io_A_Valid_6_delay_36_6;
    io_A_Valid_6_delay_38_4 <= io_A_Valid_6_delay_37_5;
    io_A_Valid_6_delay_39_3 <= io_A_Valid_6_delay_38_4;
    io_A_Valid_6_delay_40_2 <= io_A_Valid_6_delay_39_3;
    io_A_Valid_6_delay_41_1 <= io_A_Valid_6_delay_40_2;
    io_A_Valid_6_delay_42 <= io_A_Valid_6_delay_41_1;
    io_B_Valid_42_delay_1_5 <= io_B_Valid_42;
    io_B_Valid_42_delay_2_4 <= io_B_Valid_42_delay_1_5;
    io_B_Valid_42_delay_3_3 <= io_B_Valid_42_delay_2_4;
    io_B_Valid_42_delay_4_2 <= io_B_Valid_42_delay_3_3;
    io_B_Valid_42_delay_5_1 <= io_B_Valid_42_delay_4_2;
    io_B_Valid_42_delay_6 <= io_B_Valid_42_delay_5_1;
    io_A_Valid_6_delay_1_42 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_41 <= io_A_Valid_6_delay_1_42;
    io_A_Valid_6_delay_3_40 <= io_A_Valid_6_delay_2_41;
    io_A_Valid_6_delay_4_39 <= io_A_Valid_6_delay_3_40;
    io_A_Valid_6_delay_5_38 <= io_A_Valid_6_delay_4_39;
    io_A_Valid_6_delay_6_37 <= io_A_Valid_6_delay_5_38;
    io_A_Valid_6_delay_7_36 <= io_A_Valid_6_delay_6_37;
    io_A_Valid_6_delay_8_35 <= io_A_Valid_6_delay_7_36;
    io_A_Valid_6_delay_9_34 <= io_A_Valid_6_delay_8_35;
    io_A_Valid_6_delay_10_33 <= io_A_Valid_6_delay_9_34;
    io_A_Valid_6_delay_11_32 <= io_A_Valid_6_delay_10_33;
    io_A_Valid_6_delay_12_31 <= io_A_Valid_6_delay_11_32;
    io_A_Valid_6_delay_13_30 <= io_A_Valid_6_delay_12_31;
    io_A_Valid_6_delay_14_29 <= io_A_Valid_6_delay_13_30;
    io_A_Valid_6_delay_15_28 <= io_A_Valid_6_delay_14_29;
    io_A_Valid_6_delay_16_27 <= io_A_Valid_6_delay_15_28;
    io_A_Valid_6_delay_17_26 <= io_A_Valid_6_delay_16_27;
    io_A_Valid_6_delay_18_25 <= io_A_Valid_6_delay_17_26;
    io_A_Valid_6_delay_19_24 <= io_A_Valid_6_delay_18_25;
    io_A_Valid_6_delay_20_23 <= io_A_Valid_6_delay_19_24;
    io_A_Valid_6_delay_21_22 <= io_A_Valid_6_delay_20_23;
    io_A_Valid_6_delay_22_21 <= io_A_Valid_6_delay_21_22;
    io_A_Valid_6_delay_23_20 <= io_A_Valid_6_delay_22_21;
    io_A_Valid_6_delay_24_19 <= io_A_Valid_6_delay_23_20;
    io_A_Valid_6_delay_25_18 <= io_A_Valid_6_delay_24_19;
    io_A_Valid_6_delay_26_17 <= io_A_Valid_6_delay_25_18;
    io_A_Valid_6_delay_27_16 <= io_A_Valid_6_delay_26_17;
    io_A_Valid_6_delay_28_15 <= io_A_Valid_6_delay_27_16;
    io_A_Valid_6_delay_29_14 <= io_A_Valid_6_delay_28_15;
    io_A_Valid_6_delay_30_13 <= io_A_Valid_6_delay_29_14;
    io_A_Valid_6_delay_31_12 <= io_A_Valid_6_delay_30_13;
    io_A_Valid_6_delay_32_11 <= io_A_Valid_6_delay_31_12;
    io_A_Valid_6_delay_33_10 <= io_A_Valid_6_delay_32_11;
    io_A_Valid_6_delay_34_9 <= io_A_Valid_6_delay_33_10;
    io_A_Valid_6_delay_35_8 <= io_A_Valid_6_delay_34_9;
    io_A_Valid_6_delay_36_7 <= io_A_Valid_6_delay_35_8;
    io_A_Valid_6_delay_37_6 <= io_A_Valid_6_delay_36_7;
    io_A_Valid_6_delay_38_5 <= io_A_Valid_6_delay_37_6;
    io_A_Valid_6_delay_39_4 <= io_A_Valid_6_delay_38_5;
    io_A_Valid_6_delay_40_3 <= io_A_Valid_6_delay_39_4;
    io_A_Valid_6_delay_41_2 <= io_A_Valid_6_delay_40_3;
    io_A_Valid_6_delay_42_1 <= io_A_Valid_6_delay_41_2;
    io_A_Valid_6_delay_43 <= io_A_Valid_6_delay_42_1;
    io_B_Valid_43_delay_1_5 <= io_B_Valid_43;
    io_B_Valid_43_delay_2_4 <= io_B_Valid_43_delay_1_5;
    io_B_Valid_43_delay_3_3 <= io_B_Valid_43_delay_2_4;
    io_B_Valid_43_delay_4_2 <= io_B_Valid_43_delay_3_3;
    io_B_Valid_43_delay_5_1 <= io_B_Valid_43_delay_4_2;
    io_B_Valid_43_delay_6 <= io_B_Valid_43_delay_5_1;
    io_A_Valid_6_delay_1_43 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_42 <= io_A_Valid_6_delay_1_43;
    io_A_Valid_6_delay_3_41 <= io_A_Valid_6_delay_2_42;
    io_A_Valid_6_delay_4_40 <= io_A_Valid_6_delay_3_41;
    io_A_Valid_6_delay_5_39 <= io_A_Valid_6_delay_4_40;
    io_A_Valid_6_delay_6_38 <= io_A_Valid_6_delay_5_39;
    io_A_Valid_6_delay_7_37 <= io_A_Valid_6_delay_6_38;
    io_A_Valid_6_delay_8_36 <= io_A_Valid_6_delay_7_37;
    io_A_Valid_6_delay_9_35 <= io_A_Valid_6_delay_8_36;
    io_A_Valid_6_delay_10_34 <= io_A_Valid_6_delay_9_35;
    io_A_Valid_6_delay_11_33 <= io_A_Valid_6_delay_10_34;
    io_A_Valid_6_delay_12_32 <= io_A_Valid_6_delay_11_33;
    io_A_Valid_6_delay_13_31 <= io_A_Valid_6_delay_12_32;
    io_A_Valid_6_delay_14_30 <= io_A_Valid_6_delay_13_31;
    io_A_Valid_6_delay_15_29 <= io_A_Valid_6_delay_14_30;
    io_A_Valid_6_delay_16_28 <= io_A_Valid_6_delay_15_29;
    io_A_Valid_6_delay_17_27 <= io_A_Valid_6_delay_16_28;
    io_A_Valid_6_delay_18_26 <= io_A_Valid_6_delay_17_27;
    io_A_Valid_6_delay_19_25 <= io_A_Valid_6_delay_18_26;
    io_A_Valid_6_delay_20_24 <= io_A_Valid_6_delay_19_25;
    io_A_Valid_6_delay_21_23 <= io_A_Valid_6_delay_20_24;
    io_A_Valid_6_delay_22_22 <= io_A_Valid_6_delay_21_23;
    io_A_Valid_6_delay_23_21 <= io_A_Valid_6_delay_22_22;
    io_A_Valid_6_delay_24_20 <= io_A_Valid_6_delay_23_21;
    io_A_Valid_6_delay_25_19 <= io_A_Valid_6_delay_24_20;
    io_A_Valid_6_delay_26_18 <= io_A_Valid_6_delay_25_19;
    io_A_Valid_6_delay_27_17 <= io_A_Valid_6_delay_26_18;
    io_A_Valid_6_delay_28_16 <= io_A_Valid_6_delay_27_17;
    io_A_Valid_6_delay_29_15 <= io_A_Valid_6_delay_28_16;
    io_A_Valid_6_delay_30_14 <= io_A_Valid_6_delay_29_15;
    io_A_Valid_6_delay_31_13 <= io_A_Valid_6_delay_30_14;
    io_A_Valid_6_delay_32_12 <= io_A_Valid_6_delay_31_13;
    io_A_Valid_6_delay_33_11 <= io_A_Valid_6_delay_32_12;
    io_A_Valid_6_delay_34_10 <= io_A_Valid_6_delay_33_11;
    io_A_Valid_6_delay_35_9 <= io_A_Valid_6_delay_34_10;
    io_A_Valid_6_delay_36_8 <= io_A_Valid_6_delay_35_9;
    io_A_Valid_6_delay_37_7 <= io_A_Valid_6_delay_36_8;
    io_A_Valid_6_delay_38_6 <= io_A_Valid_6_delay_37_7;
    io_A_Valid_6_delay_39_5 <= io_A_Valid_6_delay_38_6;
    io_A_Valid_6_delay_40_4 <= io_A_Valid_6_delay_39_5;
    io_A_Valid_6_delay_41_3 <= io_A_Valid_6_delay_40_4;
    io_A_Valid_6_delay_42_2 <= io_A_Valid_6_delay_41_3;
    io_A_Valid_6_delay_43_1 <= io_A_Valid_6_delay_42_2;
    io_A_Valid_6_delay_44 <= io_A_Valid_6_delay_43_1;
    io_B_Valid_44_delay_1_5 <= io_B_Valid_44;
    io_B_Valid_44_delay_2_4 <= io_B_Valid_44_delay_1_5;
    io_B_Valid_44_delay_3_3 <= io_B_Valid_44_delay_2_4;
    io_B_Valid_44_delay_4_2 <= io_B_Valid_44_delay_3_3;
    io_B_Valid_44_delay_5_1 <= io_B_Valid_44_delay_4_2;
    io_B_Valid_44_delay_6 <= io_B_Valid_44_delay_5_1;
    io_A_Valid_6_delay_1_44 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_43 <= io_A_Valid_6_delay_1_44;
    io_A_Valid_6_delay_3_42 <= io_A_Valid_6_delay_2_43;
    io_A_Valid_6_delay_4_41 <= io_A_Valid_6_delay_3_42;
    io_A_Valid_6_delay_5_40 <= io_A_Valid_6_delay_4_41;
    io_A_Valid_6_delay_6_39 <= io_A_Valid_6_delay_5_40;
    io_A_Valid_6_delay_7_38 <= io_A_Valid_6_delay_6_39;
    io_A_Valid_6_delay_8_37 <= io_A_Valid_6_delay_7_38;
    io_A_Valid_6_delay_9_36 <= io_A_Valid_6_delay_8_37;
    io_A_Valid_6_delay_10_35 <= io_A_Valid_6_delay_9_36;
    io_A_Valid_6_delay_11_34 <= io_A_Valid_6_delay_10_35;
    io_A_Valid_6_delay_12_33 <= io_A_Valid_6_delay_11_34;
    io_A_Valid_6_delay_13_32 <= io_A_Valid_6_delay_12_33;
    io_A_Valid_6_delay_14_31 <= io_A_Valid_6_delay_13_32;
    io_A_Valid_6_delay_15_30 <= io_A_Valid_6_delay_14_31;
    io_A_Valid_6_delay_16_29 <= io_A_Valid_6_delay_15_30;
    io_A_Valid_6_delay_17_28 <= io_A_Valid_6_delay_16_29;
    io_A_Valid_6_delay_18_27 <= io_A_Valid_6_delay_17_28;
    io_A_Valid_6_delay_19_26 <= io_A_Valid_6_delay_18_27;
    io_A_Valid_6_delay_20_25 <= io_A_Valid_6_delay_19_26;
    io_A_Valid_6_delay_21_24 <= io_A_Valid_6_delay_20_25;
    io_A_Valid_6_delay_22_23 <= io_A_Valid_6_delay_21_24;
    io_A_Valid_6_delay_23_22 <= io_A_Valid_6_delay_22_23;
    io_A_Valid_6_delay_24_21 <= io_A_Valid_6_delay_23_22;
    io_A_Valid_6_delay_25_20 <= io_A_Valid_6_delay_24_21;
    io_A_Valid_6_delay_26_19 <= io_A_Valid_6_delay_25_20;
    io_A_Valid_6_delay_27_18 <= io_A_Valid_6_delay_26_19;
    io_A_Valid_6_delay_28_17 <= io_A_Valid_6_delay_27_18;
    io_A_Valid_6_delay_29_16 <= io_A_Valid_6_delay_28_17;
    io_A_Valid_6_delay_30_15 <= io_A_Valid_6_delay_29_16;
    io_A_Valid_6_delay_31_14 <= io_A_Valid_6_delay_30_15;
    io_A_Valid_6_delay_32_13 <= io_A_Valid_6_delay_31_14;
    io_A_Valid_6_delay_33_12 <= io_A_Valid_6_delay_32_13;
    io_A_Valid_6_delay_34_11 <= io_A_Valid_6_delay_33_12;
    io_A_Valid_6_delay_35_10 <= io_A_Valid_6_delay_34_11;
    io_A_Valid_6_delay_36_9 <= io_A_Valid_6_delay_35_10;
    io_A_Valid_6_delay_37_8 <= io_A_Valid_6_delay_36_9;
    io_A_Valid_6_delay_38_7 <= io_A_Valid_6_delay_37_8;
    io_A_Valid_6_delay_39_6 <= io_A_Valid_6_delay_38_7;
    io_A_Valid_6_delay_40_5 <= io_A_Valid_6_delay_39_6;
    io_A_Valid_6_delay_41_4 <= io_A_Valid_6_delay_40_5;
    io_A_Valid_6_delay_42_3 <= io_A_Valid_6_delay_41_4;
    io_A_Valid_6_delay_43_2 <= io_A_Valid_6_delay_42_3;
    io_A_Valid_6_delay_44_1 <= io_A_Valid_6_delay_43_2;
    io_A_Valid_6_delay_45 <= io_A_Valid_6_delay_44_1;
    io_B_Valid_45_delay_1_5 <= io_B_Valid_45;
    io_B_Valid_45_delay_2_4 <= io_B_Valid_45_delay_1_5;
    io_B_Valid_45_delay_3_3 <= io_B_Valid_45_delay_2_4;
    io_B_Valid_45_delay_4_2 <= io_B_Valid_45_delay_3_3;
    io_B_Valid_45_delay_5_1 <= io_B_Valid_45_delay_4_2;
    io_B_Valid_45_delay_6 <= io_B_Valid_45_delay_5_1;
    io_A_Valid_6_delay_1_45 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_44 <= io_A_Valid_6_delay_1_45;
    io_A_Valid_6_delay_3_43 <= io_A_Valid_6_delay_2_44;
    io_A_Valid_6_delay_4_42 <= io_A_Valid_6_delay_3_43;
    io_A_Valid_6_delay_5_41 <= io_A_Valid_6_delay_4_42;
    io_A_Valid_6_delay_6_40 <= io_A_Valid_6_delay_5_41;
    io_A_Valid_6_delay_7_39 <= io_A_Valid_6_delay_6_40;
    io_A_Valid_6_delay_8_38 <= io_A_Valid_6_delay_7_39;
    io_A_Valid_6_delay_9_37 <= io_A_Valid_6_delay_8_38;
    io_A_Valid_6_delay_10_36 <= io_A_Valid_6_delay_9_37;
    io_A_Valid_6_delay_11_35 <= io_A_Valid_6_delay_10_36;
    io_A_Valid_6_delay_12_34 <= io_A_Valid_6_delay_11_35;
    io_A_Valid_6_delay_13_33 <= io_A_Valid_6_delay_12_34;
    io_A_Valid_6_delay_14_32 <= io_A_Valid_6_delay_13_33;
    io_A_Valid_6_delay_15_31 <= io_A_Valid_6_delay_14_32;
    io_A_Valid_6_delay_16_30 <= io_A_Valid_6_delay_15_31;
    io_A_Valid_6_delay_17_29 <= io_A_Valid_6_delay_16_30;
    io_A_Valid_6_delay_18_28 <= io_A_Valid_6_delay_17_29;
    io_A_Valid_6_delay_19_27 <= io_A_Valid_6_delay_18_28;
    io_A_Valid_6_delay_20_26 <= io_A_Valid_6_delay_19_27;
    io_A_Valid_6_delay_21_25 <= io_A_Valid_6_delay_20_26;
    io_A_Valid_6_delay_22_24 <= io_A_Valid_6_delay_21_25;
    io_A_Valid_6_delay_23_23 <= io_A_Valid_6_delay_22_24;
    io_A_Valid_6_delay_24_22 <= io_A_Valid_6_delay_23_23;
    io_A_Valid_6_delay_25_21 <= io_A_Valid_6_delay_24_22;
    io_A_Valid_6_delay_26_20 <= io_A_Valid_6_delay_25_21;
    io_A_Valid_6_delay_27_19 <= io_A_Valid_6_delay_26_20;
    io_A_Valid_6_delay_28_18 <= io_A_Valid_6_delay_27_19;
    io_A_Valid_6_delay_29_17 <= io_A_Valid_6_delay_28_18;
    io_A_Valid_6_delay_30_16 <= io_A_Valid_6_delay_29_17;
    io_A_Valid_6_delay_31_15 <= io_A_Valid_6_delay_30_16;
    io_A_Valid_6_delay_32_14 <= io_A_Valid_6_delay_31_15;
    io_A_Valid_6_delay_33_13 <= io_A_Valid_6_delay_32_14;
    io_A_Valid_6_delay_34_12 <= io_A_Valid_6_delay_33_13;
    io_A_Valid_6_delay_35_11 <= io_A_Valid_6_delay_34_12;
    io_A_Valid_6_delay_36_10 <= io_A_Valid_6_delay_35_11;
    io_A_Valid_6_delay_37_9 <= io_A_Valid_6_delay_36_10;
    io_A_Valid_6_delay_38_8 <= io_A_Valid_6_delay_37_9;
    io_A_Valid_6_delay_39_7 <= io_A_Valid_6_delay_38_8;
    io_A_Valid_6_delay_40_6 <= io_A_Valid_6_delay_39_7;
    io_A_Valid_6_delay_41_5 <= io_A_Valid_6_delay_40_6;
    io_A_Valid_6_delay_42_4 <= io_A_Valid_6_delay_41_5;
    io_A_Valid_6_delay_43_3 <= io_A_Valid_6_delay_42_4;
    io_A_Valid_6_delay_44_2 <= io_A_Valid_6_delay_43_3;
    io_A_Valid_6_delay_45_1 <= io_A_Valid_6_delay_44_2;
    io_A_Valid_6_delay_46 <= io_A_Valid_6_delay_45_1;
    io_B_Valid_46_delay_1_5 <= io_B_Valid_46;
    io_B_Valid_46_delay_2_4 <= io_B_Valid_46_delay_1_5;
    io_B_Valid_46_delay_3_3 <= io_B_Valid_46_delay_2_4;
    io_B_Valid_46_delay_4_2 <= io_B_Valid_46_delay_3_3;
    io_B_Valid_46_delay_5_1 <= io_B_Valid_46_delay_4_2;
    io_B_Valid_46_delay_6 <= io_B_Valid_46_delay_5_1;
    io_A_Valid_6_delay_1_46 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_45 <= io_A_Valid_6_delay_1_46;
    io_A_Valid_6_delay_3_44 <= io_A_Valid_6_delay_2_45;
    io_A_Valid_6_delay_4_43 <= io_A_Valid_6_delay_3_44;
    io_A_Valid_6_delay_5_42 <= io_A_Valid_6_delay_4_43;
    io_A_Valid_6_delay_6_41 <= io_A_Valid_6_delay_5_42;
    io_A_Valid_6_delay_7_40 <= io_A_Valid_6_delay_6_41;
    io_A_Valid_6_delay_8_39 <= io_A_Valid_6_delay_7_40;
    io_A_Valid_6_delay_9_38 <= io_A_Valid_6_delay_8_39;
    io_A_Valid_6_delay_10_37 <= io_A_Valid_6_delay_9_38;
    io_A_Valid_6_delay_11_36 <= io_A_Valid_6_delay_10_37;
    io_A_Valid_6_delay_12_35 <= io_A_Valid_6_delay_11_36;
    io_A_Valid_6_delay_13_34 <= io_A_Valid_6_delay_12_35;
    io_A_Valid_6_delay_14_33 <= io_A_Valid_6_delay_13_34;
    io_A_Valid_6_delay_15_32 <= io_A_Valid_6_delay_14_33;
    io_A_Valid_6_delay_16_31 <= io_A_Valid_6_delay_15_32;
    io_A_Valid_6_delay_17_30 <= io_A_Valid_6_delay_16_31;
    io_A_Valid_6_delay_18_29 <= io_A_Valid_6_delay_17_30;
    io_A_Valid_6_delay_19_28 <= io_A_Valid_6_delay_18_29;
    io_A_Valid_6_delay_20_27 <= io_A_Valid_6_delay_19_28;
    io_A_Valid_6_delay_21_26 <= io_A_Valid_6_delay_20_27;
    io_A_Valid_6_delay_22_25 <= io_A_Valid_6_delay_21_26;
    io_A_Valid_6_delay_23_24 <= io_A_Valid_6_delay_22_25;
    io_A_Valid_6_delay_24_23 <= io_A_Valid_6_delay_23_24;
    io_A_Valid_6_delay_25_22 <= io_A_Valid_6_delay_24_23;
    io_A_Valid_6_delay_26_21 <= io_A_Valid_6_delay_25_22;
    io_A_Valid_6_delay_27_20 <= io_A_Valid_6_delay_26_21;
    io_A_Valid_6_delay_28_19 <= io_A_Valid_6_delay_27_20;
    io_A_Valid_6_delay_29_18 <= io_A_Valid_6_delay_28_19;
    io_A_Valid_6_delay_30_17 <= io_A_Valid_6_delay_29_18;
    io_A_Valid_6_delay_31_16 <= io_A_Valid_6_delay_30_17;
    io_A_Valid_6_delay_32_15 <= io_A_Valid_6_delay_31_16;
    io_A_Valid_6_delay_33_14 <= io_A_Valid_6_delay_32_15;
    io_A_Valid_6_delay_34_13 <= io_A_Valid_6_delay_33_14;
    io_A_Valid_6_delay_35_12 <= io_A_Valid_6_delay_34_13;
    io_A_Valid_6_delay_36_11 <= io_A_Valid_6_delay_35_12;
    io_A_Valid_6_delay_37_10 <= io_A_Valid_6_delay_36_11;
    io_A_Valid_6_delay_38_9 <= io_A_Valid_6_delay_37_10;
    io_A_Valid_6_delay_39_8 <= io_A_Valid_6_delay_38_9;
    io_A_Valid_6_delay_40_7 <= io_A_Valid_6_delay_39_8;
    io_A_Valid_6_delay_41_6 <= io_A_Valid_6_delay_40_7;
    io_A_Valid_6_delay_42_5 <= io_A_Valid_6_delay_41_6;
    io_A_Valid_6_delay_43_4 <= io_A_Valid_6_delay_42_5;
    io_A_Valid_6_delay_44_3 <= io_A_Valid_6_delay_43_4;
    io_A_Valid_6_delay_45_2 <= io_A_Valid_6_delay_44_3;
    io_A_Valid_6_delay_46_1 <= io_A_Valid_6_delay_45_2;
    io_A_Valid_6_delay_47 <= io_A_Valid_6_delay_46_1;
    io_B_Valid_47_delay_1_5 <= io_B_Valid_47;
    io_B_Valid_47_delay_2_4 <= io_B_Valid_47_delay_1_5;
    io_B_Valid_47_delay_3_3 <= io_B_Valid_47_delay_2_4;
    io_B_Valid_47_delay_4_2 <= io_B_Valid_47_delay_3_3;
    io_B_Valid_47_delay_5_1 <= io_B_Valid_47_delay_4_2;
    io_B_Valid_47_delay_6 <= io_B_Valid_47_delay_5_1;
    io_A_Valid_6_delay_1_47 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_46 <= io_A_Valid_6_delay_1_47;
    io_A_Valid_6_delay_3_45 <= io_A_Valid_6_delay_2_46;
    io_A_Valid_6_delay_4_44 <= io_A_Valid_6_delay_3_45;
    io_A_Valid_6_delay_5_43 <= io_A_Valid_6_delay_4_44;
    io_A_Valid_6_delay_6_42 <= io_A_Valid_6_delay_5_43;
    io_A_Valid_6_delay_7_41 <= io_A_Valid_6_delay_6_42;
    io_A_Valid_6_delay_8_40 <= io_A_Valid_6_delay_7_41;
    io_A_Valid_6_delay_9_39 <= io_A_Valid_6_delay_8_40;
    io_A_Valid_6_delay_10_38 <= io_A_Valid_6_delay_9_39;
    io_A_Valid_6_delay_11_37 <= io_A_Valid_6_delay_10_38;
    io_A_Valid_6_delay_12_36 <= io_A_Valid_6_delay_11_37;
    io_A_Valid_6_delay_13_35 <= io_A_Valid_6_delay_12_36;
    io_A_Valid_6_delay_14_34 <= io_A_Valid_6_delay_13_35;
    io_A_Valid_6_delay_15_33 <= io_A_Valid_6_delay_14_34;
    io_A_Valid_6_delay_16_32 <= io_A_Valid_6_delay_15_33;
    io_A_Valid_6_delay_17_31 <= io_A_Valid_6_delay_16_32;
    io_A_Valid_6_delay_18_30 <= io_A_Valid_6_delay_17_31;
    io_A_Valid_6_delay_19_29 <= io_A_Valid_6_delay_18_30;
    io_A_Valid_6_delay_20_28 <= io_A_Valid_6_delay_19_29;
    io_A_Valid_6_delay_21_27 <= io_A_Valid_6_delay_20_28;
    io_A_Valid_6_delay_22_26 <= io_A_Valid_6_delay_21_27;
    io_A_Valid_6_delay_23_25 <= io_A_Valid_6_delay_22_26;
    io_A_Valid_6_delay_24_24 <= io_A_Valid_6_delay_23_25;
    io_A_Valid_6_delay_25_23 <= io_A_Valid_6_delay_24_24;
    io_A_Valid_6_delay_26_22 <= io_A_Valid_6_delay_25_23;
    io_A_Valid_6_delay_27_21 <= io_A_Valid_6_delay_26_22;
    io_A_Valid_6_delay_28_20 <= io_A_Valid_6_delay_27_21;
    io_A_Valid_6_delay_29_19 <= io_A_Valid_6_delay_28_20;
    io_A_Valid_6_delay_30_18 <= io_A_Valid_6_delay_29_19;
    io_A_Valid_6_delay_31_17 <= io_A_Valid_6_delay_30_18;
    io_A_Valid_6_delay_32_16 <= io_A_Valid_6_delay_31_17;
    io_A_Valid_6_delay_33_15 <= io_A_Valid_6_delay_32_16;
    io_A_Valid_6_delay_34_14 <= io_A_Valid_6_delay_33_15;
    io_A_Valid_6_delay_35_13 <= io_A_Valid_6_delay_34_14;
    io_A_Valid_6_delay_36_12 <= io_A_Valid_6_delay_35_13;
    io_A_Valid_6_delay_37_11 <= io_A_Valid_6_delay_36_12;
    io_A_Valid_6_delay_38_10 <= io_A_Valid_6_delay_37_11;
    io_A_Valid_6_delay_39_9 <= io_A_Valid_6_delay_38_10;
    io_A_Valid_6_delay_40_8 <= io_A_Valid_6_delay_39_9;
    io_A_Valid_6_delay_41_7 <= io_A_Valid_6_delay_40_8;
    io_A_Valid_6_delay_42_6 <= io_A_Valid_6_delay_41_7;
    io_A_Valid_6_delay_43_5 <= io_A_Valid_6_delay_42_6;
    io_A_Valid_6_delay_44_4 <= io_A_Valid_6_delay_43_5;
    io_A_Valid_6_delay_45_3 <= io_A_Valid_6_delay_44_4;
    io_A_Valid_6_delay_46_2 <= io_A_Valid_6_delay_45_3;
    io_A_Valid_6_delay_47_1 <= io_A_Valid_6_delay_46_2;
    io_A_Valid_6_delay_48 <= io_A_Valid_6_delay_47_1;
    io_B_Valid_48_delay_1_5 <= io_B_Valid_48;
    io_B_Valid_48_delay_2_4 <= io_B_Valid_48_delay_1_5;
    io_B_Valid_48_delay_3_3 <= io_B_Valid_48_delay_2_4;
    io_B_Valid_48_delay_4_2 <= io_B_Valid_48_delay_3_3;
    io_B_Valid_48_delay_5_1 <= io_B_Valid_48_delay_4_2;
    io_B_Valid_48_delay_6 <= io_B_Valid_48_delay_5_1;
    io_A_Valid_6_delay_1_48 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_47 <= io_A_Valid_6_delay_1_48;
    io_A_Valid_6_delay_3_46 <= io_A_Valid_6_delay_2_47;
    io_A_Valid_6_delay_4_45 <= io_A_Valid_6_delay_3_46;
    io_A_Valid_6_delay_5_44 <= io_A_Valid_6_delay_4_45;
    io_A_Valid_6_delay_6_43 <= io_A_Valid_6_delay_5_44;
    io_A_Valid_6_delay_7_42 <= io_A_Valid_6_delay_6_43;
    io_A_Valid_6_delay_8_41 <= io_A_Valid_6_delay_7_42;
    io_A_Valid_6_delay_9_40 <= io_A_Valid_6_delay_8_41;
    io_A_Valid_6_delay_10_39 <= io_A_Valid_6_delay_9_40;
    io_A_Valid_6_delay_11_38 <= io_A_Valid_6_delay_10_39;
    io_A_Valid_6_delay_12_37 <= io_A_Valid_6_delay_11_38;
    io_A_Valid_6_delay_13_36 <= io_A_Valid_6_delay_12_37;
    io_A_Valid_6_delay_14_35 <= io_A_Valid_6_delay_13_36;
    io_A_Valid_6_delay_15_34 <= io_A_Valid_6_delay_14_35;
    io_A_Valid_6_delay_16_33 <= io_A_Valid_6_delay_15_34;
    io_A_Valid_6_delay_17_32 <= io_A_Valid_6_delay_16_33;
    io_A_Valid_6_delay_18_31 <= io_A_Valid_6_delay_17_32;
    io_A_Valid_6_delay_19_30 <= io_A_Valid_6_delay_18_31;
    io_A_Valid_6_delay_20_29 <= io_A_Valid_6_delay_19_30;
    io_A_Valid_6_delay_21_28 <= io_A_Valid_6_delay_20_29;
    io_A_Valid_6_delay_22_27 <= io_A_Valid_6_delay_21_28;
    io_A_Valid_6_delay_23_26 <= io_A_Valid_6_delay_22_27;
    io_A_Valid_6_delay_24_25 <= io_A_Valid_6_delay_23_26;
    io_A_Valid_6_delay_25_24 <= io_A_Valid_6_delay_24_25;
    io_A_Valid_6_delay_26_23 <= io_A_Valid_6_delay_25_24;
    io_A_Valid_6_delay_27_22 <= io_A_Valid_6_delay_26_23;
    io_A_Valid_6_delay_28_21 <= io_A_Valid_6_delay_27_22;
    io_A_Valid_6_delay_29_20 <= io_A_Valid_6_delay_28_21;
    io_A_Valid_6_delay_30_19 <= io_A_Valid_6_delay_29_20;
    io_A_Valid_6_delay_31_18 <= io_A_Valid_6_delay_30_19;
    io_A_Valid_6_delay_32_17 <= io_A_Valid_6_delay_31_18;
    io_A_Valid_6_delay_33_16 <= io_A_Valid_6_delay_32_17;
    io_A_Valid_6_delay_34_15 <= io_A_Valid_6_delay_33_16;
    io_A_Valid_6_delay_35_14 <= io_A_Valid_6_delay_34_15;
    io_A_Valid_6_delay_36_13 <= io_A_Valid_6_delay_35_14;
    io_A_Valid_6_delay_37_12 <= io_A_Valid_6_delay_36_13;
    io_A_Valid_6_delay_38_11 <= io_A_Valid_6_delay_37_12;
    io_A_Valid_6_delay_39_10 <= io_A_Valid_6_delay_38_11;
    io_A_Valid_6_delay_40_9 <= io_A_Valid_6_delay_39_10;
    io_A_Valid_6_delay_41_8 <= io_A_Valid_6_delay_40_9;
    io_A_Valid_6_delay_42_7 <= io_A_Valid_6_delay_41_8;
    io_A_Valid_6_delay_43_6 <= io_A_Valid_6_delay_42_7;
    io_A_Valid_6_delay_44_5 <= io_A_Valid_6_delay_43_6;
    io_A_Valid_6_delay_45_4 <= io_A_Valid_6_delay_44_5;
    io_A_Valid_6_delay_46_3 <= io_A_Valid_6_delay_45_4;
    io_A_Valid_6_delay_47_2 <= io_A_Valid_6_delay_46_3;
    io_A_Valid_6_delay_48_1 <= io_A_Valid_6_delay_47_2;
    io_A_Valid_6_delay_49 <= io_A_Valid_6_delay_48_1;
    io_B_Valid_49_delay_1_5 <= io_B_Valid_49;
    io_B_Valid_49_delay_2_4 <= io_B_Valid_49_delay_1_5;
    io_B_Valid_49_delay_3_3 <= io_B_Valid_49_delay_2_4;
    io_B_Valid_49_delay_4_2 <= io_B_Valid_49_delay_3_3;
    io_B_Valid_49_delay_5_1 <= io_B_Valid_49_delay_4_2;
    io_B_Valid_49_delay_6 <= io_B_Valid_49_delay_5_1;
    io_A_Valid_6_delay_1_49 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_48 <= io_A_Valid_6_delay_1_49;
    io_A_Valid_6_delay_3_47 <= io_A_Valid_6_delay_2_48;
    io_A_Valid_6_delay_4_46 <= io_A_Valid_6_delay_3_47;
    io_A_Valid_6_delay_5_45 <= io_A_Valid_6_delay_4_46;
    io_A_Valid_6_delay_6_44 <= io_A_Valid_6_delay_5_45;
    io_A_Valid_6_delay_7_43 <= io_A_Valid_6_delay_6_44;
    io_A_Valid_6_delay_8_42 <= io_A_Valid_6_delay_7_43;
    io_A_Valid_6_delay_9_41 <= io_A_Valid_6_delay_8_42;
    io_A_Valid_6_delay_10_40 <= io_A_Valid_6_delay_9_41;
    io_A_Valid_6_delay_11_39 <= io_A_Valid_6_delay_10_40;
    io_A_Valid_6_delay_12_38 <= io_A_Valid_6_delay_11_39;
    io_A_Valid_6_delay_13_37 <= io_A_Valid_6_delay_12_38;
    io_A_Valid_6_delay_14_36 <= io_A_Valid_6_delay_13_37;
    io_A_Valid_6_delay_15_35 <= io_A_Valid_6_delay_14_36;
    io_A_Valid_6_delay_16_34 <= io_A_Valid_6_delay_15_35;
    io_A_Valid_6_delay_17_33 <= io_A_Valid_6_delay_16_34;
    io_A_Valid_6_delay_18_32 <= io_A_Valid_6_delay_17_33;
    io_A_Valid_6_delay_19_31 <= io_A_Valid_6_delay_18_32;
    io_A_Valid_6_delay_20_30 <= io_A_Valid_6_delay_19_31;
    io_A_Valid_6_delay_21_29 <= io_A_Valid_6_delay_20_30;
    io_A_Valid_6_delay_22_28 <= io_A_Valid_6_delay_21_29;
    io_A_Valid_6_delay_23_27 <= io_A_Valid_6_delay_22_28;
    io_A_Valid_6_delay_24_26 <= io_A_Valid_6_delay_23_27;
    io_A_Valid_6_delay_25_25 <= io_A_Valid_6_delay_24_26;
    io_A_Valid_6_delay_26_24 <= io_A_Valid_6_delay_25_25;
    io_A_Valid_6_delay_27_23 <= io_A_Valid_6_delay_26_24;
    io_A_Valid_6_delay_28_22 <= io_A_Valid_6_delay_27_23;
    io_A_Valid_6_delay_29_21 <= io_A_Valid_6_delay_28_22;
    io_A_Valid_6_delay_30_20 <= io_A_Valid_6_delay_29_21;
    io_A_Valid_6_delay_31_19 <= io_A_Valid_6_delay_30_20;
    io_A_Valid_6_delay_32_18 <= io_A_Valid_6_delay_31_19;
    io_A_Valid_6_delay_33_17 <= io_A_Valid_6_delay_32_18;
    io_A_Valid_6_delay_34_16 <= io_A_Valid_6_delay_33_17;
    io_A_Valid_6_delay_35_15 <= io_A_Valid_6_delay_34_16;
    io_A_Valid_6_delay_36_14 <= io_A_Valid_6_delay_35_15;
    io_A_Valid_6_delay_37_13 <= io_A_Valid_6_delay_36_14;
    io_A_Valid_6_delay_38_12 <= io_A_Valid_6_delay_37_13;
    io_A_Valid_6_delay_39_11 <= io_A_Valid_6_delay_38_12;
    io_A_Valid_6_delay_40_10 <= io_A_Valid_6_delay_39_11;
    io_A_Valid_6_delay_41_9 <= io_A_Valid_6_delay_40_10;
    io_A_Valid_6_delay_42_8 <= io_A_Valid_6_delay_41_9;
    io_A_Valid_6_delay_43_7 <= io_A_Valid_6_delay_42_8;
    io_A_Valid_6_delay_44_6 <= io_A_Valid_6_delay_43_7;
    io_A_Valid_6_delay_45_5 <= io_A_Valid_6_delay_44_6;
    io_A_Valid_6_delay_46_4 <= io_A_Valid_6_delay_45_5;
    io_A_Valid_6_delay_47_3 <= io_A_Valid_6_delay_46_4;
    io_A_Valid_6_delay_48_2 <= io_A_Valid_6_delay_47_3;
    io_A_Valid_6_delay_49_1 <= io_A_Valid_6_delay_48_2;
    io_A_Valid_6_delay_50 <= io_A_Valid_6_delay_49_1;
    io_B_Valid_50_delay_1_5 <= io_B_Valid_50;
    io_B_Valid_50_delay_2_4 <= io_B_Valid_50_delay_1_5;
    io_B_Valid_50_delay_3_3 <= io_B_Valid_50_delay_2_4;
    io_B_Valid_50_delay_4_2 <= io_B_Valid_50_delay_3_3;
    io_B_Valid_50_delay_5_1 <= io_B_Valid_50_delay_4_2;
    io_B_Valid_50_delay_6 <= io_B_Valid_50_delay_5_1;
    io_A_Valid_6_delay_1_50 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_49 <= io_A_Valid_6_delay_1_50;
    io_A_Valid_6_delay_3_48 <= io_A_Valid_6_delay_2_49;
    io_A_Valid_6_delay_4_47 <= io_A_Valid_6_delay_3_48;
    io_A_Valid_6_delay_5_46 <= io_A_Valid_6_delay_4_47;
    io_A_Valid_6_delay_6_45 <= io_A_Valid_6_delay_5_46;
    io_A_Valid_6_delay_7_44 <= io_A_Valid_6_delay_6_45;
    io_A_Valid_6_delay_8_43 <= io_A_Valid_6_delay_7_44;
    io_A_Valid_6_delay_9_42 <= io_A_Valid_6_delay_8_43;
    io_A_Valid_6_delay_10_41 <= io_A_Valid_6_delay_9_42;
    io_A_Valid_6_delay_11_40 <= io_A_Valid_6_delay_10_41;
    io_A_Valid_6_delay_12_39 <= io_A_Valid_6_delay_11_40;
    io_A_Valid_6_delay_13_38 <= io_A_Valid_6_delay_12_39;
    io_A_Valid_6_delay_14_37 <= io_A_Valid_6_delay_13_38;
    io_A_Valid_6_delay_15_36 <= io_A_Valid_6_delay_14_37;
    io_A_Valid_6_delay_16_35 <= io_A_Valid_6_delay_15_36;
    io_A_Valid_6_delay_17_34 <= io_A_Valid_6_delay_16_35;
    io_A_Valid_6_delay_18_33 <= io_A_Valid_6_delay_17_34;
    io_A_Valid_6_delay_19_32 <= io_A_Valid_6_delay_18_33;
    io_A_Valid_6_delay_20_31 <= io_A_Valid_6_delay_19_32;
    io_A_Valid_6_delay_21_30 <= io_A_Valid_6_delay_20_31;
    io_A_Valid_6_delay_22_29 <= io_A_Valid_6_delay_21_30;
    io_A_Valid_6_delay_23_28 <= io_A_Valid_6_delay_22_29;
    io_A_Valid_6_delay_24_27 <= io_A_Valid_6_delay_23_28;
    io_A_Valid_6_delay_25_26 <= io_A_Valid_6_delay_24_27;
    io_A_Valid_6_delay_26_25 <= io_A_Valid_6_delay_25_26;
    io_A_Valid_6_delay_27_24 <= io_A_Valid_6_delay_26_25;
    io_A_Valid_6_delay_28_23 <= io_A_Valid_6_delay_27_24;
    io_A_Valid_6_delay_29_22 <= io_A_Valid_6_delay_28_23;
    io_A_Valid_6_delay_30_21 <= io_A_Valid_6_delay_29_22;
    io_A_Valid_6_delay_31_20 <= io_A_Valid_6_delay_30_21;
    io_A_Valid_6_delay_32_19 <= io_A_Valid_6_delay_31_20;
    io_A_Valid_6_delay_33_18 <= io_A_Valid_6_delay_32_19;
    io_A_Valid_6_delay_34_17 <= io_A_Valid_6_delay_33_18;
    io_A_Valid_6_delay_35_16 <= io_A_Valid_6_delay_34_17;
    io_A_Valid_6_delay_36_15 <= io_A_Valid_6_delay_35_16;
    io_A_Valid_6_delay_37_14 <= io_A_Valid_6_delay_36_15;
    io_A_Valid_6_delay_38_13 <= io_A_Valid_6_delay_37_14;
    io_A_Valid_6_delay_39_12 <= io_A_Valid_6_delay_38_13;
    io_A_Valid_6_delay_40_11 <= io_A_Valid_6_delay_39_12;
    io_A_Valid_6_delay_41_10 <= io_A_Valid_6_delay_40_11;
    io_A_Valid_6_delay_42_9 <= io_A_Valid_6_delay_41_10;
    io_A_Valid_6_delay_43_8 <= io_A_Valid_6_delay_42_9;
    io_A_Valid_6_delay_44_7 <= io_A_Valid_6_delay_43_8;
    io_A_Valid_6_delay_45_6 <= io_A_Valid_6_delay_44_7;
    io_A_Valid_6_delay_46_5 <= io_A_Valid_6_delay_45_6;
    io_A_Valid_6_delay_47_4 <= io_A_Valid_6_delay_46_5;
    io_A_Valid_6_delay_48_3 <= io_A_Valid_6_delay_47_4;
    io_A_Valid_6_delay_49_2 <= io_A_Valid_6_delay_48_3;
    io_A_Valid_6_delay_50_1 <= io_A_Valid_6_delay_49_2;
    io_A_Valid_6_delay_51 <= io_A_Valid_6_delay_50_1;
    io_B_Valid_51_delay_1_5 <= io_B_Valid_51;
    io_B_Valid_51_delay_2_4 <= io_B_Valid_51_delay_1_5;
    io_B_Valid_51_delay_3_3 <= io_B_Valid_51_delay_2_4;
    io_B_Valid_51_delay_4_2 <= io_B_Valid_51_delay_3_3;
    io_B_Valid_51_delay_5_1 <= io_B_Valid_51_delay_4_2;
    io_B_Valid_51_delay_6 <= io_B_Valid_51_delay_5_1;
    io_A_Valid_6_delay_1_51 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_50 <= io_A_Valid_6_delay_1_51;
    io_A_Valid_6_delay_3_49 <= io_A_Valid_6_delay_2_50;
    io_A_Valid_6_delay_4_48 <= io_A_Valid_6_delay_3_49;
    io_A_Valid_6_delay_5_47 <= io_A_Valid_6_delay_4_48;
    io_A_Valid_6_delay_6_46 <= io_A_Valid_6_delay_5_47;
    io_A_Valid_6_delay_7_45 <= io_A_Valid_6_delay_6_46;
    io_A_Valid_6_delay_8_44 <= io_A_Valid_6_delay_7_45;
    io_A_Valid_6_delay_9_43 <= io_A_Valid_6_delay_8_44;
    io_A_Valid_6_delay_10_42 <= io_A_Valid_6_delay_9_43;
    io_A_Valid_6_delay_11_41 <= io_A_Valid_6_delay_10_42;
    io_A_Valid_6_delay_12_40 <= io_A_Valid_6_delay_11_41;
    io_A_Valid_6_delay_13_39 <= io_A_Valid_6_delay_12_40;
    io_A_Valid_6_delay_14_38 <= io_A_Valid_6_delay_13_39;
    io_A_Valid_6_delay_15_37 <= io_A_Valid_6_delay_14_38;
    io_A_Valid_6_delay_16_36 <= io_A_Valid_6_delay_15_37;
    io_A_Valid_6_delay_17_35 <= io_A_Valid_6_delay_16_36;
    io_A_Valid_6_delay_18_34 <= io_A_Valid_6_delay_17_35;
    io_A_Valid_6_delay_19_33 <= io_A_Valid_6_delay_18_34;
    io_A_Valid_6_delay_20_32 <= io_A_Valid_6_delay_19_33;
    io_A_Valid_6_delay_21_31 <= io_A_Valid_6_delay_20_32;
    io_A_Valid_6_delay_22_30 <= io_A_Valid_6_delay_21_31;
    io_A_Valid_6_delay_23_29 <= io_A_Valid_6_delay_22_30;
    io_A_Valid_6_delay_24_28 <= io_A_Valid_6_delay_23_29;
    io_A_Valid_6_delay_25_27 <= io_A_Valid_6_delay_24_28;
    io_A_Valid_6_delay_26_26 <= io_A_Valid_6_delay_25_27;
    io_A_Valid_6_delay_27_25 <= io_A_Valid_6_delay_26_26;
    io_A_Valid_6_delay_28_24 <= io_A_Valid_6_delay_27_25;
    io_A_Valid_6_delay_29_23 <= io_A_Valid_6_delay_28_24;
    io_A_Valid_6_delay_30_22 <= io_A_Valid_6_delay_29_23;
    io_A_Valid_6_delay_31_21 <= io_A_Valid_6_delay_30_22;
    io_A_Valid_6_delay_32_20 <= io_A_Valid_6_delay_31_21;
    io_A_Valid_6_delay_33_19 <= io_A_Valid_6_delay_32_20;
    io_A_Valid_6_delay_34_18 <= io_A_Valid_6_delay_33_19;
    io_A_Valid_6_delay_35_17 <= io_A_Valid_6_delay_34_18;
    io_A_Valid_6_delay_36_16 <= io_A_Valid_6_delay_35_17;
    io_A_Valid_6_delay_37_15 <= io_A_Valid_6_delay_36_16;
    io_A_Valid_6_delay_38_14 <= io_A_Valid_6_delay_37_15;
    io_A_Valid_6_delay_39_13 <= io_A_Valid_6_delay_38_14;
    io_A_Valid_6_delay_40_12 <= io_A_Valid_6_delay_39_13;
    io_A_Valid_6_delay_41_11 <= io_A_Valid_6_delay_40_12;
    io_A_Valid_6_delay_42_10 <= io_A_Valid_6_delay_41_11;
    io_A_Valid_6_delay_43_9 <= io_A_Valid_6_delay_42_10;
    io_A_Valid_6_delay_44_8 <= io_A_Valid_6_delay_43_9;
    io_A_Valid_6_delay_45_7 <= io_A_Valid_6_delay_44_8;
    io_A_Valid_6_delay_46_6 <= io_A_Valid_6_delay_45_7;
    io_A_Valid_6_delay_47_5 <= io_A_Valid_6_delay_46_6;
    io_A_Valid_6_delay_48_4 <= io_A_Valid_6_delay_47_5;
    io_A_Valid_6_delay_49_3 <= io_A_Valid_6_delay_48_4;
    io_A_Valid_6_delay_50_2 <= io_A_Valid_6_delay_49_3;
    io_A_Valid_6_delay_51_1 <= io_A_Valid_6_delay_50_2;
    io_A_Valid_6_delay_52 <= io_A_Valid_6_delay_51_1;
    io_B_Valid_52_delay_1_5 <= io_B_Valid_52;
    io_B_Valid_52_delay_2_4 <= io_B_Valid_52_delay_1_5;
    io_B_Valid_52_delay_3_3 <= io_B_Valid_52_delay_2_4;
    io_B_Valid_52_delay_4_2 <= io_B_Valid_52_delay_3_3;
    io_B_Valid_52_delay_5_1 <= io_B_Valid_52_delay_4_2;
    io_B_Valid_52_delay_6 <= io_B_Valid_52_delay_5_1;
    io_A_Valid_6_delay_1_52 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_51 <= io_A_Valid_6_delay_1_52;
    io_A_Valid_6_delay_3_50 <= io_A_Valid_6_delay_2_51;
    io_A_Valid_6_delay_4_49 <= io_A_Valid_6_delay_3_50;
    io_A_Valid_6_delay_5_48 <= io_A_Valid_6_delay_4_49;
    io_A_Valid_6_delay_6_47 <= io_A_Valid_6_delay_5_48;
    io_A_Valid_6_delay_7_46 <= io_A_Valid_6_delay_6_47;
    io_A_Valid_6_delay_8_45 <= io_A_Valid_6_delay_7_46;
    io_A_Valid_6_delay_9_44 <= io_A_Valid_6_delay_8_45;
    io_A_Valid_6_delay_10_43 <= io_A_Valid_6_delay_9_44;
    io_A_Valid_6_delay_11_42 <= io_A_Valid_6_delay_10_43;
    io_A_Valid_6_delay_12_41 <= io_A_Valid_6_delay_11_42;
    io_A_Valid_6_delay_13_40 <= io_A_Valid_6_delay_12_41;
    io_A_Valid_6_delay_14_39 <= io_A_Valid_6_delay_13_40;
    io_A_Valid_6_delay_15_38 <= io_A_Valid_6_delay_14_39;
    io_A_Valid_6_delay_16_37 <= io_A_Valid_6_delay_15_38;
    io_A_Valid_6_delay_17_36 <= io_A_Valid_6_delay_16_37;
    io_A_Valid_6_delay_18_35 <= io_A_Valid_6_delay_17_36;
    io_A_Valid_6_delay_19_34 <= io_A_Valid_6_delay_18_35;
    io_A_Valid_6_delay_20_33 <= io_A_Valid_6_delay_19_34;
    io_A_Valid_6_delay_21_32 <= io_A_Valid_6_delay_20_33;
    io_A_Valid_6_delay_22_31 <= io_A_Valid_6_delay_21_32;
    io_A_Valid_6_delay_23_30 <= io_A_Valid_6_delay_22_31;
    io_A_Valid_6_delay_24_29 <= io_A_Valid_6_delay_23_30;
    io_A_Valid_6_delay_25_28 <= io_A_Valid_6_delay_24_29;
    io_A_Valid_6_delay_26_27 <= io_A_Valid_6_delay_25_28;
    io_A_Valid_6_delay_27_26 <= io_A_Valid_6_delay_26_27;
    io_A_Valid_6_delay_28_25 <= io_A_Valid_6_delay_27_26;
    io_A_Valid_6_delay_29_24 <= io_A_Valid_6_delay_28_25;
    io_A_Valid_6_delay_30_23 <= io_A_Valid_6_delay_29_24;
    io_A_Valid_6_delay_31_22 <= io_A_Valid_6_delay_30_23;
    io_A_Valid_6_delay_32_21 <= io_A_Valid_6_delay_31_22;
    io_A_Valid_6_delay_33_20 <= io_A_Valid_6_delay_32_21;
    io_A_Valid_6_delay_34_19 <= io_A_Valid_6_delay_33_20;
    io_A_Valid_6_delay_35_18 <= io_A_Valid_6_delay_34_19;
    io_A_Valid_6_delay_36_17 <= io_A_Valid_6_delay_35_18;
    io_A_Valid_6_delay_37_16 <= io_A_Valid_6_delay_36_17;
    io_A_Valid_6_delay_38_15 <= io_A_Valid_6_delay_37_16;
    io_A_Valid_6_delay_39_14 <= io_A_Valid_6_delay_38_15;
    io_A_Valid_6_delay_40_13 <= io_A_Valid_6_delay_39_14;
    io_A_Valid_6_delay_41_12 <= io_A_Valid_6_delay_40_13;
    io_A_Valid_6_delay_42_11 <= io_A_Valid_6_delay_41_12;
    io_A_Valid_6_delay_43_10 <= io_A_Valid_6_delay_42_11;
    io_A_Valid_6_delay_44_9 <= io_A_Valid_6_delay_43_10;
    io_A_Valid_6_delay_45_8 <= io_A_Valid_6_delay_44_9;
    io_A_Valid_6_delay_46_7 <= io_A_Valid_6_delay_45_8;
    io_A_Valid_6_delay_47_6 <= io_A_Valid_6_delay_46_7;
    io_A_Valid_6_delay_48_5 <= io_A_Valid_6_delay_47_6;
    io_A_Valid_6_delay_49_4 <= io_A_Valid_6_delay_48_5;
    io_A_Valid_6_delay_50_3 <= io_A_Valid_6_delay_49_4;
    io_A_Valid_6_delay_51_2 <= io_A_Valid_6_delay_50_3;
    io_A_Valid_6_delay_52_1 <= io_A_Valid_6_delay_51_2;
    io_A_Valid_6_delay_53 <= io_A_Valid_6_delay_52_1;
    io_B_Valid_53_delay_1_5 <= io_B_Valid_53;
    io_B_Valid_53_delay_2_4 <= io_B_Valid_53_delay_1_5;
    io_B_Valid_53_delay_3_3 <= io_B_Valid_53_delay_2_4;
    io_B_Valid_53_delay_4_2 <= io_B_Valid_53_delay_3_3;
    io_B_Valid_53_delay_5_1 <= io_B_Valid_53_delay_4_2;
    io_B_Valid_53_delay_6 <= io_B_Valid_53_delay_5_1;
    io_A_Valid_6_delay_1_53 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_52 <= io_A_Valid_6_delay_1_53;
    io_A_Valid_6_delay_3_51 <= io_A_Valid_6_delay_2_52;
    io_A_Valid_6_delay_4_50 <= io_A_Valid_6_delay_3_51;
    io_A_Valid_6_delay_5_49 <= io_A_Valid_6_delay_4_50;
    io_A_Valid_6_delay_6_48 <= io_A_Valid_6_delay_5_49;
    io_A_Valid_6_delay_7_47 <= io_A_Valid_6_delay_6_48;
    io_A_Valid_6_delay_8_46 <= io_A_Valid_6_delay_7_47;
    io_A_Valid_6_delay_9_45 <= io_A_Valid_6_delay_8_46;
    io_A_Valid_6_delay_10_44 <= io_A_Valid_6_delay_9_45;
    io_A_Valid_6_delay_11_43 <= io_A_Valid_6_delay_10_44;
    io_A_Valid_6_delay_12_42 <= io_A_Valid_6_delay_11_43;
    io_A_Valid_6_delay_13_41 <= io_A_Valid_6_delay_12_42;
    io_A_Valid_6_delay_14_40 <= io_A_Valid_6_delay_13_41;
    io_A_Valid_6_delay_15_39 <= io_A_Valid_6_delay_14_40;
    io_A_Valid_6_delay_16_38 <= io_A_Valid_6_delay_15_39;
    io_A_Valid_6_delay_17_37 <= io_A_Valid_6_delay_16_38;
    io_A_Valid_6_delay_18_36 <= io_A_Valid_6_delay_17_37;
    io_A_Valid_6_delay_19_35 <= io_A_Valid_6_delay_18_36;
    io_A_Valid_6_delay_20_34 <= io_A_Valid_6_delay_19_35;
    io_A_Valid_6_delay_21_33 <= io_A_Valid_6_delay_20_34;
    io_A_Valid_6_delay_22_32 <= io_A_Valid_6_delay_21_33;
    io_A_Valid_6_delay_23_31 <= io_A_Valid_6_delay_22_32;
    io_A_Valid_6_delay_24_30 <= io_A_Valid_6_delay_23_31;
    io_A_Valid_6_delay_25_29 <= io_A_Valid_6_delay_24_30;
    io_A_Valid_6_delay_26_28 <= io_A_Valid_6_delay_25_29;
    io_A_Valid_6_delay_27_27 <= io_A_Valid_6_delay_26_28;
    io_A_Valid_6_delay_28_26 <= io_A_Valid_6_delay_27_27;
    io_A_Valid_6_delay_29_25 <= io_A_Valid_6_delay_28_26;
    io_A_Valid_6_delay_30_24 <= io_A_Valid_6_delay_29_25;
    io_A_Valid_6_delay_31_23 <= io_A_Valid_6_delay_30_24;
    io_A_Valid_6_delay_32_22 <= io_A_Valid_6_delay_31_23;
    io_A_Valid_6_delay_33_21 <= io_A_Valid_6_delay_32_22;
    io_A_Valid_6_delay_34_20 <= io_A_Valid_6_delay_33_21;
    io_A_Valid_6_delay_35_19 <= io_A_Valid_6_delay_34_20;
    io_A_Valid_6_delay_36_18 <= io_A_Valid_6_delay_35_19;
    io_A_Valid_6_delay_37_17 <= io_A_Valid_6_delay_36_18;
    io_A_Valid_6_delay_38_16 <= io_A_Valid_6_delay_37_17;
    io_A_Valid_6_delay_39_15 <= io_A_Valid_6_delay_38_16;
    io_A_Valid_6_delay_40_14 <= io_A_Valid_6_delay_39_15;
    io_A_Valid_6_delay_41_13 <= io_A_Valid_6_delay_40_14;
    io_A_Valid_6_delay_42_12 <= io_A_Valid_6_delay_41_13;
    io_A_Valid_6_delay_43_11 <= io_A_Valid_6_delay_42_12;
    io_A_Valid_6_delay_44_10 <= io_A_Valid_6_delay_43_11;
    io_A_Valid_6_delay_45_9 <= io_A_Valid_6_delay_44_10;
    io_A_Valid_6_delay_46_8 <= io_A_Valid_6_delay_45_9;
    io_A_Valid_6_delay_47_7 <= io_A_Valid_6_delay_46_8;
    io_A_Valid_6_delay_48_6 <= io_A_Valid_6_delay_47_7;
    io_A_Valid_6_delay_49_5 <= io_A_Valid_6_delay_48_6;
    io_A_Valid_6_delay_50_4 <= io_A_Valid_6_delay_49_5;
    io_A_Valid_6_delay_51_3 <= io_A_Valid_6_delay_50_4;
    io_A_Valid_6_delay_52_2 <= io_A_Valid_6_delay_51_3;
    io_A_Valid_6_delay_53_1 <= io_A_Valid_6_delay_52_2;
    io_A_Valid_6_delay_54 <= io_A_Valid_6_delay_53_1;
    io_B_Valid_54_delay_1_5 <= io_B_Valid_54;
    io_B_Valid_54_delay_2_4 <= io_B_Valid_54_delay_1_5;
    io_B_Valid_54_delay_3_3 <= io_B_Valid_54_delay_2_4;
    io_B_Valid_54_delay_4_2 <= io_B_Valid_54_delay_3_3;
    io_B_Valid_54_delay_5_1 <= io_B_Valid_54_delay_4_2;
    io_B_Valid_54_delay_6 <= io_B_Valid_54_delay_5_1;
    io_A_Valid_6_delay_1_54 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_53 <= io_A_Valid_6_delay_1_54;
    io_A_Valid_6_delay_3_52 <= io_A_Valid_6_delay_2_53;
    io_A_Valid_6_delay_4_51 <= io_A_Valid_6_delay_3_52;
    io_A_Valid_6_delay_5_50 <= io_A_Valid_6_delay_4_51;
    io_A_Valid_6_delay_6_49 <= io_A_Valid_6_delay_5_50;
    io_A_Valid_6_delay_7_48 <= io_A_Valid_6_delay_6_49;
    io_A_Valid_6_delay_8_47 <= io_A_Valid_6_delay_7_48;
    io_A_Valid_6_delay_9_46 <= io_A_Valid_6_delay_8_47;
    io_A_Valid_6_delay_10_45 <= io_A_Valid_6_delay_9_46;
    io_A_Valid_6_delay_11_44 <= io_A_Valid_6_delay_10_45;
    io_A_Valid_6_delay_12_43 <= io_A_Valid_6_delay_11_44;
    io_A_Valid_6_delay_13_42 <= io_A_Valid_6_delay_12_43;
    io_A_Valid_6_delay_14_41 <= io_A_Valid_6_delay_13_42;
    io_A_Valid_6_delay_15_40 <= io_A_Valid_6_delay_14_41;
    io_A_Valid_6_delay_16_39 <= io_A_Valid_6_delay_15_40;
    io_A_Valid_6_delay_17_38 <= io_A_Valid_6_delay_16_39;
    io_A_Valid_6_delay_18_37 <= io_A_Valid_6_delay_17_38;
    io_A_Valid_6_delay_19_36 <= io_A_Valid_6_delay_18_37;
    io_A_Valid_6_delay_20_35 <= io_A_Valid_6_delay_19_36;
    io_A_Valid_6_delay_21_34 <= io_A_Valid_6_delay_20_35;
    io_A_Valid_6_delay_22_33 <= io_A_Valid_6_delay_21_34;
    io_A_Valid_6_delay_23_32 <= io_A_Valid_6_delay_22_33;
    io_A_Valid_6_delay_24_31 <= io_A_Valid_6_delay_23_32;
    io_A_Valid_6_delay_25_30 <= io_A_Valid_6_delay_24_31;
    io_A_Valid_6_delay_26_29 <= io_A_Valid_6_delay_25_30;
    io_A_Valid_6_delay_27_28 <= io_A_Valid_6_delay_26_29;
    io_A_Valid_6_delay_28_27 <= io_A_Valid_6_delay_27_28;
    io_A_Valid_6_delay_29_26 <= io_A_Valid_6_delay_28_27;
    io_A_Valid_6_delay_30_25 <= io_A_Valid_6_delay_29_26;
    io_A_Valid_6_delay_31_24 <= io_A_Valid_6_delay_30_25;
    io_A_Valid_6_delay_32_23 <= io_A_Valid_6_delay_31_24;
    io_A_Valid_6_delay_33_22 <= io_A_Valid_6_delay_32_23;
    io_A_Valid_6_delay_34_21 <= io_A_Valid_6_delay_33_22;
    io_A_Valid_6_delay_35_20 <= io_A_Valid_6_delay_34_21;
    io_A_Valid_6_delay_36_19 <= io_A_Valid_6_delay_35_20;
    io_A_Valid_6_delay_37_18 <= io_A_Valid_6_delay_36_19;
    io_A_Valid_6_delay_38_17 <= io_A_Valid_6_delay_37_18;
    io_A_Valid_6_delay_39_16 <= io_A_Valid_6_delay_38_17;
    io_A_Valid_6_delay_40_15 <= io_A_Valid_6_delay_39_16;
    io_A_Valid_6_delay_41_14 <= io_A_Valid_6_delay_40_15;
    io_A_Valid_6_delay_42_13 <= io_A_Valid_6_delay_41_14;
    io_A_Valid_6_delay_43_12 <= io_A_Valid_6_delay_42_13;
    io_A_Valid_6_delay_44_11 <= io_A_Valid_6_delay_43_12;
    io_A_Valid_6_delay_45_10 <= io_A_Valid_6_delay_44_11;
    io_A_Valid_6_delay_46_9 <= io_A_Valid_6_delay_45_10;
    io_A_Valid_6_delay_47_8 <= io_A_Valid_6_delay_46_9;
    io_A_Valid_6_delay_48_7 <= io_A_Valid_6_delay_47_8;
    io_A_Valid_6_delay_49_6 <= io_A_Valid_6_delay_48_7;
    io_A_Valid_6_delay_50_5 <= io_A_Valid_6_delay_49_6;
    io_A_Valid_6_delay_51_4 <= io_A_Valid_6_delay_50_5;
    io_A_Valid_6_delay_52_3 <= io_A_Valid_6_delay_51_4;
    io_A_Valid_6_delay_53_2 <= io_A_Valid_6_delay_52_3;
    io_A_Valid_6_delay_54_1 <= io_A_Valid_6_delay_53_2;
    io_A_Valid_6_delay_55 <= io_A_Valid_6_delay_54_1;
    io_B_Valid_55_delay_1_5 <= io_B_Valid_55;
    io_B_Valid_55_delay_2_4 <= io_B_Valid_55_delay_1_5;
    io_B_Valid_55_delay_3_3 <= io_B_Valid_55_delay_2_4;
    io_B_Valid_55_delay_4_2 <= io_B_Valid_55_delay_3_3;
    io_B_Valid_55_delay_5_1 <= io_B_Valid_55_delay_4_2;
    io_B_Valid_55_delay_6 <= io_B_Valid_55_delay_5_1;
    io_A_Valid_6_delay_1_55 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_54 <= io_A_Valid_6_delay_1_55;
    io_A_Valid_6_delay_3_53 <= io_A_Valid_6_delay_2_54;
    io_A_Valid_6_delay_4_52 <= io_A_Valid_6_delay_3_53;
    io_A_Valid_6_delay_5_51 <= io_A_Valid_6_delay_4_52;
    io_A_Valid_6_delay_6_50 <= io_A_Valid_6_delay_5_51;
    io_A_Valid_6_delay_7_49 <= io_A_Valid_6_delay_6_50;
    io_A_Valid_6_delay_8_48 <= io_A_Valid_6_delay_7_49;
    io_A_Valid_6_delay_9_47 <= io_A_Valid_6_delay_8_48;
    io_A_Valid_6_delay_10_46 <= io_A_Valid_6_delay_9_47;
    io_A_Valid_6_delay_11_45 <= io_A_Valid_6_delay_10_46;
    io_A_Valid_6_delay_12_44 <= io_A_Valid_6_delay_11_45;
    io_A_Valid_6_delay_13_43 <= io_A_Valid_6_delay_12_44;
    io_A_Valid_6_delay_14_42 <= io_A_Valid_6_delay_13_43;
    io_A_Valid_6_delay_15_41 <= io_A_Valid_6_delay_14_42;
    io_A_Valid_6_delay_16_40 <= io_A_Valid_6_delay_15_41;
    io_A_Valid_6_delay_17_39 <= io_A_Valid_6_delay_16_40;
    io_A_Valid_6_delay_18_38 <= io_A_Valid_6_delay_17_39;
    io_A_Valid_6_delay_19_37 <= io_A_Valid_6_delay_18_38;
    io_A_Valid_6_delay_20_36 <= io_A_Valid_6_delay_19_37;
    io_A_Valid_6_delay_21_35 <= io_A_Valid_6_delay_20_36;
    io_A_Valid_6_delay_22_34 <= io_A_Valid_6_delay_21_35;
    io_A_Valid_6_delay_23_33 <= io_A_Valid_6_delay_22_34;
    io_A_Valid_6_delay_24_32 <= io_A_Valid_6_delay_23_33;
    io_A_Valid_6_delay_25_31 <= io_A_Valid_6_delay_24_32;
    io_A_Valid_6_delay_26_30 <= io_A_Valid_6_delay_25_31;
    io_A_Valid_6_delay_27_29 <= io_A_Valid_6_delay_26_30;
    io_A_Valid_6_delay_28_28 <= io_A_Valid_6_delay_27_29;
    io_A_Valid_6_delay_29_27 <= io_A_Valid_6_delay_28_28;
    io_A_Valid_6_delay_30_26 <= io_A_Valid_6_delay_29_27;
    io_A_Valid_6_delay_31_25 <= io_A_Valid_6_delay_30_26;
    io_A_Valid_6_delay_32_24 <= io_A_Valid_6_delay_31_25;
    io_A_Valid_6_delay_33_23 <= io_A_Valid_6_delay_32_24;
    io_A_Valid_6_delay_34_22 <= io_A_Valid_6_delay_33_23;
    io_A_Valid_6_delay_35_21 <= io_A_Valid_6_delay_34_22;
    io_A_Valid_6_delay_36_20 <= io_A_Valid_6_delay_35_21;
    io_A_Valid_6_delay_37_19 <= io_A_Valid_6_delay_36_20;
    io_A_Valid_6_delay_38_18 <= io_A_Valid_6_delay_37_19;
    io_A_Valid_6_delay_39_17 <= io_A_Valid_6_delay_38_18;
    io_A_Valid_6_delay_40_16 <= io_A_Valid_6_delay_39_17;
    io_A_Valid_6_delay_41_15 <= io_A_Valid_6_delay_40_16;
    io_A_Valid_6_delay_42_14 <= io_A_Valid_6_delay_41_15;
    io_A_Valid_6_delay_43_13 <= io_A_Valid_6_delay_42_14;
    io_A_Valid_6_delay_44_12 <= io_A_Valid_6_delay_43_13;
    io_A_Valid_6_delay_45_11 <= io_A_Valid_6_delay_44_12;
    io_A_Valid_6_delay_46_10 <= io_A_Valid_6_delay_45_11;
    io_A_Valid_6_delay_47_9 <= io_A_Valid_6_delay_46_10;
    io_A_Valid_6_delay_48_8 <= io_A_Valid_6_delay_47_9;
    io_A_Valid_6_delay_49_7 <= io_A_Valid_6_delay_48_8;
    io_A_Valid_6_delay_50_6 <= io_A_Valid_6_delay_49_7;
    io_A_Valid_6_delay_51_5 <= io_A_Valid_6_delay_50_6;
    io_A_Valid_6_delay_52_4 <= io_A_Valid_6_delay_51_5;
    io_A_Valid_6_delay_53_3 <= io_A_Valid_6_delay_52_4;
    io_A_Valid_6_delay_54_2 <= io_A_Valid_6_delay_53_3;
    io_A_Valid_6_delay_55_1 <= io_A_Valid_6_delay_54_2;
    io_A_Valid_6_delay_56 <= io_A_Valid_6_delay_55_1;
    io_B_Valid_56_delay_1_5 <= io_B_Valid_56;
    io_B_Valid_56_delay_2_4 <= io_B_Valid_56_delay_1_5;
    io_B_Valid_56_delay_3_3 <= io_B_Valid_56_delay_2_4;
    io_B_Valid_56_delay_4_2 <= io_B_Valid_56_delay_3_3;
    io_B_Valid_56_delay_5_1 <= io_B_Valid_56_delay_4_2;
    io_B_Valid_56_delay_6 <= io_B_Valid_56_delay_5_1;
    io_A_Valid_6_delay_1_56 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_55 <= io_A_Valid_6_delay_1_56;
    io_A_Valid_6_delay_3_54 <= io_A_Valid_6_delay_2_55;
    io_A_Valid_6_delay_4_53 <= io_A_Valid_6_delay_3_54;
    io_A_Valid_6_delay_5_52 <= io_A_Valid_6_delay_4_53;
    io_A_Valid_6_delay_6_51 <= io_A_Valid_6_delay_5_52;
    io_A_Valid_6_delay_7_50 <= io_A_Valid_6_delay_6_51;
    io_A_Valid_6_delay_8_49 <= io_A_Valid_6_delay_7_50;
    io_A_Valid_6_delay_9_48 <= io_A_Valid_6_delay_8_49;
    io_A_Valid_6_delay_10_47 <= io_A_Valid_6_delay_9_48;
    io_A_Valid_6_delay_11_46 <= io_A_Valid_6_delay_10_47;
    io_A_Valid_6_delay_12_45 <= io_A_Valid_6_delay_11_46;
    io_A_Valid_6_delay_13_44 <= io_A_Valid_6_delay_12_45;
    io_A_Valid_6_delay_14_43 <= io_A_Valid_6_delay_13_44;
    io_A_Valid_6_delay_15_42 <= io_A_Valid_6_delay_14_43;
    io_A_Valid_6_delay_16_41 <= io_A_Valid_6_delay_15_42;
    io_A_Valid_6_delay_17_40 <= io_A_Valid_6_delay_16_41;
    io_A_Valid_6_delay_18_39 <= io_A_Valid_6_delay_17_40;
    io_A_Valid_6_delay_19_38 <= io_A_Valid_6_delay_18_39;
    io_A_Valid_6_delay_20_37 <= io_A_Valid_6_delay_19_38;
    io_A_Valid_6_delay_21_36 <= io_A_Valid_6_delay_20_37;
    io_A_Valid_6_delay_22_35 <= io_A_Valid_6_delay_21_36;
    io_A_Valid_6_delay_23_34 <= io_A_Valid_6_delay_22_35;
    io_A_Valid_6_delay_24_33 <= io_A_Valid_6_delay_23_34;
    io_A_Valid_6_delay_25_32 <= io_A_Valid_6_delay_24_33;
    io_A_Valid_6_delay_26_31 <= io_A_Valid_6_delay_25_32;
    io_A_Valid_6_delay_27_30 <= io_A_Valid_6_delay_26_31;
    io_A_Valid_6_delay_28_29 <= io_A_Valid_6_delay_27_30;
    io_A_Valid_6_delay_29_28 <= io_A_Valid_6_delay_28_29;
    io_A_Valid_6_delay_30_27 <= io_A_Valid_6_delay_29_28;
    io_A_Valid_6_delay_31_26 <= io_A_Valid_6_delay_30_27;
    io_A_Valid_6_delay_32_25 <= io_A_Valid_6_delay_31_26;
    io_A_Valid_6_delay_33_24 <= io_A_Valid_6_delay_32_25;
    io_A_Valid_6_delay_34_23 <= io_A_Valid_6_delay_33_24;
    io_A_Valid_6_delay_35_22 <= io_A_Valid_6_delay_34_23;
    io_A_Valid_6_delay_36_21 <= io_A_Valid_6_delay_35_22;
    io_A_Valid_6_delay_37_20 <= io_A_Valid_6_delay_36_21;
    io_A_Valid_6_delay_38_19 <= io_A_Valid_6_delay_37_20;
    io_A_Valid_6_delay_39_18 <= io_A_Valid_6_delay_38_19;
    io_A_Valid_6_delay_40_17 <= io_A_Valid_6_delay_39_18;
    io_A_Valid_6_delay_41_16 <= io_A_Valid_6_delay_40_17;
    io_A_Valid_6_delay_42_15 <= io_A_Valid_6_delay_41_16;
    io_A_Valid_6_delay_43_14 <= io_A_Valid_6_delay_42_15;
    io_A_Valid_6_delay_44_13 <= io_A_Valid_6_delay_43_14;
    io_A_Valid_6_delay_45_12 <= io_A_Valid_6_delay_44_13;
    io_A_Valid_6_delay_46_11 <= io_A_Valid_6_delay_45_12;
    io_A_Valid_6_delay_47_10 <= io_A_Valid_6_delay_46_11;
    io_A_Valid_6_delay_48_9 <= io_A_Valid_6_delay_47_10;
    io_A_Valid_6_delay_49_8 <= io_A_Valid_6_delay_48_9;
    io_A_Valid_6_delay_50_7 <= io_A_Valid_6_delay_49_8;
    io_A_Valid_6_delay_51_6 <= io_A_Valid_6_delay_50_7;
    io_A_Valid_6_delay_52_5 <= io_A_Valid_6_delay_51_6;
    io_A_Valid_6_delay_53_4 <= io_A_Valid_6_delay_52_5;
    io_A_Valid_6_delay_54_3 <= io_A_Valid_6_delay_53_4;
    io_A_Valid_6_delay_55_2 <= io_A_Valid_6_delay_54_3;
    io_A_Valid_6_delay_56_1 <= io_A_Valid_6_delay_55_2;
    io_A_Valid_6_delay_57 <= io_A_Valid_6_delay_56_1;
    io_B_Valid_57_delay_1_5 <= io_B_Valid_57;
    io_B_Valid_57_delay_2_4 <= io_B_Valid_57_delay_1_5;
    io_B_Valid_57_delay_3_3 <= io_B_Valid_57_delay_2_4;
    io_B_Valid_57_delay_4_2 <= io_B_Valid_57_delay_3_3;
    io_B_Valid_57_delay_5_1 <= io_B_Valid_57_delay_4_2;
    io_B_Valid_57_delay_6 <= io_B_Valid_57_delay_5_1;
    io_A_Valid_6_delay_1_57 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_56 <= io_A_Valid_6_delay_1_57;
    io_A_Valid_6_delay_3_55 <= io_A_Valid_6_delay_2_56;
    io_A_Valid_6_delay_4_54 <= io_A_Valid_6_delay_3_55;
    io_A_Valid_6_delay_5_53 <= io_A_Valid_6_delay_4_54;
    io_A_Valid_6_delay_6_52 <= io_A_Valid_6_delay_5_53;
    io_A_Valid_6_delay_7_51 <= io_A_Valid_6_delay_6_52;
    io_A_Valid_6_delay_8_50 <= io_A_Valid_6_delay_7_51;
    io_A_Valid_6_delay_9_49 <= io_A_Valid_6_delay_8_50;
    io_A_Valid_6_delay_10_48 <= io_A_Valid_6_delay_9_49;
    io_A_Valid_6_delay_11_47 <= io_A_Valid_6_delay_10_48;
    io_A_Valid_6_delay_12_46 <= io_A_Valid_6_delay_11_47;
    io_A_Valid_6_delay_13_45 <= io_A_Valid_6_delay_12_46;
    io_A_Valid_6_delay_14_44 <= io_A_Valid_6_delay_13_45;
    io_A_Valid_6_delay_15_43 <= io_A_Valid_6_delay_14_44;
    io_A_Valid_6_delay_16_42 <= io_A_Valid_6_delay_15_43;
    io_A_Valid_6_delay_17_41 <= io_A_Valid_6_delay_16_42;
    io_A_Valid_6_delay_18_40 <= io_A_Valid_6_delay_17_41;
    io_A_Valid_6_delay_19_39 <= io_A_Valid_6_delay_18_40;
    io_A_Valid_6_delay_20_38 <= io_A_Valid_6_delay_19_39;
    io_A_Valid_6_delay_21_37 <= io_A_Valid_6_delay_20_38;
    io_A_Valid_6_delay_22_36 <= io_A_Valid_6_delay_21_37;
    io_A_Valid_6_delay_23_35 <= io_A_Valid_6_delay_22_36;
    io_A_Valid_6_delay_24_34 <= io_A_Valid_6_delay_23_35;
    io_A_Valid_6_delay_25_33 <= io_A_Valid_6_delay_24_34;
    io_A_Valid_6_delay_26_32 <= io_A_Valid_6_delay_25_33;
    io_A_Valid_6_delay_27_31 <= io_A_Valid_6_delay_26_32;
    io_A_Valid_6_delay_28_30 <= io_A_Valid_6_delay_27_31;
    io_A_Valid_6_delay_29_29 <= io_A_Valid_6_delay_28_30;
    io_A_Valid_6_delay_30_28 <= io_A_Valid_6_delay_29_29;
    io_A_Valid_6_delay_31_27 <= io_A_Valid_6_delay_30_28;
    io_A_Valid_6_delay_32_26 <= io_A_Valid_6_delay_31_27;
    io_A_Valid_6_delay_33_25 <= io_A_Valid_6_delay_32_26;
    io_A_Valid_6_delay_34_24 <= io_A_Valid_6_delay_33_25;
    io_A_Valid_6_delay_35_23 <= io_A_Valid_6_delay_34_24;
    io_A_Valid_6_delay_36_22 <= io_A_Valid_6_delay_35_23;
    io_A_Valid_6_delay_37_21 <= io_A_Valid_6_delay_36_22;
    io_A_Valid_6_delay_38_20 <= io_A_Valid_6_delay_37_21;
    io_A_Valid_6_delay_39_19 <= io_A_Valid_6_delay_38_20;
    io_A_Valid_6_delay_40_18 <= io_A_Valid_6_delay_39_19;
    io_A_Valid_6_delay_41_17 <= io_A_Valid_6_delay_40_18;
    io_A_Valid_6_delay_42_16 <= io_A_Valid_6_delay_41_17;
    io_A_Valid_6_delay_43_15 <= io_A_Valid_6_delay_42_16;
    io_A_Valid_6_delay_44_14 <= io_A_Valid_6_delay_43_15;
    io_A_Valid_6_delay_45_13 <= io_A_Valid_6_delay_44_14;
    io_A_Valid_6_delay_46_12 <= io_A_Valid_6_delay_45_13;
    io_A_Valid_6_delay_47_11 <= io_A_Valid_6_delay_46_12;
    io_A_Valid_6_delay_48_10 <= io_A_Valid_6_delay_47_11;
    io_A_Valid_6_delay_49_9 <= io_A_Valid_6_delay_48_10;
    io_A_Valid_6_delay_50_8 <= io_A_Valid_6_delay_49_9;
    io_A_Valid_6_delay_51_7 <= io_A_Valid_6_delay_50_8;
    io_A_Valid_6_delay_52_6 <= io_A_Valid_6_delay_51_7;
    io_A_Valid_6_delay_53_5 <= io_A_Valid_6_delay_52_6;
    io_A_Valid_6_delay_54_4 <= io_A_Valid_6_delay_53_5;
    io_A_Valid_6_delay_55_3 <= io_A_Valid_6_delay_54_4;
    io_A_Valid_6_delay_56_2 <= io_A_Valid_6_delay_55_3;
    io_A_Valid_6_delay_57_1 <= io_A_Valid_6_delay_56_2;
    io_A_Valid_6_delay_58 <= io_A_Valid_6_delay_57_1;
    io_B_Valid_58_delay_1_5 <= io_B_Valid_58;
    io_B_Valid_58_delay_2_4 <= io_B_Valid_58_delay_1_5;
    io_B_Valid_58_delay_3_3 <= io_B_Valid_58_delay_2_4;
    io_B_Valid_58_delay_4_2 <= io_B_Valid_58_delay_3_3;
    io_B_Valid_58_delay_5_1 <= io_B_Valid_58_delay_4_2;
    io_B_Valid_58_delay_6 <= io_B_Valid_58_delay_5_1;
    io_A_Valid_6_delay_1_58 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_57 <= io_A_Valid_6_delay_1_58;
    io_A_Valid_6_delay_3_56 <= io_A_Valid_6_delay_2_57;
    io_A_Valid_6_delay_4_55 <= io_A_Valid_6_delay_3_56;
    io_A_Valid_6_delay_5_54 <= io_A_Valid_6_delay_4_55;
    io_A_Valid_6_delay_6_53 <= io_A_Valid_6_delay_5_54;
    io_A_Valid_6_delay_7_52 <= io_A_Valid_6_delay_6_53;
    io_A_Valid_6_delay_8_51 <= io_A_Valid_6_delay_7_52;
    io_A_Valid_6_delay_9_50 <= io_A_Valid_6_delay_8_51;
    io_A_Valid_6_delay_10_49 <= io_A_Valid_6_delay_9_50;
    io_A_Valid_6_delay_11_48 <= io_A_Valid_6_delay_10_49;
    io_A_Valid_6_delay_12_47 <= io_A_Valid_6_delay_11_48;
    io_A_Valid_6_delay_13_46 <= io_A_Valid_6_delay_12_47;
    io_A_Valid_6_delay_14_45 <= io_A_Valid_6_delay_13_46;
    io_A_Valid_6_delay_15_44 <= io_A_Valid_6_delay_14_45;
    io_A_Valid_6_delay_16_43 <= io_A_Valid_6_delay_15_44;
    io_A_Valid_6_delay_17_42 <= io_A_Valid_6_delay_16_43;
    io_A_Valid_6_delay_18_41 <= io_A_Valid_6_delay_17_42;
    io_A_Valid_6_delay_19_40 <= io_A_Valid_6_delay_18_41;
    io_A_Valid_6_delay_20_39 <= io_A_Valid_6_delay_19_40;
    io_A_Valid_6_delay_21_38 <= io_A_Valid_6_delay_20_39;
    io_A_Valid_6_delay_22_37 <= io_A_Valid_6_delay_21_38;
    io_A_Valid_6_delay_23_36 <= io_A_Valid_6_delay_22_37;
    io_A_Valid_6_delay_24_35 <= io_A_Valid_6_delay_23_36;
    io_A_Valid_6_delay_25_34 <= io_A_Valid_6_delay_24_35;
    io_A_Valid_6_delay_26_33 <= io_A_Valid_6_delay_25_34;
    io_A_Valid_6_delay_27_32 <= io_A_Valid_6_delay_26_33;
    io_A_Valid_6_delay_28_31 <= io_A_Valid_6_delay_27_32;
    io_A_Valid_6_delay_29_30 <= io_A_Valid_6_delay_28_31;
    io_A_Valid_6_delay_30_29 <= io_A_Valid_6_delay_29_30;
    io_A_Valid_6_delay_31_28 <= io_A_Valid_6_delay_30_29;
    io_A_Valid_6_delay_32_27 <= io_A_Valid_6_delay_31_28;
    io_A_Valid_6_delay_33_26 <= io_A_Valid_6_delay_32_27;
    io_A_Valid_6_delay_34_25 <= io_A_Valid_6_delay_33_26;
    io_A_Valid_6_delay_35_24 <= io_A_Valid_6_delay_34_25;
    io_A_Valid_6_delay_36_23 <= io_A_Valid_6_delay_35_24;
    io_A_Valid_6_delay_37_22 <= io_A_Valid_6_delay_36_23;
    io_A_Valid_6_delay_38_21 <= io_A_Valid_6_delay_37_22;
    io_A_Valid_6_delay_39_20 <= io_A_Valid_6_delay_38_21;
    io_A_Valid_6_delay_40_19 <= io_A_Valid_6_delay_39_20;
    io_A_Valid_6_delay_41_18 <= io_A_Valid_6_delay_40_19;
    io_A_Valid_6_delay_42_17 <= io_A_Valid_6_delay_41_18;
    io_A_Valid_6_delay_43_16 <= io_A_Valid_6_delay_42_17;
    io_A_Valid_6_delay_44_15 <= io_A_Valid_6_delay_43_16;
    io_A_Valid_6_delay_45_14 <= io_A_Valid_6_delay_44_15;
    io_A_Valid_6_delay_46_13 <= io_A_Valid_6_delay_45_14;
    io_A_Valid_6_delay_47_12 <= io_A_Valid_6_delay_46_13;
    io_A_Valid_6_delay_48_11 <= io_A_Valid_6_delay_47_12;
    io_A_Valid_6_delay_49_10 <= io_A_Valid_6_delay_48_11;
    io_A_Valid_6_delay_50_9 <= io_A_Valid_6_delay_49_10;
    io_A_Valid_6_delay_51_8 <= io_A_Valid_6_delay_50_9;
    io_A_Valid_6_delay_52_7 <= io_A_Valid_6_delay_51_8;
    io_A_Valid_6_delay_53_6 <= io_A_Valid_6_delay_52_7;
    io_A_Valid_6_delay_54_5 <= io_A_Valid_6_delay_53_6;
    io_A_Valid_6_delay_55_4 <= io_A_Valid_6_delay_54_5;
    io_A_Valid_6_delay_56_3 <= io_A_Valid_6_delay_55_4;
    io_A_Valid_6_delay_57_2 <= io_A_Valid_6_delay_56_3;
    io_A_Valid_6_delay_58_1 <= io_A_Valid_6_delay_57_2;
    io_A_Valid_6_delay_59 <= io_A_Valid_6_delay_58_1;
    io_B_Valid_59_delay_1_5 <= io_B_Valid_59;
    io_B_Valid_59_delay_2_4 <= io_B_Valid_59_delay_1_5;
    io_B_Valid_59_delay_3_3 <= io_B_Valid_59_delay_2_4;
    io_B_Valid_59_delay_4_2 <= io_B_Valid_59_delay_3_3;
    io_B_Valid_59_delay_5_1 <= io_B_Valid_59_delay_4_2;
    io_B_Valid_59_delay_6 <= io_B_Valid_59_delay_5_1;
    io_A_Valid_6_delay_1_59 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_58 <= io_A_Valid_6_delay_1_59;
    io_A_Valid_6_delay_3_57 <= io_A_Valid_6_delay_2_58;
    io_A_Valid_6_delay_4_56 <= io_A_Valid_6_delay_3_57;
    io_A_Valid_6_delay_5_55 <= io_A_Valid_6_delay_4_56;
    io_A_Valid_6_delay_6_54 <= io_A_Valid_6_delay_5_55;
    io_A_Valid_6_delay_7_53 <= io_A_Valid_6_delay_6_54;
    io_A_Valid_6_delay_8_52 <= io_A_Valid_6_delay_7_53;
    io_A_Valid_6_delay_9_51 <= io_A_Valid_6_delay_8_52;
    io_A_Valid_6_delay_10_50 <= io_A_Valid_6_delay_9_51;
    io_A_Valid_6_delay_11_49 <= io_A_Valid_6_delay_10_50;
    io_A_Valid_6_delay_12_48 <= io_A_Valid_6_delay_11_49;
    io_A_Valid_6_delay_13_47 <= io_A_Valid_6_delay_12_48;
    io_A_Valid_6_delay_14_46 <= io_A_Valid_6_delay_13_47;
    io_A_Valid_6_delay_15_45 <= io_A_Valid_6_delay_14_46;
    io_A_Valid_6_delay_16_44 <= io_A_Valid_6_delay_15_45;
    io_A_Valid_6_delay_17_43 <= io_A_Valid_6_delay_16_44;
    io_A_Valid_6_delay_18_42 <= io_A_Valid_6_delay_17_43;
    io_A_Valid_6_delay_19_41 <= io_A_Valid_6_delay_18_42;
    io_A_Valid_6_delay_20_40 <= io_A_Valid_6_delay_19_41;
    io_A_Valid_6_delay_21_39 <= io_A_Valid_6_delay_20_40;
    io_A_Valid_6_delay_22_38 <= io_A_Valid_6_delay_21_39;
    io_A_Valid_6_delay_23_37 <= io_A_Valid_6_delay_22_38;
    io_A_Valid_6_delay_24_36 <= io_A_Valid_6_delay_23_37;
    io_A_Valid_6_delay_25_35 <= io_A_Valid_6_delay_24_36;
    io_A_Valid_6_delay_26_34 <= io_A_Valid_6_delay_25_35;
    io_A_Valid_6_delay_27_33 <= io_A_Valid_6_delay_26_34;
    io_A_Valid_6_delay_28_32 <= io_A_Valid_6_delay_27_33;
    io_A_Valid_6_delay_29_31 <= io_A_Valid_6_delay_28_32;
    io_A_Valid_6_delay_30_30 <= io_A_Valid_6_delay_29_31;
    io_A_Valid_6_delay_31_29 <= io_A_Valid_6_delay_30_30;
    io_A_Valid_6_delay_32_28 <= io_A_Valid_6_delay_31_29;
    io_A_Valid_6_delay_33_27 <= io_A_Valid_6_delay_32_28;
    io_A_Valid_6_delay_34_26 <= io_A_Valid_6_delay_33_27;
    io_A_Valid_6_delay_35_25 <= io_A_Valid_6_delay_34_26;
    io_A_Valid_6_delay_36_24 <= io_A_Valid_6_delay_35_25;
    io_A_Valid_6_delay_37_23 <= io_A_Valid_6_delay_36_24;
    io_A_Valid_6_delay_38_22 <= io_A_Valid_6_delay_37_23;
    io_A_Valid_6_delay_39_21 <= io_A_Valid_6_delay_38_22;
    io_A_Valid_6_delay_40_20 <= io_A_Valid_6_delay_39_21;
    io_A_Valid_6_delay_41_19 <= io_A_Valid_6_delay_40_20;
    io_A_Valid_6_delay_42_18 <= io_A_Valid_6_delay_41_19;
    io_A_Valid_6_delay_43_17 <= io_A_Valid_6_delay_42_18;
    io_A_Valid_6_delay_44_16 <= io_A_Valid_6_delay_43_17;
    io_A_Valid_6_delay_45_15 <= io_A_Valid_6_delay_44_16;
    io_A_Valid_6_delay_46_14 <= io_A_Valid_6_delay_45_15;
    io_A_Valid_6_delay_47_13 <= io_A_Valid_6_delay_46_14;
    io_A_Valid_6_delay_48_12 <= io_A_Valid_6_delay_47_13;
    io_A_Valid_6_delay_49_11 <= io_A_Valid_6_delay_48_12;
    io_A_Valid_6_delay_50_10 <= io_A_Valid_6_delay_49_11;
    io_A_Valid_6_delay_51_9 <= io_A_Valid_6_delay_50_10;
    io_A_Valid_6_delay_52_8 <= io_A_Valid_6_delay_51_9;
    io_A_Valid_6_delay_53_7 <= io_A_Valid_6_delay_52_8;
    io_A_Valid_6_delay_54_6 <= io_A_Valid_6_delay_53_7;
    io_A_Valid_6_delay_55_5 <= io_A_Valid_6_delay_54_6;
    io_A_Valid_6_delay_56_4 <= io_A_Valid_6_delay_55_5;
    io_A_Valid_6_delay_57_3 <= io_A_Valid_6_delay_56_4;
    io_A_Valid_6_delay_58_2 <= io_A_Valid_6_delay_57_3;
    io_A_Valid_6_delay_59_1 <= io_A_Valid_6_delay_58_2;
    io_A_Valid_6_delay_60 <= io_A_Valid_6_delay_59_1;
    io_B_Valid_60_delay_1_5 <= io_B_Valid_60;
    io_B_Valid_60_delay_2_4 <= io_B_Valid_60_delay_1_5;
    io_B_Valid_60_delay_3_3 <= io_B_Valid_60_delay_2_4;
    io_B_Valid_60_delay_4_2 <= io_B_Valid_60_delay_3_3;
    io_B_Valid_60_delay_5_1 <= io_B_Valid_60_delay_4_2;
    io_B_Valid_60_delay_6 <= io_B_Valid_60_delay_5_1;
    io_A_Valid_6_delay_1_60 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_59 <= io_A_Valid_6_delay_1_60;
    io_A_Valid_6_delay_3_58 <= io_A_Valid_6_delay_2_59;
    io_A_Valid_6_delay_4_57 <= io_A_Valid_6_delay_3_58;
    io_A_Valid_6_delay_5_56 <= io_A_Valid_6_delay_4_57;
    io_A_Valid_6_delay_6_55 <= io_A_Valid_6_delay_5_56;
    io_A_Valid_6_delay_7_54 <= io_A_Valid_6_delay_6_55;
    io_A_Valid_6_delay_8_53 <= io_A_Valid_6_delay_7_54;
    io_A_Valid_6_delay_9_52 <= io_A_Valid_6_delay_8_53;
    io_A_Valid_6_delay_10_51 <= io_A_Valid_6_delay_9_52;
    io_A_Valid_6_delay_11_50 <= io_A_Valid_6_delay_10_51;
    io_A_Valid_6_delay_12_49 <= io_A_Valid_6_delay_11_50;
    io_A_Valid_6_delay_13_48 <= io_A_Valid_6_delay_12_49;
    io_A_Valid_6_delay_14_47 <= io_A_Valid_6_delay_13_48;
    io_A_Valid_6_delay_15_46 <= io_A_Valid_6_delay_14_47;
    io_A_Valid_6_delay_16_45 <= io_A_Valid_6_delay_15_46;
    io_A_Valid_6_delay_17_44 <= io_A_Valid_6_delay_16_45;
    io_A_Valid_6_delay_18_43 <= io_A_Valid_6_delay_17_44;
    io_A_Valid_6_delay_19_42 <= io_A_Valid_6_delay_18_43;
    io_A_Valid_6_delay_20_41 <= io_A_Valid_6_delay_19_42;
    io_A_Valid_6_delay_21_40 <= io_A_Valid_6_delay_20_41;
    io_A_Valid_6_delay_22_39 <= io_A_Valid_6_delay_21_40;
    io_A_Valid_6_delay_23_38 <= io_A_Valid_6_delay_22_39;
    io_A_Valid_6_delay_24_37 <= io_A_Valid_6_delay_23_38;
    io_A_Valid_6_delay_25_36 <= io_A_Valid_6_delay_24_37;
    io_A_Valid_6_delay_26_35 <= io_A_Valid_6_delay_25_36;
    io_A_Valid_6_delay_27_34 <= io_A_Valid_6_delay_26_35;
    io_A_Valid_6_delay_28_33 <= io_A_Valid_6_delay_27_34;
    io_A_Valid_6_delay_29_32 <= io_A_Valid_6_delay_28_33;
    io_A_Valid_6_delay_30_31 <= io_A_Valid_6_delay_29_32;
    io_A_Valid_6_delay_31_30 <= io_A_Valid_6_delay_30_31;
    io_A_Valid_6_delay_32_29 <= io_A_Valid_6_delay_31_30;
    io_A_Valid_6_delay_33_28 <= io_A_Valid_6_delay_32_29;
    io_A_Valid_6_delay_34_27 <= io_A_Valid_6_delay_33_28;
    io_A_Valid_6_delay_35_26 <= io_A_Valid_6_delay_34_27;
    io_A_Valid_6_delay_36_25 <= io_A_Valid_6_delay_35_26;
    io_A_Valid_6_delay_37_24 <= io_A_Valid_6_delay_36_25;
    io_A_Valid_6_delay_38_23 <= io_A_Valid_6_delay_37_24;
    io_A_Valid_6_delay_39_22 <= io_A_Valid_6_delay_38_23;
    io_A_Valid_6_delay_40_21 <= io_A_Valid_6_delay_39_22;
    io_A_Valid_6_delay_41_20 <= io_A_Valid_6_delay_40_21;
    io_A_Valid_6_delay_42_19 <= io_A_Valid_6_delay_41_20;
    io_A_Valid_6_delay_43_18 <= io_A_Valid_6_delay_42_19;
    io_A_Valid_6_delay_44_17 <= io_A_Valid_6_delay_43_18;
    io_A_Valid_6_delay_45_16 <= io_A_Valid_6_delay_44_17;
    io_A_Valid_6_delay_46_15 <= io_A_Valid_6_delay_45_16;
    io_A_Valid_6_delay_47_14 <= io_A_Valid_6_delay_46_15;
    io_A_Valid_6_delay_48_13 <= io_A_Valid_6_delay_47_14;
    io_A_Valid_6_delay_49_12 <= io_A_Valid_6_delay_48_13;
    io_A_Valid_6_delay_50_11 <= io_A_Valid_6_delay_49_12;
    io_A_Valid_6_delay_51_10 <= io_A_Valid_6_delay_50_11;
    io_A_Valid_6_delay_52_9 <= io_A_Valid_6_delay_51_10;
    io_A_Valid_6_delay_53_8 <= io_A_Valid_6_delay_52_9;
    io_A_Valid_6_delay_54_7 <= io_A_Valid_6_delay_53_8;
    io_A_Valid_6_delay_55_6 <= io_A_Valid_6_delay_54_7;
    io_A_Valid_6_delay_56_5 <= io_A_Valid_6_delay_55_6;
    io_A_Valid_6_delay_57_4 <= io_A_Valid_6_delay_56_5;
    io_A_Valid_6_delay_58_3 <= io_A_Valid_6_delay_57_4;
    io_A_Valid_6_delay_59_2 <= io_A_Valid_6_delay_58_3;
    io_A_Valid_6_delay_60_1 <= io_A_Valid_6_delay_59_2;
    io_A_Valid_6_delay_61 <= io_A_Valid_6_delay_60_1;
    io_B_Valid_61_delay_1_5 <= io_B_Valid_61;
    io_B_Valid_61_delay_2_4 <= io_B_Valid_61_delay_1_5;
    io_B_Valid_61_delay_3_3 <= io_B_Valid_61_delay_2_4;
    io_B_Valid_61_delay_4_2 <= io_B_Valid_61_delay_3_3;
    io_B_Valid_61_delay_5_1 <= io_B_Valid_61_delay_4_2;
    io_B_Valid_61_delay_6 <= io_B_Valid_61_delay_5_1;
    io_A_Valid_6_delay_1_61 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_60 <= io_A_Valid_6_delay_1_61;
    io_A_Valid_6_delay_3_59 <= io_A_Valid_6_delay_2_60;
    io_A_Valid_6_delay_4_58 <= io_A_Valid_6_delay_3_59;
    io_A_Valid_6_delay_5_57 <= io_A_Valid_6_delay_4_58;
    io_A_Valid_6_delay_6_56 <= io_A_Valid_6_delay_5_57;
    io_A_Valid_6_delay_7_55 <= io_A_Valid_6_delay_6_56;
    io_A_Valid_6_delay_8_54 <= io_A_Valid_6_delay_7_55;
    io_A_Valid_6_delay_9_53 <= io_A_Valid_6_delay_8_54;
    io_A_Valid_6_delay_10_52 <= io_A_Valid_6_delay_9_53;
    io_A_Valid_6_delay_11_51 <= io_A_Valid_6_delay_10_52;
    io_A_Valid_6_delay_12_50 <= io_A_Valid_6_delay_11_51;
    io_A_Valid_6_delay_13_49 <= io_A_Valid_6_delay_12_50;
    io_A_Valid_6_delay_14_48 <= io_A_Valid_6_delay_13_49;
    io_A_Valid_6_delay_15_47 <= io_A_Valid_6_delay_14_48;
    io_A_Valid_6_delay_16_46 <= io_A_Valid_6_delay_15_47;
    io_A_Valid_6_delay_17_45 <= io_A_Valid_6_delay_16_46;
    io_A_Valid_6_delay_18_44 <= io_A_Valid_6_delay_17_45;
    io_A_Valid_6_delay_19_43 <= io_A_Valid_6_delay_18_44;
    io_A_Valid_6_delay_20_42 <= io_A_Valid_6_delay_19_43;
    io_A_Valid_6_delay_21_41 <= io_A_Valid_6_delay_20_42;
    io_A_Valid_6_delay_22_40 <= io_A_Valid_6_delay_21_41;
    io_A_Valid_6_delay_23_39 <= io_A_Valid_6_delay_22_40;
    io_A_Valid_6_delay_24_38 <= io_A_Valid_6_delay_23_39;
    io_A_Valid_6_delay_25_37 <= io_A_Valid_6_delay_24_38;
    io_A_Valid_6_delay_26_36 <= io_A_Valid_6_delay_25_37;
    io_A_Valid_6_delay_27_35 <= io_A_Valid_6_delay_26_36;
    io_A_Valid_6_delay_28_34 <= io_A_Valid_6_delay_27_35;
    io_A_Valid_6_delay_29_33 <= io_A_Valid_6_delay_28_34;
    io_A_Valid_6_delay_30_32 <= io_A_Valid_6_delay_29_33;
    io_A_Valid_6_delay_31_31 <= io_A_Valid_6_delay_30_32;
    io_A_Valid_6_delay_32_30 <= io_A_Valid_6_delay_31_31;
    io_A_Valid_6_delay_33_29 <= io_A_Valid_6_delay_32_30;
    io_A_Valid_6_delay_34_28 <= io_A_Valid_6_delay_33_29;
    io_A_Valid_6_delay_35_27 <= io_A_Valid_6_delay_34_28;
    io_A_Valid_6_delay_36_26 <= io_A_Valid_6_delay_35_27;
    io_A_Valid_6_delay_37_25 <= io_A_Valid_6_delay_36_26;
    io_A_Valid_6_delay_38_24 <= io_A_Valid_6_delay_37_25;
    io_A_Valid_6_delay_39_23 <= io_A_Valid_6_delay_38_24;
    io_A_Valid_6_delay_40_22 <= io_A_Valid_6_delay_39_23;
    io_A_Valid_6_delay_41_21 <= io_A_Valid_6_delay_40_22;
    io_A_Valid_6_delay_42_20 <= io_A_Valid_6_delay_41_21;
    io_A_Valid_6_delay_43_19 <= io_A_Valid_6_delay_42_20;
    io_A_Valid_6_delay_44_18 <= io_A_Valid_6_delay_43_19;
    io_A_Valid_6_delay_45_17 <= io_A_Valid_6_delay_44_18;
    io_A_Valid_6_delay_46_16 <= io_A_Valid_6_delay_45_17;
    io_A_Valid_6_delay_47_15 <= io_A_Valid_6_delay_46_16;
    io_A_Valid_6_delay_48_14 <= io_A_Valid_6_delay_47_15;
    io_A_Valid_6_delay_49_13 <= io_A_Valid_6_delay_48_14;
    io_A_Valid_6_delay_50_12 <= io_A_Valid_6_delay_49_13;
    io_A_Valid_6_delay_51_11 <= io_A_Valid_6_delay_50_12;
    io_A_Valid_6_delay_52_10 <= io_A_Valid_6_delay_51_11;
    io_A_Valid_6_delay_53_9 <= io_A_Valid_6_delay_52_10;
    io_A_Valid_6_delay_54_8 <= io_A_Valid_6_delay_53_9;
    io_A_Valid_6_delay_55_7 <= io_A_Valid_6_delay_54_8;
    io_A_Valid_6_delay_56_6 <= io_A_Valid_6_delay_55_7;
    io_A_Valid_6_delay_57_5 <= io_A_Valid_6_delay_56_6;
    io_A_Valid_6_delay_58_4 <= io_A_Valid_6_delay_57_5;
    io_A_Valid_6_delay_59_3 <= io_A_Valid_6_delay_58_4;
    io_A_Valid_6_delay_60_2 <= io_A_Valid_6_delay_59_3;
    io_A_Valid_6_delay_61_1 <= io_A_Valid_6_delay_60_2;
    io_A_Valid_6_delay_62 <= io_A_Valid_6_delay_61_1;
    io_B_Valid_62_delay_1_5 <= io_B_Valid_62;
    io_B_Valid_62_delay_2_4 <= io_B_Valid_62_delay_1_5;
    io_B_Valid_62_delay_3_3 <= io_B_Valid_62_delay_2_4;
    io_B_Valid_62_delay_4_2 <= io_B_Valid_62_delay_3_3;
    io_B_Valid_62_delay_5_1 <= io_B_Valid_62_delay_4_2;
    io_B_Valid_62_delay_6 <= io_B_Valid_62_delay_5_1;
    io_A_Valid_6_delay_1_62 <= io_A_Valid_6;
    io_A_Valid_6_delay_2_61 <= io_A_Valid_6_delay_1_62;
    io_A_Valid_6_delay_3_60 <= io_A_Valid_6_delay_2_61;
    io_A_Valid_6_delay_4_59 <= io_A_Valid_6_delay_3_60;
    io_A_Valid_6_delay_5_58 <= io_A_Valid_6_delay_4_59;
    io_A_Valid_6_delay_6_57 <= io_A_Valid_6_delay_5_58;
    io_A_Valid_6_delay_7_56 <= io_A_Valid_6_delay_6_57;
    io_A_Valid_6_delay_8_55 <= io_A_Valid_6_delay_7_56;
    io_A_Valid_6_delay_9_54 <= io_A_Valid_6_delay_8_55;
    io_A_Valid_6_delay_10_53 <= io_A_Valid_6_delay_9_54;
    io_A_Valid_6_delay_11_52 <= io_A_Valid_6_delay_10_53;
    io_A_Valid_6_delay_12_51 <= io_A_Valid_6_delay_11_52;
    io_A_Valid_6_delay_13_50 <= io_A_Valid_6_delay_12_51;
    io_A_Valid_6_delay_14_49 <= io_A_Valid_6_delay_13_50;
    io_A_Valid_6_delay_15_48 <= io_A_Valid_6_delay_14_49;
    io_A_Valid_6_delay_16_47 <= io_A_Valid_6_delay_15_48;
    io_A_Valid_6_delay_17_46 <= io_A_Valid_6_delay_16_47;
    io_A_Valid_6_delay_18_45 <= io_A_Valid_6_delay_17_46;
    io_A_Valid_6_delay_19_44 <= io_A_Valid_6_delay_18_45;
    io_A_Valid_6_delay_20_43 <= io_A_Valid_6_delay_19_44;
    io_A_Valid_6_delay_21_42 <= io_A_Valid_6_delay_20_43;
    io_A_Valid_6_delay_22_41 <= io_A_Valid_6_delay_21_42;
    io_A_Valid_6_delay_23_40 <= io_A_Valid_6_delay_22_41;
    io_A_Valid_6_delay_24_39 <= io_A_Valid_6_delay_23_40;
    io_A_Valid_6_delay_25_38 <= io_A_Valid_6_delay_24_39;
    io_A_Valid_6_delay_26_37 <= io_A_Valid_6_delay_25_38;
    io_A_Valid_6_delay_27_36 <= io_A_Valid_6_delay_26_37;
    io_A_Valid_6_delay_28_35 <= io_A_Valid_6_delay_27_36;
    io_A_Valid_6_delay_29_34 <= io_A_Valid_6_delay_28_35;
    io_A_Valid_6_delay_30_33 <= io_A_Valid_6_delay_29_34;
    io_A_Valid_6_delay_31_32 <= io_A_Valid_6_delay_30_33;
    io_A_Valid_6_delay_32_31 <= io_A_Valid_6_delay_31_32;
    io_A_Valid_6_delay_33_30 <= io_A_Valid_6_delay_32_31;
    io_A_Valid_6_delay_34_29 <= io_A_Valid_6_delay_33_30;
    io_A_Valid_6_delay_35_28 <= io_A_Valid_6_delay_34_29;
    io_A_Valid_6_delay_36_27 <= io_A_Valid_6_delay_35_28;
    io_A_Valid_6_delay_37_26 <= io_A_Valid_6_delay_36_27;
    io_A_Valid_6_delay_38_25 <= io_A_Valid_6_delay_37_26;
    io_A_Valid_6_delay_39_24 <= io_A_Valid_6_delay_38_25;
    io_A_Valid_6_delay_40_23 <= io_A_Valid_6_delay_39_24;
    io_A_Valid_6_delay_41_22 <= io_A_Valid_6_delay_40_23;
    io_A_Valid_6_delay_42_21 <= io_A_Valid_6_delay_41_22;
    io_A_Valid_6_delay_43_20 <= io_A_Valid_6_delay_42_21;
    io_A_Valid_6_delay_44_19 <= io_A_Valid_6_delay_43_20;
    io_A_Valid_6_delay_45_18 <= io_A_Valid_6_delay_44_19;
    io_A_Valid_6_delay_46_17 <= io_A_Valid_6_delay_45_18;
    io_A_Valid_6_delay_47_16 <= io_A_Valid_6_delay_46_17;
    io_A_Valid_6_delay_48_15 <= io_A_Valid_6_delay_47_16;
    io_A_Valid_6_delay_49_14 <= io_A_Valid_6_delay_48_15;
    io_A_Valid_6_delay_50_13 <= io_A_Valid_6_delay_49_14;
    io_A_Valid_6_delay_51_12 <= io_A_Valid_6_delay_50_13;
    io_A_Valid_6_delay_52_11 <= io_A_Valid_6_delay_51_12;
    io_A_Valid_6_delay_53_10 <= io_A_Valid_6_delay_52_11;
    io_A_Valid_6_delay_54_9 <= io_A_Valid_6_delay_53_10;
    io_A_Valid_6_delay_55_8 <= io_A_Valid_6_delay_54_9;
    io_A_Valid_6_delay_56_7 <= io_A_Valid_6_delay_55_8;
    io_A_Valid_6_delay_57_6 <= io_A_Valid_6_delay_56_7;
    io_A_Valid_6_delay_58_5 <= io_A_Valid_6_delay_57_6;
    io_A_Valid_6_delay_59_4 <= io_A_Valid_6_delay_58_5;
    io_A_Valid_6_delay_60_3 <= io_A_Valid_6_delay_59_4;
    io_A_Valid_6_delay_61_2 <= io_A_Valid_6_delay_60_3;
    io_A_Valid_6_delay_62_1 <= io_A_Valid_6_delay_61_2;
    io_A_Valid_6_delay_63 <= io_A_Valid_6_delay_62_1;
    io_B_Valid_63_delay_1_5 <= io_B_Valid_63;
    io_B_Valid_63_delay_2_4 <= io_B_Valid_63_delay_1_5;
    io_B_Valid_63_delay_3_3 <= io_B_Valid_63_delay_2_4;
    io_B_Valid_63_delay_4_2 <= io_B_Valid_63_delay_3_3;
    io_B_Valid_63_delay_5_1 <= io_B_Valid_63_delay_4_2;
    io_B_Valid_63_delay_6 <= io_B_Valid_63_delay_5_1;
    io_B_Valid_0_delay_1_6 <= io_B_Valid_0;
    io_B_Valid_0_delay_2_5 <= io_B_Valid_0_delay_1_6;
    io_B_Valid_0_delay_3_4 <= io_B_Valid_0_delay_2_5;
    io_B_Valid_0_delay_4_3 <= io_B_Valid_0_delay_3_4;
    io_B_Valid_0_delay_5_2 <= io_B_Valid_0_delay_4_3;
    io_B_Valid_0_delay_6_1 <= io_B_Valid_0_delay_5_2;
    io_B_Valid_0_delay_7 <= io_B_Valid_0_delay_6_1;
    io_A_Valid_7_delay_1 <= io_A_Valid_7;
    io_B_Valid_1_delay_1_6 <= io_B_Valid_1;
    io_B_Valid_1_delay_2_5 <= io_B_Valid_1_delay_1_6;
    io_B_Valid_1_delay_3_4 <= io_B_Valid_1_delay_2_5;
    io_B_Valid_1_delay_4_3 <= io_B_Valid_1_delay_3_4;
    io_B_Valid_1_delay_5_2 <= io_B_Valid_1_delay_4_3;
    io_B_Valid_1_delay_6_1 <= io_B_Valid_1_delay_5_2;
    io_B_Valid_1_delay_7 <= io_B_Valid_1_delay_6_1;
    io_A_Valid_7_delay_1_1 <= io_A_Valid_7;
    io_A_Valid_7_delay_2 <= io_A_Valid_7_delay_1_1;
    io_B_Valid_2_delay_1_6 <= io_B_Valid_2;
    io_B_Valid_2_delay_2_5 <= io_B_Valid_2_delay_1_6;
    io_B_Valid_2_delay_3_4 <= io_B_Valid_2_delay_2_5;
    io_B_Valid_2_delay_4_3 <= io_B_Valid_2_delay_3_4;
    io_B_Valid_2_delay_5_2 <= io_B_Valid_2_delay_4_3;
    io_B_Valid_2_delay_6_1 <= io_B_Valid_2_delay_5_2;
    io_B_Valid_2_delay_7 <= io_B_Valid_2_delay_6_1;
    io_A_Valid_7_delay_1_2 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_1 <= io_A_Valid_7_delay_1_2;
    io_A_Valid_7_delay_3 <= io_A_Valid_7_delay_2_1;
    io_B_Valid_3_delay_1_6 <= io_B_Valid_3;
    io_B_Valid_3_delay_2_5 <= io_B_Valid_3_delay_1_6;
    io_B_Valid_3_delay_3_4 <= io_B_Valid_3_delay_2_5;
    io_B_Valid_3_delay_4_3 <= io_B_Valid_3_delay_3_4;
    io_B_Valid_3_delay_5_2 <= io_B_Valid_3_delay_4_3;
    io_B_Valid_3_delay_6_1 <= io_B_Valid_3_delay_5_2;
    io_B_Valid_3_delay_7 <= io_B_Valid_3_delay_6_1;
    io_A_Valid_7_delay_1_3 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_2 <= io_A_Valid_7_delay_1_3;
    io_A_Valid_7_delay_3_1 <= io_A_Valid_7_delay_2_2;
    io_A_Valid_7_delay_4 <= io_A_Valid_7_delay_3_1;
    io_B_Valid_4_delay_1_6 <= io_B_Valid_4;
    io_B_Valid_4_delay_2_5 <= io_B_Valid_4_delay_1_6;
    io_B_Valid_4_delay_3_4 <= io_B_Valid_4_delay_2_5;
    io_B_Valid_4_delay_4_3 <= io_B_Valid_4_delay_3_4;
    io_B_Valid_4_delay_5_2 <= io_B_Valid_4_delay_4_3;
    io_B_Valid_4_delay_6_1 <= io_B_Valid_4_delay_5_2;
    io_B_Valid_4_delay_7 <= io_B_Valid_4_delay_6_1;
    io_A_Valid_7_delay_1_4 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_3 <= io_A_Valid_7_delay_1_4;
    io_A_Valid_7_delay_3_2 <= io_A_Valid_7_delay_2_3;
    io_A_Valid_7_delay_4_1 <= io_A_Valid_7_delay_3_2;
    io_A_Valid_7_delay_5 <= io_A_Valid_7_delay_4_1;
    io_B_Valid_5_delay_1_6 <= io_B_Valid_5;
    io_B_Valid_5_delay_2_5 <= io_B_Valid_5_delay_1_6;
    io_B_Valid_5_delay_3_4 <= io_B_Valid_5_delay_2_5;
    io_B_Valid_5_delay_4_3 <= io_B_Valid_5_delay_3_4;
    io_B_Valid_5_delay_5_2 <= io_B_Valid_5_delay_4_3;
    io_B_Valid_5_delay_6_1 <= io_B_Valid_5_delay_5_2;
    io_B_Valid_5_delay_7 <= io_B_Valid_5_delay_6_1;
    io_A_Valid_7_delay_1_5 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_4 <= io_A_Valid_7_delay_1_5;
    io_A_Valid_7_delay_3_3 <= io_A_Valid_7_delay_2_4;
    io_A_Valid_7_delay_4_2 <= io_A_Valid_7_delay_3_3;
    io_A_Valid_7_delay_5_1 <= io_A_Valid_7_delay_4_2;
    io_A_Valid_7_delay_6 <= io_A_Valid_7_delay_5_1;
    io_B_Valid_6_delay_1_6 <= io_B_Valid_6;
    io_B_Valid_6_delay_2_5 <= io_B_Valid_6_delay_1_6;
    io_B_Valid_6_delay_3_4 <= io_B_Valid_6_delay_2_5;
    io_B_Valid_6_delay_4_3 <= io_B_Valid_6_delay_3_4;
    io_B_Valid_6_delay_5_2 <= io_B_Valid_6_delay_4_3;
    io_B_Valid_6_delay_6_1 <= io_B_Valid_6_delay_5_2;
    io_B_Valid_6_delay_7 <= io_B_Valid_6_delay_6_1;
    io_A_Valid_7_delay_1_6 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_5 <= io_A_Valid_7_delay_1_6;
    io_A_Valid_7_delay_3_4 <= io_A_Valid_7_delay_2_5;
    io_A_Valid_7_delay_4_3 <= io_A_Valid_7_delay_3_4;
    io_A_Valid_7_delay_5_2 <= io_A_Valid_7_delay_4_3;
    io_A_Valid_7_delay_6_1 <= io_A_Valid_7_delay_5_2;
    io_A_Valid_7_delay_7 <= io_A_Valid_7_delay_6_1;
    io_B_Valid_7_delay_1_6 <= io_B_Valid_7;
    io_B_Valid_7_delay_2_5 <= io_B_Valid_7_delay_1_6;
    io_B_Valid_7_delay_3_4 <= io_B_Valid_7_delay_2_5;
    io_B_Valid_7_delay_4_3 <= io_B_Valid_7_delay_3_4;
    io_B_Valid_7_delay_5_2 <= io_B_Valid_7_delay_4_3;
    io_B_Valid_7_delay_6_1 <= io_B_Valid_7_delay_5_2;
    io_B_Valid_7_delay_7 <= io_B_Valid_7_delay_6_1;
    io_A_Valid_7_delay_1_7 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_6 <= io_A_Valid_7_delay_1_7;
    io_A_Valid_7_delay_3_5 <= io_A_Valid_7_delay_2_6;
    io_A_Valid_7_delay_4_4 <= io_A_Valid_7_delay_3_5;
    io_A_Valid_7_delay_5_3 <= io_A_Valid_7_delay_4_4;
    io_A_Valid_7_delay_6_2 <= io_A_Valid_7_delay_5_3;
    io_A_Valid_7_delay_7_1 <= io_A_Valid_7_delay_6_2;
    io_A_Valid_7_delay_8 <= io_A_Valid_7_delay_7_1;
    io_B_Valid_8_delay_1_6 <= io_B_Valid_8;
    io_B_Valid_8_delay_2_5 <= io_B_Valid_8_delay_1_6;
    io_B_Valid_8_delay_3_4 <= io_B_Valid_8_delay_2_5;
    io_B_Valid_8_delay_4_3 <= io_B_Valid_8_delay_3_4;
    io_B_Valid_8_delay_5_2 <= io_B_Valid_8_delay_4_3;
    io_B_Valid_8_delay_6_1 <= io_B_Valid_8_delay_5_2;
    io_B_Valid_8_delay_7 <= io_B_Valid_8_delay_6_1;
    io_A_Valid_7_delay_1_8 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_7 <= io_A_Valid_7_delay_1_8;
    io_A_Valid_7_delay_3_6 <= io_A_Valid_7_delay_2_7;
    io_A_Valid_7_delay_4_5 <= io_A_Valid_7_delay_3_6;
    io_A_Valid_7_delay_5_4 <= io_A_Valid_7_delay_4_5;
    io_A_Valid_7_delay_6_3 <= io_A_Valid_7_delay_5_4;
    io_A_Valid_7_delay_7_2 <= io_A_Valid_7_delay_6_3;
    io_A_Valid_7_delay_8_1 <= io_A_Valid_7_delay_7_2;
    io_A_Valid_7_delay_9 <= io_A_Valid_7_delay_8_1;
    io_B_Valid_9_delay_1_6 <= io_B_Valid_9;
    io_B_Valid_9_delay_2_5 <= io_B_Valid_9_delay_1_6;
    io_B_Valid_9_delay_3_4 <= io_B_Valid_9_delay_2_5;
    io_B_Valid_9_delay_4_3 <= io_B_Valid_9_delay_3_4;
    io_B_Valid_9_delay_5_2 <= io_B_Valid_9_delay_4_3;
    io_B_Valid_9_delay_6_1 <= io_B_Valid_9_delay_5_2;
    io_B_Valid_9_delay_7 <= io_B_Valid_9_delay_6_1;
    io_A_Valid_7_delay_1_9 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_8 <= io_A_Valid_7_delay_1_9;
    io_A_Valid_7_delay_3_7 <= io_A_Valid_7_delay_2_8;
    io_A_Valid_7_delay_4_6 <= io_A_Valid_7_delay_3_7;
    io_A_Valid_7_delay_5_5 <= io_A_Valid_7_delay_4_6;
    io_A_Valid_7_delay_6_4 <= io_A_Valid_7_delay_5_5;
    io_A_Valid_7_delay_7_3 <= io_A_Valid_7_delay_6_4;
    io_A_Valid_7_delay_8_2 <= io_A_Valid_7_delay_7_3;
    io_A_Valid_7_delay_9_1 <= io_A_Valid_7_delay_8_2;
    io_A_Valid_7_delay_10 <= io_A_Valid_7_delay_9_1;
    io_B_Valid_10_delay_1_6 <= io_B_Valid_10;
    io_B_Valid_10_delay_2_5 <= io_B_Valid_10_delay_1_6;
    io_B_Valid_10_delay_3_4 <= io_B_Valid_10_delay_2_5;
    io_B_Valid_10_delay_4_3 <= io_B_Valid_10_delay_3_4;
    io_B_Valid_10_delay_5_2 <= io_B_Valid_10_delay_4_3;
    io_B_Valid_10_delay_6_1 <= io_B_Valid_10_delay_5_2;
    io_B_Valid_10_delay_7 <= io_B_Valid_10_delay_6_1;
    io_A_Valid_7_delay_1_10 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_9 <= io_A_Valid_7_delay_1_10;
    io_A_Valid_7_delay_3_8 <= io_A_Valid_7_delay_2_9;
    io_A_Valid_7_delay_4_7 <= io_A_Valid_7_delay_3_8;
    io_A_Valid_7_delay_5_6 <= io_A_Valid_7_delay_4_7;
    io_A_Valid_7_delay_6_5 <= io_A_Valid_7_delay_5_6;
    io_A_Valid_7_delay_7_4 <= io_A_Valid_7_delay_6_5;
    io_A_Valid_7_delay_8_3 <= io_A_Valid_7_delay_7_4;
    io_A_Valid_7_delay_9_2 <= io_A_Valid_7_delay_8_3;
    io_A_Valid_7_delay_10_1 <= io_A_Valid_7_delay_9_2;
    io_A_Valid_7_delay_11 <= io_A_Valid_7_delay_10_1;
    io_B_Valid_11_delay_1_6 <= io_B_Valid_11;
    io_B_Valid_11_delay_2_5 <= io_B_Valid_11_delay_1_6;
    io_B_Valid_11_delay_3_4 <= io_B_Valid_11_delay_2_5;
    io_B_Valid_11_delay_4_3 <= io_B_Valid_11_delay_3_4;
    io_B_Valid_11_delay_5_2 <= io_B_Valid_11_delay_4_3;
    io_B_Valid_11_delay_6_1 <= io_B_Valid_11_delay_5_2;
    io_B_Valid_11_delay_7 <= io_B_Valid_11_delay_6_1;
    io_A_Valid_7_delay_1_11 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_10 <= io_A_Valid_7_delay_1_11;
    io_A_Valid_7_delay_3_9 <= io_A_Valid_7_delay_2_10;
    io_A_Valid_7_delay_4_8 <= io_A_Valid_7_delay_3_9;
    io_A_Valid_7_delay_5_7 <= io_A_Valid_7_delay_4_8;
    io_A_Valid_7_delay_6_6 <= io_A_Valid_7_delay_5_7;
    io_A_Valid_7_delay_7_5 <= io_A_Valid_7_delay_6_6;
    io_A_Valid_7_delay_8_4 <= io_A_Valid_7_delay_7_5;
    io_A_Valid_7_delay_9_3 <= io_A_Valid_7_delay_8_4;
    io_A_Valid_7_delay_10_2 <= io_A_Valid_7_delay_9_3;
    io_A_Valid_7_delay_11_1 <= io_A_Valid_7_delay_10_2;
    io_A_Valid_7_delay_12 <= io_A_Valid_7_delay_11_1;
    io_B_Valid_12_delay_1_6 <= io_B_Valid_12;
    io_B_Valid_12_delay_2_5 <= io_B_Valid_12_delay_1_6;
    io_B_Valid_12_delay_3_4 <= io_B_Valid_12_delay_2_5;
    io_B_Valid_12_delay_4_3 <= io_B_Valid_12_delay_3_4;
    io_B_Valid_12_delay_5_2 <= io_B_Valid_12_delay_4_3;
    io_B_Valid_12_delay_6_1 <= io_B_Valid_12_delay_5_2;
    io_B_Valid_12_delay_7 <= io_B_Valid_12_delay_6_1;
    io_A_Valid_7_delay_1_12 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_11 <= io_A_Valid_7_delay_1_12;
    io_A_Valid_7_delay_3_10 <= io_A_Valid_7_delay_2_11;
    io_A_Valid_7_delay_4_9 <= io_A_Valid_7_delay_3_10;
    io_A_Valid_7_delay_5_8 <= io_A_Valid_7_delay_4_9;
    io_A_Valid_7_delay_6_7 <= io_A_Valid_7_delay_5_8;
    io_A_Valid_7_delay_7_6 <= io_A_Valid_7_delay_6_7;
    io_A_Valid_7_delay_8_5 <= io_A_Valid_7_delay_7_6;
    io_A_Valid_7_delay_9_4 <= io_A_Valid_7_delay_8_5;
    io_A_Valid_7_delay_10_3 <= io_A_Valid_7_delay_9_4;
    io_A_Valid_7_delay_11_2 <= io_A_Valid_7_delay_10_3;
    io_A_Valid_7_delay_12_1 <= io_A_Valid_7_delay_11_2;
    io_A_Valid_7_delay_13 <= io_A_Valid_7_delay_12_1;
    io_B_Valid_13_delay_1_6 <= io_B_Valid_13;
    io_B_Valid_13_delay_2_5 <= io_B_Valid_13_delay_1_6;
    io_B_Valid_13_delay_3_4 <= io_B_Valid_13_delay_2_5;
    io_B_Valid_13_delay_4_3 <= io_B_Valid_13_delay_3_4;
    io_B_Valid_13_delay_5_2 <= io_B_Valid_13_delay_4_3;
    io_B_Valid_13_delay_6_1 <= io_B_Valid_13_delay_5_2;
    io_B_Valid_13_delay_7 <= io_B_Valid_13_delay_6_1;
    io_A_Valid_7_delay_1_13 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_12 <= io_A_Valid_7_delay_1_13;
    io_A_Valid_7_delay_3_11 <= io_A_Valid_7_delay_2_12;
    io_A_Valid_7_delay_4_10 <= io_A_Valid_7_delay_3_11;
    io_A_Valid_7_delay_5_9 <= io_A_Valid_7_delay_4_10;
    io_A_Valid_7_delay_6_8 <= io_A_Valid_7_delay_5_9;
    io_A_Valid_7_delay_7_7 <= io_A_Valid_7_delay_6_8;
    io_A_Valid_7_delay_8_6 <= io_A_Valid_7_delay_7_7;
    io_A_Valid_7_delay_9_5 <= io_A_Valid_7_delay_8_6;
    io_A_Valid_7_delay_10_4 <= io_A_Valid_7_delay_9_5;
    io_A_Valid_7_delay_11_3 <= io_A_Valid_7_delay_10_4;
    io_A_Valid_7_delay_12_2 <= io_A_Valid_7_delay_11_3;
    io_A_Valid_7_delay_13_1 <= io_A_Valid_7_delay_12_2;
    io_A_Valid_7_delay_14 <= io_A_Valid_7_delay_13_1;
    io_B_Valid_14_delay_1_6 <= io_B_Valid_14;
    io_B_Valid_14_delay_2_5 <= io_B_Valid_14_delay_1_6;
    io_B_Valid_14_delay_3_4 <= io_B_Valid_14_delay_2_5;
    io_B_Valid_14_delay_4_3 <= io_B_Valid_14_delay_3_4;
    io_B_Valid_14_delay_5_2 <= io_B_Valid_14_delay_4_3;
    io_B_Valid_14_delay_6_1 <= io_B_Valid_14_delay_5_2;
    io_B_Valid_14_delay_7 <= io_B_Valid_14_delay_6_1;
    io_A_Valid_7_delay_1_14 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_13 <= io_A_Valid_7_delay_1_14;
    io_A_Valid_7_delay_3_12 <= io_A_Valid_7_delay_2_13;
    io_A_Valid_7_delay_4_11 <= io_A_Valid_7_delay_3_12;
    io_A_Valid_7_delay_5_10 <= io_A_Valid_7_delay_4_11;
    io_A_Valid_7_delay_6_9 <= io_A_Valid_7_delay_5_10;
    io_A_Valid_7_delay_7_8 <= io_A_Valid_7_delay_6_9;
    io_A_Valid_7_delay_8_7 <= io_A_Valid_7_delay_7_8;
    io_A_Valid_7_delay_9_6 <= io_A_Valid_7_delay_8_7;
    io_A_Valid_7_delay_10_5 <= io_A_Valid_7_delay_9_6;
    io_A_Valid_7_delay_11_4 <= io_A_Valid_7_delay_10_5;
    io_A_Valid_7_delay_12_3 <= io_A_Valid_7_delay_11_4;
    io_A_Valid_7_delay_13_2 <= io_A_Valid_7_delay_12_3;
    io_A_Valid_7_delay_14_1 <= io_A_Valid_7_delay_13_2;
    io_A_Valid_7_delay_15 <= io_A_Valid_7_delay_14_1;
    io_B_Valid_15_delay_1_6 <= io_B_Valid_15;
    io_B_Valid_15_delay_2_5 <= io_B_Valid_15_delay_1_6;
    io_B_Valid_15_delay_3_4 <= io_B_Valid_15_delay_2_5;
    io_B_Valid_15_delay_4_3 <= io_B_Valid_15_delay_3_4;
    io_B_Valid_15_delay_5_2 <= io_B_Valid_15_delay_4_3;
    io_B_Valid_15_delay_6_1 <= io_B_Valid_15_delay_5_2;
    io_B_Valid_15_delay_7 <= io_B_Valid_15_delay_6_1;
    io_A_Valid_7_delay_1_15 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_14 <= io_A_Valid_7_delay_1_15;
    io_A_Valid_7_delay_3_13 <= io_A_Valid_7_delay_2_14;
    io_A_Valid_7_delay_4_12 <= io_A_Valid_7_delay_3_13;
    io_A_Valid_7_delay_5_11 <= io_A_Valid_7_delay_4_12;
    io_A_Valid_7_delay_6_10 <= io_A_Valid_7_delay_5_11;
    io_A_Valid_7_delay_7_9 <= io_A_Valid_7_delay_6_10;
    io_A_Valid_7_delay_8_8 <= io_A_Valid_7_delay_7_9;
    io_A_Valid_7_delay_9_7 <= io_A_Valid_7_delay_8_8;
    io_A_Valid_7_delay_10_6 <= io_A_Valid_7_delay_9_7;
    io_A_Valid_7_delay_11_5 <= io_A_Valid_7_delay_10_6;
    io_A_Valid_7_delay_12_4 <= io_A_Valid_7_delay_11_5;
    io_A_Valid_7_delay_13_3 <= io_A_Valid_7_delay_12_4;
    io_A_Valid_7_delay_14_2 <= io_A_Valid_7_delay_13_3;
    io_A_Valid_7_delay_15_1 <= io_A_Valid_7_delay_14_2;
    io_A_Valid_7_delay_16 <= io_A_Valid_7_delay_15_1;
    io_B_Valid_16_delay_1_6 <= io_B_Valid_16;
    io_B_Valid_16_delay_2_5 <= io_B_Valid_16_delay_1_6;
    io_B_Valid_16_delay_3_4 <= io_B_Valid_16_delay_2_5;
    io_B_Valid_16_delay_4_3 <= io_B_Valid_16_delay_3_4;
    io_B_Valid_16_delay_5_2 <= io_B_Valid_16_delay_4_3;
    io_B_Valid_16_delay_6_1 <= io_B_Valid_16_delay_5_2;
    io_B_Valid_16_delay_7 <= io_B_Valid_16_delay_6_1;
    io_A_Valid_7_delay_1_16 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_15 <= io_A_Valid_7_delay_1_16;
    io_A_Valid_7_delay_3_14 <= io_A_Valid_7_delay_2_15;
    io_A_Valid_7_delay_4_13 <= io_A_Valid_7_delay_3_14;
    io_A_Valid_7_delay_5_12 <= io_A_Valid_7_delay_4_13;
    io_A_Valid_7_delay_6_11 <= io_A_Valid_7_delay_5_12;
    io_A_Valid_7_delay_7_10 <= io_A_Valid_7_delay_6_11;
    io_A_Valid_7_delay_8_9 <= io_A_Valid_7_delay_7_10;
    io_A_Valid_7_delay_9_8 <= io_A_Valid_7_delay_8_9;
    io_A_Valid_7_delay_10_7 <= io_A_Valid_7_delay_9_8;
    io_A_Valid_7_delay_11_6 <= io_A_Valid_7_delay_10_7;
    io_A_Valid_7_delay_12_5 <= io_A_Valid_7_delay_11_6;
    io_A_Valid_7_delay_13_4 <= io_A_Valid_7_delay_12_5;
    io_A_Valid_7_delay_14_3 <= io_A_Valid_7_delay_13_4;
    io_A_Valid_7_delay_15_2 <= io_A_Valid_7_delay_14_3;
    io_A_Valid_7_delay_16_1 <= io_A_Valid_7_delay_15_2;
    io_A_Valid_7_delay_17 <= io_A_Valid_7_delay_16_1;
    io_B_Valid_17_delay_1_6 <= io_B_Valid_17;
    io_B_Valid_17_delay_2_5 <= io_B_Valid_17_delay_1_6;
    io_B_Valid_17_delay_3_4 <= io_B_Valid_17_delay_2_5;
    io_B_Valid_17_delay_4_3 <= io_B_Valid_17_delay_3_4;
    io_B_Valid_17_delay_5_2 <= io_B_Valid_17_delay_4_3;
    io_B_Valid_17_delay_6_1 <= io_B_Valid_17_delay_5_2;
    io_B_Valid_17_delay_7 <= io_B_Valid_17_delay_6_1;
    io_A_Valid_7_delay_1_17 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_16 <= io_A_Valid_7_delay_1_17;
    io_A_Valid_7_delay_3_15 <= io_A_Valid_7_delay_2_16;
    io_A_Valid_7_delay_4_14 <= io_A_Valid_7_delay_3_15;
    io_A_Valid_7_delay_5_13 <= io_A_Valid_7_delay_4_14;
    io_A_Valid_7_delay_6_12 <= io_A_Valid_7_delay_5_13;
    io_A_Valid_7_delay_7_11 <= io_A_Valid_7_delay_6_12;
    io_A_Valid_7_delay_8_10 <= io_A_Valid_7_delay_7_11;
    io_A_Valid_7_delay_9_9 <= io_A_Valid_7_delay_8_10;
    io_A_Valid_7_delay_10_8 <= io_A_Valid_7_delay_9_9;
    io_A_Valid_7_delay_11_7 <= io_A_Valid_7_delay_10_8;
    io_A_Valid_7_delay_12_6 <= io_A_Valid_7_delay_11_7;
    io_A_Valid_7_delay_13_5 <= io_A_Valid_7_delay_12_6;
    io_A_Valid_7_delay_14_4 <= io_A_Valid_7_delay_13_5;
    io_A_Valid_7_delay_15_3 <= io_A_Valid_7_delay_14_4;
    io_A_Valid_7_delay_16_2 <= io_A_Valid_7_delay_15_3;
    io_A_Valid_7_delay_17_1 <= io_A_Valid_7_delay_16_2;
    io_A_Valid_7_delay_18 <= io_A_Valid_7_delay_17_1;
    io_B_Valid_18_delay_1_6 <= io_B_Valid_18;
    io_B_Valid_18_delay_2_5 <= io_B_Valid_18_delay_1_6;
    io_B_Valid_18_delay_3_4 <= io_B_Valid_18_delay_2_5;
    io_B_Valid_18_delay_4_3 <= io_B_Valid_18_delay_3_4;
    io_B_Valid_18_delay_5_2 <= io_B_Valid_18_delay_4_3;
    io_B_Valid_18_delay_6_1 <= io_B_Valid_18_delay_5_2;
    io_B_Valid_18_delay_7 <= io_B_Valid_18_delay_6_1;
    io_A_Valid_7_delay_1_18 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_17 <= io_A_Valid_7_delay_1_18;
    io_A_Valid_7_delay_3_16 <= io_A_Valid_7_delay_2_17;
    io_A_Valid_7_delay_4_15 <= io_A_Valid_7_delay_3_16;
    io_A_Valid_7_delay_5_14 <= io_A_Valid_7_delay_4_15;
    io_A_Valid_7_delay_6_13 <= io_A_Valid_7_delay_5_14;
    io_A_Valid_7_delay_7_12 <= io_A_Valid_7_delay_6_13;
    io_A_Valid_7_delay_8_11 <= io_A_Valid_7_delay_7_12;
    io_A_Valid_7_delay_9_10 <= io_A_Valid_7_delay_8_11;
    io_A_Valid_7_delay_10_9 <= io_A_Valid_7_delay_9_10;
    io_A_Valid_7_delay_11_8 <= io_A_Valid_7_delay_10_9;
    io_A_Valid_7_delay_12_7 <= io_A_Valid_7_delay_11_8;
    io_A_Valid_7_delay_13_6 <= io_A_Valid_7_delay_12_7;
    io_A_Valid_7_delay_14_5 <= io_A_Valid_7_delay_13_6;
    io_A_Valid_7_delay_15_4 <= io_A_Valid_7_delay_14_5;
    io_A_Valid_7_delay_16_3 <= io_A_Valid_7_delay_15_4;
    io_A_Valid_7_delay_17_2 <= io_A_Valid_7_delay_16_3;
    io_A_Valid_7_delay_18_1 <= io_A_Valid_7_delay_17_2;
    io_A_Valid_7_delay_19 <= io_A_Valid_7_delay_18_1;
    io_B_Valid_19_delay_1_6 <= io_B_Valid_19;
    io_B_Valid_19_delay_2_5 <= io_B_Valid_19_delay_1_6;
    io_B_Valid_19_delay_3_4 <= io_B_Valid_19_delay_2_5;
    io_B_Valid_19_delay_4_3 <= io_B_Valid_19_delay_3_4;
    io_B_Valid_19_delay_5_2 <= io_B_Valid_19_delay_4_3;
    io_B_Valid_19_delay_6_1 <= io_B_Valid_19_delay_5_2;
    io_B_Valid_19_delay_7 <= io_B_Valid_19_delay_6_1;
    io_A_Valid_7_delay_1_19 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_18 <= io_A_Valid_7_delay_1_19;
    io_A_Valid_7_delay_3_17 <= io_A_Valid_7_delay_2_18;
    io_A_Valid_7_delay_4_16 <= io_A_Valid_7_delay_3_17;
    io_A_Valid_7_delay_5_15 <= io_A_Valid_7_delay_4_16;
    io_A_Valid_7_delay_6_14 <= io_A_Valid_7_delay_5_15;
    io_A_Valid_7_delay_7_13 <= io_A_Valid_7_delay_6_14;
    io_A_Valid_7_delay_8_12 <= io_A_Valid_7_delay_7_13;
    io_A_Valid_7_delay_9_11 <= io_A_Valid_7_delay_8_12;
    io_A_Valid_7_delay_10_10 <= io_A_Valid_7_delay_9_11;
    io_A_Valid_7_delay_11_9 <= io_A_Valid_7_delay_10_10;
    io_A_Valid_7_delay_12_8 <= io_A_Valid_7_delay_11_9;
    io_A_Valid_7_delay_13_7 <= io_A_Valid_7_delay_12_8;
    io_A_Valid_7_delay_14_6 <= io_A_Valid_7_delay_13_7;
    io_A_Valid_7_delay_15_5 <= io_A_Valid_7_delay_14_6;
    io_A_Valid_7_delay_16_4 <= io_A_Valid_7_delay_15_5;
    io_A_Valid_7_delay_17_3 <= io_A_Valid_7_delay_16_4;
    io_A_Valid_7_delay_18_2 <= io_A_Valid_7_delay_17_3;
    io_A_Valid_7_delay_19_1 <= io_A_Valid_7_delay_18_2;
    io_A_Valid_7_delay_20 <= io_A_Valid_7_delay_19_1;
    io_B_Valid_20_delay_1_6 <= io_B_Valid_20;
    io_B_Valid_20_delay_2_5 <= io_B_Valid_20_delay_1_6;
    io_B_Valid_20_delay_3_4 <= io_B_Valid_20_delay_2_5;
    io_B_Valid_20_delay_4_3 <= io_B_Valid_20_delay_3_4;
    io_B_Valid_20_delay_5_2 <= io_B_Valid_20_delay_4_3;
    io_B_Valid_20_delay_6_1 <= io_B_Valid_20_delay_5_2;
    io_B_Valid_20_delay_7 <= io_B_Valid_20_delay_6_1;
    io_A_Valid_7_delay_1_20 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_19 <= io_A_Valid_7_delay_1_20;
    io_A_Valid_7_delay_3_18 <= io_A_Valid_7_delay_2_19;
    io_A_Valid_7_delay_4_17 <= io_A_Valid_7_delay_3_18;
    io_A_Valid_7_delay_5_16 <= io_A_Valid_7_delay_4_17;
    io_A_Valid_7_delay_6_15 <= io_A_Valid_7_delay_5_16;
    io_A_Valid_7_delay_7_14 <= io_A_Valid_7_delay_6_15;
    io_A_Valid_7_delay_8_13 <= io_A_Valid_7_delay_7_14;
    io_A_Valid_7_delay_9_12 <= io_A_Valid_7_delay_8_13;
    io_A_Valid_7_delay_10_11 <= io_A_Valid_7_delay_9_12;
    io_A_Valid_7_delay_11_10 <= io_A_Valid_7_delay_10_11;
    io_A_Valid_7_delay_12_9 <= io_A_Valid_7_delay_11_10;
    io_A_Valid_7_delay_13_8 <= io_A_Valid_7_delay_12_9;
    io_A_Valid_7_delay_14_7 <= io_A_Valid_7_delay_13_8;
    io_A_Valid_7_delay_15_6 <= io_A_Valid_7_delay_14_7;
    io_A_Valid_7_delay_16_5 <= io_A_Valid_7_delay_15_6;
    io_A_Valid_7_delay_17_4 <= io_A_Valid_7_delay_16_5;
    io_A_Valid_7_delay_18_3 <= io_A_Valid_7_delay_17_4;
    io_A_Valid_7_delay_19_2 <= io_A_Valid_7_delay_18_3;
    io_A_Valid_7_delay_20_1 <= io_A_Valid_7_delay_19_2;
    io_A_Valid_7_delay_21 <= io_A_Valid_7_delay_20_1;
    io_B_Valid_21_delay_1_6 <= io_B_Valid_21;
    io_B_Valid_21_delay_2_5 <= io_B_Valid_21_delay_1_6;
    io_B_Valid_21_delay_3_4 <= io_B_Valid_21_delay_2_5;
    io_B_Valid_21_delay_4_3 <= io_B_Valid_21_delay_3_4;
    io_B_Valid_21_delay_5_2 <= io_B_Valid_21_delay_4_3;
    io_B_Valid_21_delay_6_1 <= io_B_Valid_21_delay_5_2;
    io_B_Valid_21_delay_7 <= io_B_Valid_21_delay_6_1;
    io_A_Valid_7_delay_1_21 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_20 <= io_A_Valid_7_delay_1_21;
    io_A_Valid_7_delay_3_19 <= io_A_Valid_7_delay_2_20;
    io_A_Valid_7_delay_4_18 <= io_A_Valid_7_delay_3_19;
    io_A_Valid_7_delay_5_17 <= io_A_Valid_7_delay_4_18;
    io_A_Valid_7_delay_6_16 <= io_A_Valid_7_delay_5_17;
    io_A_Valid_7_delay_7_15 <= io_A_Valid_7_delay_6_16;
    io_A_Valid_7_delay_8_14 <= io_A_Valid_7_delay_7_15;
    io_A_Valid_7_delay_9_13 <= io_A_Valid_7_delay_8_14;
    io_A_Valid_7_delay_10_12 <= io_A_Valid_7_delay_9_13;
    io_A_Valid_7_delay_11_11 <= io_A_Valid_7_delay_10_12;
    io_A_Valid_7_delay_12_10 <= io_A_Valid_7_delay_11_11;
    io_A_Valid_7_delay_13_9 <= io_A_Valid_7_delay_12_10;
    io_A_Valid_7_delay_14_8 <= io_A_Valid_7_delay_13_9;
    io_A_Valid_7_delay_15_7 <= io_A_Valid_7_delay_14_8;
    io_A_Valid_7_delay_16_6 <= io_A_Valid_7_delay_15_7;
    io_A_Valid_7_delay_17_5 <= io_A_Valid_7_delay_16_6;
    io_A_Valid_7_delay_18_4 <= io_A_Valid_7_delay_17_5;
    io_A_Valid_7_delay_19_3 <= io_A_Valid_7_delay_18_4;
    io_A_Valid_7_delay_20_2 <= io_A_Valid_7_delay_19_3;
    io_A_Valid_7_delay_21_1 <= io_A_Valid_7_delay_20_2;
    io_A_Valid_7_delay_22 <= io_A_Valid_7_delay_21_1;
    io_B_Valid_22_delay_1_6 <= io_B_Valid_22;
    io_B_Valid_22_delay_2_5 <= io_B_Valid_22_delay_1_6;
    io_B_Valid_22_delay_3_4 <= io_B_Valid_22_delay_2_5;
    io_B_Valid_22_delay_4_3 <= io_B_Valid_22_delay_3_4;
    io_B_Valid_22_delay_5_2 <= io_B_Valid_22_delay_4_3;
    io_B_Valid_22_delay_6_1 <= io_B_Valid_22_delay_5_2;
    io_B_Valid_22_delay_7 <= io_B_Valid_22_delay_6_1;
    io_A_Valid_7_delay_1_22 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_21 <= io_A_Valid_7_delay_1_22;
    io_A_Valid_7_delay_3_20 <= io_A_Valid_7_delay_2_21;
    io_A_Valid_7_delay_4_19 <= io_A_Valid_7_delay_3_20;
    io_A_Valid_7_delay_5_18 <= io_A_Valid_7_delay_4_19;
    io_A_Valid_7_delay_6_17 <= io_A_Valid_7_delay_5_18;
    io_A_Valid_7_delay_7_16 <= io_A_Valid_7_delay_6_17;
    io_A_Valid_7_delay_8_15 <= io_A_Valid_7_delay_7_16;
    io_A_Valid_7_delay_9_14 <= io_A_Valid_7_delay_8_15;
    io_A_Valid_7_delay_10_13 <= io_A_Valid_7_delay_9_14;
    io_A_Valid_7_delay_11_12 <= io_A_Valid_7_delay_10_13;
    io_A_Valid_7_delay_12_11 <= io_A_Valid_7_delay_11_12;
    io_A_Valid_7_delay_13_10 <= io_A_Valid_7_delay_12_11;
    io_A_Valid_7_delay_14_9 <= io_A_Valid_7_delay_13_10;
    io_A_Valid_7_delay_15_8 <= io_A_Valid_7_delay_14_9;
    io_A_Valid_7_delay_16_7 <= io_A_Valid_7_delay_15_8;
    io_A_Valid_7_delay_17_6 <= io_A_Valid_7_delay_16_7;
    io_A_Valid_7_delay_18_5 <= io_A_Valid_7_delay_17_6;
    io_A_Valid_7_delay_19_4 <= io_A_Valid_7_delay_18_5;
    io_A_Valid_7_delay_20_3 <= io_A_Valid_7_delay_19_4;
    io_A_Valid_7_delay_21_2 <= io_A_Valid_7_delay_20_3;
    io_A_Valid_7_delay_22_1 <= io_A_Valid_7_delay_21_2;
    io_A_Valid_7_delay_23 <= io_A_Valid_7_delay_22_1;
    io_B_Valid_23_delay_1_6 <= io_B_Valid_23;
    io_B_Valid_23_delay_2_5 <= io_B_Valid_23_delay_1_6;
    io_B_Valid_23_delay_3_4 <= io_B_Valid_23_delay_2_5;
    io_B_Valid_23_delay_4_3 <= io_B_Valid_23_delay_3_4;
    io_B_Valid_23_delay_5_2 <= io_B_Valid_23_delay_4_3;
    io_B_Valid_23_delay_6_1 <= io_B_Valid_23_delay_5_2;
    io_B_Valid_23_delay_7 <= io_B_Valid_23_delay_6_1;
    io_A_Valid_7_delay_1_23 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_22 <= io_A_Valid_7_delay_1_23;
    io_A_Valid_7_delay_3_21 <= io_A_Valid_7_delay_2_22;
    io_A_Valid_7_delay_4_20 <= io_A_Valid_7_delay_3_21;
    io_A_Valid_7_delay_5_19 <= io_A_Valid_7_delay_4_20;
    io_A_Valid_7_delay_6_18 <= io_A_Valid_7_delay_5_19;
    io_A_Valid_7_delay_7_17 <= io_A_Valid_7_delay_6_18;
    io_A_Valid_7_delay_8_16 <= io_A_Valid_7_delay_7_17;
    io_A_Valid_7_delay_9_15 <= io_A_Valid_7_delay_8_16;
    io_A_Valid_7_delay_10_14 <= io_A_Valid_7_delay_9_15;
    io_A_Valid_7_delay_11_13 <= io_A_Valid_7_delay_10_14;
    io_A_Valid_7_delay_12_12 <= io_A_Valid_7_delay_11_13;
    io_A_Valid_7_delay_13_11 <= io_A_Valid_7_delay_12_12;
    io_A_Valid_7_delay_14_10 <= io_A_Valid_7_delay_13_11;
    io_A_Valid_7_delay_15_9 <= io_A_Valid_7_delay_14_10;
    io_A_Valid_7_delay_16_8 <= io_A_Valid_7_delay_15_9;
    io_A_Valid_7_delay_17_7 <= io_A_Valid_7_delay_16_8;
    io_A_Valid_7_delay_18_6 <= io_A_Valid_7_delay_17_7;
    io_A_Valid_7_delay_19_5 <= io_A_Valid_7_delay_18_6;
    io_A_Valid_7_delay_20_4 <= io_A_Valid_7_delay_19_5;
    io_A_Valid_7_delay_21_3 <= io_A_Valid_7_delay_20_4;
    io_A_Valid_7_delay_22_2 <= io_A_Valid_7_delay_21_3;
    io_A_Valid_7_delay_23_1 <= io_A_Valid_7_delay_22_2;
    io_A_Valid_7_delay_24 <= io_A_Valid_7_delay_23_1;
    io_B_Valid_24_delay_1_6 <= io_B_Valid_24;
    io_B_Valid_24_delay_2_5 <= io_B_Valid_24_delay_1_6;
    io_B_Valid_24_delay_3_4 <= io_B_Valid_24_delay_2_5;
    io_B_Valid_24_delay_4_3 <= io_B_Valid_24_delay_3_4;
    io_B_Valid_24_delay_5_2 <= io_B_Valid_24_delay_4_3;
    io_B_Valid_24_delay_6_1 <= io_B_Valid_24_delay_5_2;
    io_B_Valid_24_delay_7 <= io_B_Valid_24_delay_6_1;
    io_A_Valid_7_delay_1_24 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_23 <= io_A_Valid_7_delay_1_24;
    io_A_Valid_7_delay_3_22 <= io_A_Valid_7_delay_2_23;
    io_A_Valid_7_delay_4_21 <= io_A_Valid_7_delay_3_22;
    io_A_Valid_7_delay_5_20 <= io_A_Valid_7_delay_4_21;
    io_A_Valid_7_delay_6_19 <= io_A_Valid_7_delay_5_20;
    io_A_Valid_7_delay_7_18 <= io_A_Valid_7_delay_6_19;
    io_A_Valid_7_delay_8_17 <= io_A_Valid_7_delay_7_18;
    io_A_Valid_7_delay_9_16 <= io_A_Valid_7_delay_8_17;
    io_A_Valid_7_delay_10_15 <= io_A_Valid_7_delay_9_16;
    io_A_Valid_7_delay_11_14 <= io_A_Valid_7_delay_10_15;
    io_A_Valid_7_delay_12_13 <= io_A_Valid_7_delay_11_14;
    io_A_Valid_7_delay_13_12 <= io_A_Valid_7_delay_12_13;
    io_A_Valid_7_delay_14_11 <= io_A_Valid_7_delay_13_12;
    io_A_Valid_7_delay_15_10 <= io_A_Valid_7_delay_14_11;
    io_A_Valid_7_delay_16_9 <= io_A_Valid_7_delay_15_10;
    io_A_Valid_7_delay_17_8 <= io_A_Valid_7_delay_16_9;
    io_A_Valid_7_delay_18_7 <= io_A_Valid_7_delay_17_8;
    io_A_Valid_7_delay_19_6 <= io_A_Valid_7_delay_18_7;
    io_A_Valid_7_delay_20_5 <= io_A_Valid_7_delay_19_6;
    io_A_Valid_7_delay_21_4 <= io_A_Valid_7_delay_20_5;
    io_A_Valid_7_delay_22_3 <= io_A_Valid_7_delay_21_4;
    io_A_Valid_7_delay_23_2 <= io_A_Valid_7_delay_22_3;
    io_A_Valid_7_delay_24_1 <= io_A_Valid_7_delay_23_2;
    io_A_Valid_7_delay_25 <= io_A_Valid_7_delay_24_1;
    io_B_Valid_25_delay_1_6 <= io_B_Valid_25;
    io_B_Valid_25_delay_2_5 <= io_B_Valid_25_delay_1_6;
    io_B_Valid_25_delay_3_4 <= io_B_Valid_25_delay_2_5;
    io_B_Valid_25_delay_4_3 <= io_B_Valid_25_delay_3_4;
    io_B_Valid_25_delay_5_2 <= io_B_Valid_25_delay_4_3;
    io_B_Valid_25_delay_6_1 <= io_B_Valid_25_delay_5_2;
    io_B_Valid_25_delay_7 <= io_B_Valid_25_delay_6_1;
    io_A_Valid_7_delay_1_25 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_24 <= io_A_Valid_7_delay_1_25;
    io_A_Valid_7_delay_3_23 <= io_A_Valid_7_delay_2_24;
    io_A_Valid_7_delay_4_22 <= io_A_Valid_7_delay_3_23;
    io_A_Valid_7_delay_5_21 <= io_A_Valid_7_delay_4_22;
    io_A_Valid_7_delay_6_20 <= io_A_Valid_7_delay_5_21;
    io_A_Valid_7_delay_7_19 <= io_A_Valid_7_delay_6_20;
    io_A_Valid_7_delay_8_18 <= io_A_Valid_7_delay_7_19;
    io_A_Valid_7_delay_9_17 <= io_A_Valid_7_delay_8_18;
    io_A_Valid_7_delay_10_16 <= io_A_Valid_7_delay_9_17;
    io_A_Valid_7_delay_11_15 <= io_A_Valid_7_delay_10_16;
    io_A_Valid_7_delay_12_14 <= io_A_Valid_7_delay_11_15;
    io_A_Valid_7_delay_13_13 <= io_A_Valid_7_delay_12_14;
    io_A_Valid_7_delay_14_12 <= io_A_Valid_7_delay_13_13;
    io_A_Valid_7_delay_15_11 <= io_A_Valid_7_delay_14_12;
    io_A_Valid_7_delay_16_10 <= io_A_Valid_7_delay_15_11;
    io_A_Valid_7_delay_17_9 <= io_A_Valid_7_delay_16_10;
    io_A_Valid_7_delay_18_8 <= io_A_Valid_7_delay_17_9;
    io_A_Valid_7_delay_19_7 <= io_A_Valid_7_delay_18_8;
    io_A_Valid_7_delay_20_6 <= io_A_Valid_7_delay_19_7;
    io_A_Valid_7_delay_21_5 <= io_A_Valid_7_delay_20_6;
    io_A_Valid_7_delay_22_4 <= io_A_Valid_7_delay_21_5;
    io_A_Valid_7_delay_23_3 <= io_A_Valid_7_delay_22_4;
    io_A_Valid_7_delay_24_2 <= io_A_Valid_7_delay_23_3;
    io_A_Valid_7_delay_25_1 <= io_A_Valid_7_delay_24_2;
    io_A_Valid_7_delay_26 <= io_A_Valid_7_delay_25_1;
    io_B_Valid_26_delay_1_6 <= io_B_Valid_26;
    io_B_Valid_26_delay_2_5 <= io_B_Valid_26_delay_1_6;
    io_B_Valid_26_delay_3_4 <= io_B_Valid_26_delay_2_5;
    io_B_Valid_26_delay_4_3 <= io_B_Valid_26_delay_3_4;
    io_B_Valid_26_delay_5_2 <= io_B_Valid_26_delay_4_3;
    io_B_Valid_26_delay_6_1 <= io_B_Valid_26_delay_5_2;
    io_B_Valid_26_delay_7 <= io_B_Valid_26_delay_6_1;
    io_A_Valid_7_delay_1_26 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_25 <= io_A_Valid_7_delay_1_26;
    io_A_Valid_7_delay_3_24 <= io_A_Valid_7_delay_2_25;
    io_A_Valid_7_delay_4_23 <= io_A_Valid_7_delay_3_24;
    io_A_Valid_7_delay_5_22 <= io_A_Valid_7_delay_4_23;
    io_A_Valid_7_delay_6_21 <= io_A_Valid_7_delay_5_22;
    io_A_Valid_7_delay_7_20 <= io_A_Valid_7_delay_6_21;
    io_A_Valid_7_delay_8_19 <= io_A_Valid_7_delay_7_20;
    io_A_Valid_7_delay_9_18 <= io_A_Valid_7_delay_8_19;
    io_A_Valid_7_delay_10_17 <= io_A_Valid_7_delay_9_18;
    io_A_Valid_7_delay_11_16 <= io_A_Valid_7_delay_10_17;
    io_A_Valid_7_delay_12_15 <= io_A_Valid_7_delay_11_16;
    io_A_Valid_7_delay_13_14 <= io_A_Valid_7_delay_12_15;
    io_A_Valid_7_delay_14_13 <= io_A_Valid_7_delay_13_14;
    io_A_Valid_7_delay_15_12 <= io_A_Valid_7_delay_14_13;
    io_A_Valid_7_delay_16_11 <= io_A_Valid_7_delay_15_12;
    io_A_Valid_7_delay_17_10 <= io_A_Valid_7_delay_16_11;
    io_A_Valid_7_delay_18_9 <= io_A_Valid_7_delay_17_10;
    io_A_Valid_7_delay_19_8 <= io_A_Valid_7_delay_18_9;
    io_A_Valid_7_delay_20_7 <= io_A_Valid_7_delay_19_8;
    io_A_Valid_7_delay_21_6 <= io_A_Valid_7_delay_20_7;
    io_A_Valid_7_delay_22_5 <= io_A_Valid_7_delay_21_6;
    io_A_Valid_7_delay_23_4 <= io_A_Valid_7_delay_22_5;
    io_A_Valid_7_delay_24_3 <= io_A_Valid_7_delay_23_4;
    io_A_Valid_7_delay_25_2 <= io_A_Valid_7_delay_24_3;
    io_A_Valid_7_delay_26_1 <= io_A_Valid_7_delay_25_2;
    io_A_Valid_7_delay_27 <= io_A_Valid_7_delay_26_1;
    io_B_Valid_27_delay_1_6 <= io_B_Valid_27;
    io_B_Valid_27_delay_2_5 <= io_B_Valid_27_delay_1_6;
    io_B_Valid_27_delay_3_4 <= io_B_Valid_27_delay_2_5;
    io_B_Valid_27_delay_4_3 <= io_B_Valid_27_delay_3_4;
    io_B_Valid_27_delay_5_2 <= io_B_Valid_27_delay_4_3;
    io_B_Valid_27_delay_6_1 <= io_B_Valid_27_delay_5_2;
    io_B_Valid_27_delay_7 <= io_B_Valid_27_delay_6_1;
    io_A_Valid_7_delay_1_27 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_26 <= io_A_Valid_7_delay_1_27;
    io_A_Valid_7_delay_3_25 <= io_A_Valid_7_delay_2_26;
    io_A_Valid_7_delay_4_24 <= io_A_Valid_7_delay_3_25;
    io_A_Valid_7_delay_5_23 <= io_A_Valid_7_delay_4_24;
    io_A_Valid_7_delay_6_22 <= io_A_Valid_7_delay_5_23;
    io_A_Valid_7_delay_7_21 <= io_A_Valid_7_delay_6_22;
    io_A_Valid_7_delay_8_20 <= io_A_Valid_7_delay_7_21;
    io_A_Valid_7_delay_9_19 <= io_A_Valid_7_delay_8_20;
    io_A_Valid_7_delay_10_18 <= io_A_Valid_7_delay_9_19;
    io_A_Valid_7_delay_11_17 <= io_A_Valid_7_delay_10_18;
    io_A_Valid_7_delay_12_16 <= io_A_Valid_7_delay_11_17;
    io_A_Valid_7_delay_13_15 <= io_A_Valid_7_delay_12_16;
    io_A_Valid_7_delay_14_14 <= io_A_Valid_7_delay_13_15;
    io_A_Valid_7_delay_15_13 <= io_A_Valid_7_delay_14_14;
    io_A_Valid_7_delay_16_12 <= io_A_Valid_7_delay_15_13;
    io_A_Valid_7_delay_17_11 <= io_A_Valid_7_delay_16_12;
    io_A_Valid_7_delay_18_10 <= io_A_Valid_7_delay_17_11;
    io_A_Valid_7_delay_19_9 <= io_A_Valid_7_delay_18_10;
    io_A_Valid_7_delay_20_8 <= io_A_Valid_7_delay_19_9;
    io_A_Valid_7_delay_21_7 <= io_A_Valid_7_delay_20_8;
    io_A_Valid_7_delay_22_6 <= io_A_Valid_7_delay_21_7;
    io_A_Valid_7_delay_23_5 <= io_A_Valid_7_delay_22_6;
    io_A_Valid_7_delay_24_4 <= io_A_Valid_7_delay_23_5;
    io_A_Valid_7_delay_25_3 <= io_A_Valid_7_delay_24_4;
    io_A_Valid_7_delay_26_2 <= io_A_Valid_7_delay_25_3;
    io_A_Valid_7_delay_27_1 <= io_A_Valid_7_delay_26_2;
    io_A_Valid_7_delay_28 <= io_A_Valid_7_delay_27_1;
    io_B_Valid_28_delay_1_6 <= io_B_Valid_28;
    io_B_Valid_28_delay_2_5 <= io_B_Valid_28_delay_1_6;
    io_B_Valid_28_delay_3_4 <= io_B_Valid_28_delay_2_5;
    io_B_Valid_28_delay_4_3 <= io_B_Valid_28_delay_3_4;
    io_B_Valid_28_delay_5_2 <= io_B_Valid_28_delay_4_3;
    io_B_Valid_28_delay_6_1 <= io_B_Valid_28_delay_5_2;
    io_B_Valid_28_delay_7 <= io_B_Valid_28_delay_6_1;
    io_A_Valid_7_delay_1_28 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_27 <= io_A_Valid_7_delay_1_28;
    io_A_Valid_7_delay_3_26 <= io_A_Valid_7_delay_2_27;
    io_A_Valid_7_delay_4_25 <= io_A_Valid_7_delay_3_26;
    io_A_Valid_7_delay_5_24 <= io_A_Valid_7_delay_4_25;
    io_A_Valid_7_delay_6_23 <= io_A_Valid_7_delay_5_24;
    io_A_Valid_7_delay_7_22 <= io_A_Valid_7_delay_6_23;
    io_A_Valid_7_delay_8_21 <= io_A_Valid_7_delay_7_22;
    io_A_Valid_7_delay_9_20 <= io_A_Valid_7_delay_8_21;
    io_A_Valid_7_delay_10_19 <= io_A_Valid_7_delay_9_20;
    io_A_Valid_7_delay_11_18 <= io_A_Valid_7_delay_10_19;
    io_A_Valid_7_delay_12_17 <= io_A_Valid_7_delay_11_18;
    io_A_Valid_7_delay_13_16 <= io_A_Valid_7_delay_12_17;
    io_A_Valid_7_delay_14_15 <= io_A_Valid_7_delay_13_16;
    io_A_Valid_7_delay_15_14 <= io_A_Valid_7_delay_14_15;
    io_A_Valid_7_delay_16_13 <= io_A_Valid_7_delay_15_14;
    io_A_Valid_7_delay_17_12 <= io_A_Valid_7_delay_16_13;
    io_A_Valid_7_delay_18_11 <= io_A_Valid_7_delay_17_12;
    io_A_Valid_7_delay_19_10 <= io_A_Valid_7_delay_18_11;
    io_A_Valid_7_delay_20_9 <= io_A_Valid_7_delay_19_10;
    io_A_Valid_7_delay_21_8 <= io_A_Valid_7_delay_20_9;
    io_A_Valid_7_delay_22_7 <= io_A_Valid_7_delay_21_8;
    io_A_Valid_7_delay_23_6 <= io_A_Valid_7_delay_22_7;
    io_A_Valid_7_delay_24_5 <= io_A_Valid_7_delay_23_6;
    io_A_Valid_7_delay_25_4 <= io_A_Valid_7_delay_24_5;
    io_A_Valid_7_delay_26_3 <= io_A_Valid_7_delay_25_4;
    io_A_Valid_7_delay_27_2 <= io_A_Valid_7_delay_26_3;
    io_A_Valid_7_delay_28_1 <= io_A_Valid_7_delay_27_2;
    io_A_Valid_7_delay_29 <= io_A_Valid_7_delay_28_1;
    io_B_Valid_29_delay_1_6 <= io_B_Valid_29;
    io_B_Valid_29_delay_2_5 <= io_B_Valid_29_delay_1_6;
    io_B_Valid_29_delay_3_4 <= io_B_Valid_29_delay_2_5;
    io_B_Valid_29_delay_4_3 <= io_B_Valid_29_delay_3_4;
    io_B_Valid_29_delay_5_2 <= io_B_Valid_29_delay_4_3;
    io_B_Valid_29_delay_6_1 <= io_B_Valid_29_delay_5_2;
    io_B_Valid_29_delay_7 <= io_B_Valid_29_delay_6_1;
    io_A_Valid_7_delay_1_29 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_28 <= io_A_Valid_7_delay_1_29;
    io_A_Valid_7_delay_3_27 <= io_A_Valid_7_delay_2_28;
    io_A_Valid_7_delay_4_26 <= io_A_Valid_7_delay_3_27;
    io_A_Valid_7_delay_5_25 <= io_A_Valid_7_delay_4_26;
    io_A_Valid_7_delay_6_24 <= io_A_Valid_7_delay_5_25;
    io_A_Valid_7_delay_7_23 <= io_A_Valid_7_delay_6_24;
    io_A_Valid_7_delay_8_22 <= io_A_Valid_7_delay_7_23;
    io_A_Valid_7_delay_9_21 <= io_A_Valid_7_delay_8_22;
    io_A_Valid_7_delay_10_20 <= io_A_Valid_7_delay_9_21;
    io_A_Valid_7_delay_11_19 <= io_A_Valid_7_delay_10_20;
    io_A_Valid_7_delay_12_18 <= io_A_Valid_7_delay_11_19;
    io_A_Valid_7_delay_13_17 <= io_A_Valid_7_delay_12_18;
    io_A_Valid_7_delay_14_16 <= io_A_Valid_7_delay_13_17;
    io_A_Valid_7_delay_15_15 <= io_A_Valid_7_delay_14_16;
    io_A_Valid_7_delay_16_14 <= io_A_Valid_7_delay_15_15;
    io_A_Valid_7_delay_17_13 <= io_A_Valid_7_delay_16_14;
    io_A_Valid_7_delay_18_12 <= io_A_Valid_7_delay_17_13;
    io_A_Valid_7_delay_19_11 <= io_A_Valid_7_delay_18_12;
    io_A_Valid_7_delay_20_10 <= io_A_Valid_7_delay_19_11;
    io_A_Valid_7_delay_21_9 <= io_A_Valid_7_delay_20_10;
    io_A_Valid_7_delay_22_8 <= io_A_Valid_7_delay_21_9;
    io_A_Valid_7_delay_23_7 <= io_A_Valid_7_delay_22_8;
    io_A_Valid_7_delay_24_6 <= io_A_Valid_7_delay_23_7;
    io_A_Valid_7_delay_25_5 <= io_A_Valid_7_delay_24_6;
    io_A_Valid_7_delay_26_4 <= io_A_Valid_7_delay_25_5;
    io_A_Valid_7_delay_27_3 <= io_A_Valid_7_delay_26_4;
    io_A_Valid_7_delay_28_2 <= io_A_Valid_7_delay_27_3;
    io_A_Valid_7_delay_29_1 <= io_A_Valid_7_delay_28_2;
    io_A_Valid_7_delay_30 <= io_A_Valid_7_delay_29_1;
    io_B_Valid_30_delay_1_6 <= io_B_Valid_30;
    io_B_Valid_30_delay_2_5 <= io_B_Valid_30_delay_1_6;
    io_B_Valid_30_delay_3_4 <= io_B_Valid_30_delay_2_5;
    io_B_Valid_30_delay_4_3 <= io_B_Valid_30_delay_3_4;
    io_B_Valid_30_delay_5_2 <= io_B_Valid_30_delay_4_3;
    io_B_Valid_30_delay_6_1 <= io_B_Valid_30_delay_5_2;
    io_B_Valid_30_delay_7 <= io_B_Valid_30_delay_6_1;
    io_A_Valid_7_delay_1_30 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_29 <= io_A_Valid_7_delay_1_30;
    io_A_Valid_7_delay_3_28 <= io_A_Valid_7_delay_2_29;
    io_A_Valid_7_delay_4_27 <= io_A_Valid_7_delay_3_28;
    io_A_Valid_7_delay_5_26 <= io_A_Valid_7_delay_4_27;
    io_A_Valid_7_delay_6_25 <= io_A_Valid_7_delay_5_26;
    io_A_Valid_7_delay_7_24 <= io_A_Valid_7_delay_6_25;
    io_A_Valid_7_delay_8_23 <= io_A_Valid_7_delay_7_24;
    io_A_Valid_7_delay_9_22 <= io_A_Valid_7_delay_8_23;
    io_A_Valid_7_delay_10_21 <= io_A_Valid_7_delay_9_22;
    io_A_Valid_7_delay_11_20 <= io_A_Valid_7_delay_10_21;
    io_A_Valid_7_delay_12_19 <= io_A_Valid_7_delay_11_20;
    io_A_Valid_7_delay_13_18 <= io_A_Valid_7_delay_12_19;
    io_A_Valid_7_delay_14_17 <= io_A_Valid_7_delay_13_18;
    io_A_Valid_7_delay_15_16 <= io_A_Valid_7_delay_14_17;
    io_A_Valid_7_delay_16_15 <= io_A_Valid_7_delay_15_16;
    io_A_Valid_7_delay_17_14 <= io_A_Valid_7_delay_16_15;
    io_A_Valid_7_delay_18_13 <= io_A_Valid_7_delay_17_14;
    io_A_Valid_7_delay_19_12 <= io_A_Valid_7_delay_18_13;
    io_A_Valid_7_delay_20_11 <= io_A_Valid_7_delay_19_12;
    io_A_Valid_7_delay_21_10 <= io_A_Valid_7_delay_20_11;
    io_A_Valid_7_delay_22_9 <= io_A_Valid_7_delay_21_10;
    io_A_Valid_7_delay_23_8 <= io_A_Valid_7_delay_22_9;
    io_A_Valid_7_delay_24_7 <= io_A_Valid_7_delay_23_8;
    io_A_Valid_7_delay_25_6 <= io_A_Valid_7_delay_24_7;
    io_A_Valid_7_delay_26_5 <= io_A_Valid_7_delay_25_6;
    io_A_Valid_7_delay_27_4 <= io_A_Valid_7_delay_26_5;
    io_A_Valid_7_delay_28_3 <= io_A_Valid_7_delay_27_4;
    io_A_Valid_7_delay_29_2 <= io_A_Valid_7_delay_28_3;
    io_A_Valid_7_delay_30_1 <= io_A_Valid_7_delay_29_2;
    io_A_Valid_7_delay_31 <= io_A_Valid_7_delay_30_1;
    io_B_Valid_31_delay_1_6 <= io_B_Valid_31;
    io_B_Valid_31_delay_2_5 <= io_B_Valid_31_delay_1_6;
    io_B_Valid_31_delay_3_4 <= io_B_Valid_31_delay_2_5;
    io_B_Valid_31_delay_4_3 <= io_B_Valid_31_delay_3_4;
    io_B_Valid_31_delay_5_2 <= io_B_Valid_31_delay_4_3;
    io_B_Valid_31_delay_6_1 <= io_B_Valid_31_delay_5_2;
    io_B_Valid_31_delay_7 <= io_B_Valid_31_delay_6_1;
    io_A_Valid_7_delay_1_31 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_30 <= io_A_Valid_7_delay_1_31;
    io_A_Valid_7_delay_3_29 <= io_A_Valid_7_delay_2_30;
    io_A_Valid_7_delay_4_28 <= io_A_Valid_7_delay_3_29;
    io_A_Valid_7_delay_5_27 <= io_A_Valid_7_delay_4_28;
    io_A_Valid_7_delay_6_26 <= io_A_Valid_7_delay_5_27;
    io_A_Valid_7_delay_7_25 <= io_A_Valid_7_delay_6_26;
    io_A_Valid_7_delay_8_24 <= io_A_Valid_7_delay_7_25;
    io_A_Valid_7_delay_9_23 <= io_A_Valid_7_delay_8_24;
    io_A_Valid_7_delay_10_22 <= io_A_Valid_7_delay_9_23;
    io_A_Valid_7_delay_11_21 <= io_A_Valid_7_delay_10_22;
    io_A_Valid_7_delay_12_20 <= io_A_Valid_7_delay_11_21;
    io_A_Valid_7_delay_13_19 <= io_A_Valid_7_delay_12_20;
    io_A_Valid_7_delay_14_18 <= io_A_Valid_7_delay_13_19;
    io_A_Valid_7_delay_15_17 <= io_A_Valid_7_delay_14_18;
    io_A_Valid_7_delay_16_16 <= io_A_Valid_7_delay_15_17;
    io_A_Valid_7_delay_17_15 <= io_A_Valid_7_delay_16_16;
    io_A_Valid_7_delay_18_14 <= io_A_Valid_7_delay_17_15;
    io_A_Valid_7_delay_19_13 <= io_A_Valid_7_delay_18_14;
    io_A_Valid_7_delay_20_12 <= io_A_Valid_7_delay_19_13;
    io_A_Valid_7_delay_21_11 <= io_A_Valid_7_delay_20_12;
    io_A_Valid_7_delay_22_10 <= io_A_Valid_7_delay_21_11;
    io_A_Valid_7_delay_23_9 <= io_A_Valid_7_delay_22_10;
    io_A_Valid_7_delay_24_8 <= io_A_Valid_7_delay_23_9;
    io_A_Valid_7_delay_25_7 <= io_A_Valid_7_delay_24_8;
    io_A_Valid_7_delay_26_6 <= io_A_Valid_7_delay_25_7;
    io_A_Valid_7_delay_27_5 <= io_A_Valid_7_delay_26_6;
    io_A_Valid_7_delay_28_4 <= io_A_Valid_7_delay_27_5;
    io_A_Valid_7_delay_29_3 <= io_A_Valid_7_delay_28_4;
    io_A_Valid_7_delay_30_2 <= io_A_Valid_7_delay_29_3;
    io_A_Valid_7_delay_31_1 <= io_A_Valid_7_delay_30_2;
    io_A_Valid_7_delay_32 <= io_A_Valid_7_delay_31_1;
    io_B_Valid_32_delay_1_6 <= io_B_Valid_32;
    io_B_Valid_32_delay_2_5 <= io_B_Valid_32_delay_1_6;
    io_B_Valid_32_delay_3_4 <= io_B_Valid_32_delay_2_5;
    io_B_Valid_32_delay_4_3 <= io_B_Valid_32_delay_3_4;
    io_B_Valid_32_delay_5_2 <= io_B_Valid_32_delay_4_3;
    io_B_Valid_32_delay_6_1 <= io_B_Valid_32_delay_5_2;
    io_B_Valid_32_delay_7 <= io_B_Valid_32_delay_6_1;
    io_A_Valid_7_delay_1_32 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_31 <= io_A_Valid_7_delay_1_32;
    io_A_Valid_7_delay_3_30 <= io_A_Valid_7_delay_2_31;
    io_A_Valid_7_delay_4_29 <= io_A_Valid_7_delay_3_30;
    io_A_Valid_7_delay_5_28 <= io_A_Valid_7_delay_4_29;
    io_A_Valid_7_delay_6_27 <= io_A_Valid_7_delay_5_28;
    io_A_Valid_7_delay_7_26 <= io_A_Valid_7_delay_6_27;
    io_A_Valid_7_delay_8_25 <= io_A_Valid_7_delay_7_26;
    io_A_Valid_7_delay_9_24 <= io_A_Valid_7_delay_8_25;
    io_A_Valid_7_delay_10_23 <= io_A_Valid_7_delay_9_24;
    io_A_Valid_7_delay_11_22 <= io_A_Valid_7_delay_10_23;
    io_A_Valid_7_delay_12_21 <= io_A_Valid_7_delay_11_22;
    io_A_Valid_7_delay_13_20 <= io_A_Valid_7_delay_12_21;
    io_A_Valid_7_delay_14_19 <= io_A_Valid_7_delay_13_20;
    io_A_Valid_7_delay_15_18 <= io_A_Valid_7_delay_14_19;
    io_A_Valid_7_delay_16_17 <= io_A_Valid_7_delay_15_18;
    io_A_Valid_7_delay_17_16 <= io_A_Valid_7_delay_16_17;
    io_A_Valid_7_delay_18_15 <= io_A_Valid_7_delay_17_16;
    io_A_Valid_7_delay_19_14 <= io_A_Valid_7_delay_18_15;
    io_A_Valid_7_delay_20_13 <= io_A_Valid_7_delay_19_14;
    io_A_Valid_7_delay_21_12 <= io_A_Valid_7_delay_20_13;
    io_A_Valid_7_delay_22_11 <= io_A_Valid_7_delay_21_12;
    io_A_Valid_7_delay_23_10 <= io_A_Valid_7_delay_22_11;
    io_A_Valid_7_delay_24_9 <= io_A_Valid_7_delay_23_10;
    io_A_Valid_7_delay_25_8 <= io_A_Valid_7_delay_24_9;
    io_A_Valid_7_delay_26_7 <= io_A_Valid_7_delay_25_8;
    io_A_Valid_7_delay_27_6 <= io_A_Valid_7_delay_26_7;
    io_A_Valid_7_delay_28_5 <= io_A_Valid_7_delay_27_6;
    io_A_Valid_7_delay_29_4 <= io_A_Valid_7_delay_28_5;
    io_A_Valid_7_delay_30_3 <= io_A_Valid_7_delay_29_4;
    io_A_Valid_7_delay_31_2 <= io_A_Valid_7_delay_30_3;
    io_A_Valid_7_delay_32_1 <= io_A_Valid_7_delay_31_2;
    io_A_Valid_7_delay_33 <= io_A_Valid_7_delay_32_1;
    io_B_Valid_33_delay_1_6 <= io_B_Valid_33;
    io_B_Valid_33_delay_2_5 <= io_B_Valid_33_delay_1_6;
    io_B_Valid_33_delay_3_4 <= io_B_Valid_33_delay_2_5;
    io_B_Valid_33_delay_4_3 <= io_B_Valid_33_delay_3_4;
    io_B_Valid_33_delay_5_2 <= io_B_Valid_33_delay_4_3;
    io_B_Valid_33_delay_6_1 <= io_B_Valid_33_delay_5_2;
    io_B_Valid_33_delay_7 <= io_B_Valid_33_delay_6_1;
    io_A_Valid_7_delay_1_33 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_32 <= io_A_Valid_7_delay_1_33;
    io_A_Valid_7_delay_3_31 <= io_A_Valid_7_delay_2_32;
    io_A_Valid_7_delay_4_30 <= io_A_Valid_7_delay_3_31;
    io_A_Valid_7_delay_5_29 <= io_A_Valid_7_delay_4_30;
    io_A_Valid_7_delay_6_28 <= io_A_Valid_7_delay_5_29;
    io_A_Valid_7_delay_7_27 <= io_A_Valid_7_delay_6_28;
    io_A_Valid_7_delay_8_26 <= io_A_Valid_7_delay_7_27;
    io_A_Valid_7_delay_9_25 <= io_A_Valid_7_delay_8_26;
    io_A_Valid_7_delay_10_24 <= io_A_Valid_7_delay_9_25;
    io_A_Valid_7_delay_11_23 <= io_A_Valid_7_delay_10_24;
    io_A_Valid_7_delay_12_22 <= io_A_Valid_7_delay_11_23;
    io_A_Valid_7_delay_13_21 <= io_A_Valid_7_delay_12_22;
    io_A_Valid_7_delay_14_20 <= io_A_Valid_7_delay_13_21;
    io_A_Valid_7_delay_15_19 <= io_A_Valid_7_delay_14_20;
    io_A_Valid_7_delay_16_18 <= io_A_Valid_7_delay_15_19;
    io_A_Valid_7_delay_17_17 <= io_A_Valid_7_delay_16_18;
    io_A_Valid_7_delay_18_16 <= io_A_Valid_7_delay_17_17;
    io_A_Valid_7_delay_19_15 <= io_A_Valid_7_delay_18_16;
    io_A_Valid_7_delay_20_14 <= io_A_Valid_7_delay_19_15;
    io_A_Valid_7_delay_21_13 <= io_A_Valid_7_delay_20_14;
    io_A_Valid_7_delay_22_12 <= io_A_Valid_7_delay_21_13;
    io_A_Valid_7_delay_23_11 <= io_A_Valid_7_delay_22_12;
    io_A_Valid_7_delay_24_10 <= io_A_Valid_7_delay_23_11;
    io_A_Valid_7_delay_25_9 <= io_A_Valid_7_delay_24_10;
    io_A_Valid_7_delay_26_8 <= io_A_Valid_7_delay_25_9;
    io_A_Valid_7_delay_27_7 <= io_A_Valid_7_delay_26_8;
    io_A_Valid_7_delay_28_6 <= io_A_Valid_7_delay_27_7;
    io_A_Valid_7_delay_29_5 <= io_A_Valid_7_delay_28_6;
    io_A_Valid_7_delay_30_4 <= io_A_Valid_7_delay_29_5;
    io_A_Valid_7_delay_31_3 <= io_A_Valid_7_delay_30_4;
    io_A_Valid_7_delay_32_2 <= io_A_Valid_7_delay_31_3;
    io_A_Valid_7_delay_33_1 <= io_A_Valid_7_delay_32_2;
    io_A_Valid_7_delay_34 <= io_A_Valid_7_delay_33_1;
    io_B_Valid_34_delay_1_6 <= io_B_Valid_34;
    io_B_Valid_34_delay_2_5 <= io_B_Valid_34_delay_1_6;
    io_B_Valid_34_delay_3_4 <= io_B_Valid_34_delay_2_5;
    io_B_Valid_34_delay_4_3 <= io_B_Valid_34_delay_3_4;
    io_B_Valid_34_delay_5_2 <= io_B_Valid_34_delay_4_3;
    io_B_Valid_34_delay_6_1 <= io_B_Valid_34_delay_5_2;
    io_B_Valid_34_delay_7 <= io_B_Valid_34_delay_6_1;
    io_A_Valid_7_delay_1_34 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_33 <= io_A_Valid_7_delay_1_34;
    io_A_Valid_7_delay_3_32 <= io_A_Valid_7_delay_2_33;
    io_A_Valid_7_delay_4_31 <= io_A_Valid_7_delay_3_32;
    io_A_Valid_7_delay_5_30 <= io_A_Valid_7_delay_4_31;
    io_A_Valid_7_delay_6_29 <= io_A_Valid_7_delay_5_30;
    io_A_Valid_7_delay_7_28 <= io_A_Valid_7_delay_6_29;
    io_A_Valid_7_delay_8_27 <= io_A_Valid_7_delay_7_28;
    io_A_Valid_7_delay_9_26 <= io_A_Valid_7_delay_8_27;
    io_A_Valid_7_delay_10_25 <= io_A_Valid_7_delay_9_26;
    io_A_Valid_7_delay_11_24 <= io_A_Valid_7_delay_10_25;
    io_A_Valid_7_delay_12_23 <= io_A_Valid_7_delay_11_24;
    io_A_Valid_7_delay_13_22 <= io_A_Valid_7_delay_12_23;
    io_A_Valid_7_delay_14_21 <= io_A_Valid_7_delay_13_22;
    io_A_Valid_7_delay_15_20 <= io_A_Valid_7_delay_14_21;
    io_A_Valid_7_delay_16_19 <= io_A_Valid_7_delay_15_20;
    io_A_Valid_7_delay_17_18 <= io_A_Valid_7_delay_16_19;
    io_A_Valid_7_delay_18_17 <= io_A_Valid_7_delay_17_18;
    io_A_Valid_7_delay_19_16 <= io_A_Valid_7_delay_18_17;
    io_A_Valid_7_delay_20_15 <= io_A_Valid_7_delay_19_16;
    io_A_Valid_7_delay_21_14 <= io_A_Valid_7_delay_20_15;
    io_A_Valid_7_delay_22_13 <= io_A_Valid_7_delay_21_14;
    io_A_Valid_7_delay_23_12 <= io_A_Valid_7_delay_22_13;
    io_A_Valid_7_delay_24_11 <= io_A_Valid_7_delay_23_12;
    io_A_Valid_7_delay_25_10 <= io_A_Valid_7_delay_24_11;
    io_A_Valid_7_delay_26_9 <= io_A_Valid_7_delay_25_10;
    io_A_Valid_7_delay_27_8 <= io_A_Valid_7_delay_26_9;
    io_A_Valid_7_delay_28_7 <= io_A_Valid_7_delay_27_8;
    io_A_Valid_7_delay_29_6 <= io_A_Valid_7_delay_28_7;
    io_A_Valid_7_delay_30_5 <= io_A_Valid_7_delay_29_6;
    io_A_Valid_7_delay_31_4 <= io_A_Valid_7_delay_30_5;
    io_A_Valid_7_delay_32_3 <= io_A_Valid_7_delay_31_4;
    io_A_Valid_7_delay_33_2 <= io_A_Valid_7_delay_32_3;
    io_A_Valid_7_delay_34_1 <= io_A_Valid_7_delay_33_2;
    io_A_Valid_7_delay_35 <= io_A_Valid_7_delay_34_1;
    io_B_Valid_35_delay_1_6 <= io_B_Valid_35;
    io_B_Valid_35_delay_2_5 <= io_B_Valid_35_delay_1_6;
    io_B_Valid_35_delay_3_4 <= io_B_Valid_35_delay_2_5;
    io_B_Valid_35_delay_4_3 <= io_B_Valid_35_delay_3_4;
    io_B_Valid_35_delay_5_2 <= io_B_Valid_35_delay_4_3;
    io_B_Valid_35_delay_6_1 <= io_B_Valid_35_delay_5_2;
    io_B_Valid_35_delay_7 <= io_B_Valid_35_delay_6_1;
    io_A_Valid_7_delay_1_35 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_34 <= io_A_Valid_7_delay_1_35;
    io_A_Valid_7_delay_3_33 <= io_A_Valid_7_delay_2_34;
    io_A_Valid_7_delay_4_32 <= io_A_Valid_7_delay_3_33;
    io_A_Valid_7_delay_5_31 <= io_A_Valid_7_delay_4_32;
    io_A_Valid_7_delay_6_30 <= io_A_Valid_7_delay_5_31;
    io_A_Valid_7_delay_7_29 <= io_A_Valid_7_delay_6_30;
    io_A_Valid_7_delay_8_28 <= io_A_Valid_7_delay_7_29;
    io_A_Valid_7_delay_9_27 <= io_A_Valid_7_delay_8_28;
    io_A_Valid_7_delay_10_26 <= io_A_Valid_7_delay_9_27;
    io_A_Valid_7_delay_11_25 <= io_A_Valid_7_delay_10_26;
    io_A_Valid_7_delay_12_24 <= io_A_Valid_7_delay_11_25;
    io_A_Valid_7_delay_13_23 <= io_A_Valid_7_delay_12_24;
    io_A_Valid_7_delay_14_22 <= io_A_Valid_7_delay_13_23;
    io_A_Valid_7_delay_15_21 <= io_A_Valid_7_delay_14_22;
    io_A_Valid_7_delay_16_20 <= io_A_Valid_7_delay_15_21;
    io_A_Valid_7_delay_17_19 <= io_A_Valid_7_delay_16_20;
    io_A_Valid_7_delay_18_18 <= io_A_Valid_7_delay_17_19;
    io_A_Valid_7_delay_19_17 <= io_A_Valid_7_delay_18_18;
    io_A_Valid_7_delay_20_16 <= io_A_Valid_7_delay_19_17;
    io_A_Valid_7_delay_21_15 <= io_A_Valid_7_delay_20_16;
    io_A_Valid_7_delay_22_14 <= io_A_Valid_7_delay_21_15;
    io_A_Valid_7_delay_23_13 <= io_A_Valid_7_delay_22_14;
    io_A_Valid_7_delay_24_12 <= io_A_Valid_7_delay_23_13;
    io_A_Valid_7_delay_25_11 <= io_A_Valid_7_delay_24_12;
    io_A_Valid_7_delay_26_10 <= io_A_Valid_7_delay_25_11;
    io_A_Valid_7_delay_27_9 <= io_A_Valid_7_delay_26_10;
    io_A_Valid_7_delay_28_8 <= io_A_Valid_7_delay_27_9;
    io_A_Valid_7_delay_29_7 <= io_A_Valid_7_delay_28_8;
    io_A_Valid_7_delay_30_6 <= io_A_Valid_7_delay_29_7;
    io_A_Valid_7_delay_31_5 <= io_A_Valid_7_delay_30_6;
    io_A_Valid_7_delay_32_4 <= io_A_Valid_7_delay_31_5;
    io_A_Valid_7_delay_33_3 <= io_A_Valid_7_delay_32_4;
    io_A_Valid_7_delay_34_2 <= io_A_Valid_7_delay_33_3;
    io_A_Valid_7_delay_35_1 <= io_A_Valid_7_delay_34_2;
    io_A_Valid_7_delay_36 <= io_A_Valid_7_delay_35_1;
    io_B_Valid_36_delay_1_6 <= io_B_Valid_36;
    io_B_Valid_36_delay_2_5 <= io_B_Valid_36_delay_1_6;
    io_B_Valid_36_delay_3_4 <= io_B_Valid_36_delay_2_5;
    io_B_Valid_36_delay_4_3 <= io_B_Valid_36_delay_3_4;
    io_B_Valid_36_delay_5_2 <= io_B_Valid_36_delay_4_3;
    io_B_Valid_36_delay_6_1 <= io_B_Valid_36_delay_5_2;
    io_B_Valid_36_delay_7 <= io_B_Valid_36_delay_6_1;
    io_A_Valid_7_delay_1_36 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_35 <= io_A_Valid_7_delay_1_36;
    io_A_Valid_7_delay_3_34 <= io_A_Valid_7_delay_2_35;
    io_A_Valid_7_delay_4_33 <= io_A_Valid_7_delay_3_34;
    io_A_Valid_7_delay_5_32 <= io_A_Valid_7_delay_4_33;
    io_A_Valid_7_delay_6_31 <= io_A_Valid_7_delay_5_32;
    io_A_Valid_7_delay_7_30 <= io_A_Valid_7_delay_6_31;
    io_A_Valid_7_delay_8_29 <= io_A_Valid_7_delay_7_30;
    io_A_Valid_7_delay_9_28 <= io_A_Valid_7_delay_8_29;
    io_A_Valid_7_delay_10_27 <= io_A_Valid_7_delay_9_28;
    io_A_Valid_7_delay_11_26 <= io_A_Valid_7_delay_10_27;
    io_A_Valid_7_delay_12_25 <= io_A_Valid_7_delay_11_26;
    io_A_Valid_7_delay_13_24 <= io_A_Valid_7_delay_12_25;
    io_A_Valid_7_delay_14_23 <= io_A_Valid_7_delay_13_24;
    io_A_Valid_7_delay_15_22 <= io_A_Valid_7_delay_14_23;
    io_A_Valid_7_delay_16_21 <= io_A_Valid_7_delay_15_22;
    io_A_Valid_7_delay_17_20 <= io_A_Valid_7_delay_16_21;
    io_A_Valid_7_delay_18_19 <= io_A_Valid_7_delay_17_20;
    io_A_Valid_7_delay_19_18 <= io_A_Valid_7_delay_18_19;
    io_A_Valid_7_delay_20_17 <= io_A_Valid_7_delay_19_18;
    io_A_Valid_7_delay_21_16 <= io_A_Valid_7_delay_20_17;
    io_A_Valid_7_delay_22_15 <= io_A_Valid_7_delay_21_16;
    io_A_Valid_7_delay_23_14 <= io_A_Valid_7_delay_22_15;
    io_A_Valid_7_delay_24_13 <= io_A_Valid_7_delay_23_14;
    io_A_Valid_7_delay_25_12 <= io_A_Valid_7_delay_24_13;
    io_A_Valid_7_delay_26_11 <= io_A_Valid_7_delay_25_12;
    io_A_Valid_7_delay_27_10 <= io_A_Valid_7_delay_26_11;
    io_A_Valid_7_delay_28_9 <= io_A_Valid_7_delay_27_10;
    io_A_Valid_7_delay_29_8 <= io_A_Valid_7_delay_28_9;
    io_A_Valid_7_delay_30_7 <= io_A_Valid_7_delay_29_8;
    io_A_Valid_7_delay_31_6 <= io_A_Valid_7_delay_30_7;
    io_A_Valid_7_delay_32_5 <= io_A_Valid_7_delay_31_6;
    io_A_Valid_7_delay_33_4 <= io_A_Valid_7_delay_32_5;
    io_A_Valid_7_delay_34_3 <= io_A_Valid_7_delay_33_4;
    io_A_Valid_7_delay_35_2 <= io_A_Valid_7_delay_34_3;
    io_A_Valid_7_delay_36_1 <= io_A_Valid_7_delay_35_2;
    io_A_Valid_7_delay_37 <= io_A_Valid_7_delay_36_1;
    io_B_Valid_37_delay_1_6 <= io_B_Valid_37;
    io_B_Valid_37_delay_2_5 <= io_B_Valid_37_delay_1_6;
    io_B_Valid_37_delay_3_4 <= io_B_Valid_37_delay_2_5;
    io_B_Valid_37_delay_4_3 <= io_B_Valid_37_delay_3_4;
    io_B_Valid_37_delay_5_2 <= io_B_Valid_37_delay_4_3;
    io_B_Valid_37_delay_6_1 <= io_B_Valid_37_delay_5_2;
    io_B_Valid_37_delay_7 <= io_B_Valid_37_delay_6_1;
    io_A_Valid_7_delay_1_37 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_36 <= io_A_Valid_7_delay_1_37;
    io_A_Valid_7_delay_3_35 <= io_A_Valid_7_delay_2_36;
    io_A_Valid_7_delay_4_34 <= io_A_Valid_7_delay_3_35;
    io_A_Valid_7_delay_5_33 <= io_A_Valid_7_delay_4_34;
    io_A_Valid_7_delay_6_32 <= io_A_Valid_7_delay_5_33;
    io_A_Valid_7_delay_7_31 <= io_A_Valid_7_delay_6_32;
    io_A_Valid_7_delay_8_30 <= io_A_Valid_7_delay_7_31;
    io_A_Valid_7_delay_9_29 <= io_A_Valid_7_delay_8_30;
    io_A_Valid_7_delay_10_28 <= io_A_Valid_7_delay_9_29;
    io_A_Valid_7_delay_11_27 <= io_A_Valid_7_delay_10_28;
    io_A_Valid_7_delay_12_26 <= io_A_Valid_7_delay_11_27;
    io_A_Valid_7_delay_13_25 <= io_A_Valid_7_delay_12_26;
    io_A_Valid_7_delay_14_24 <= io_A_Valid_7_delay_13_25;
    io_A_Valid_7_delay_15_23 <= io_A_Valid_7_delay_14_24;
    io_A_Valid_7_delay_16_22 <= io_A_Valid_7_delay_15_23;
    io_A_Valid_7_delay_17_21 <= io_A_Valid_7_delay_16_22;
    io_A_Valid_7_delay_18_20 <= io_A_Valid_7_delay_17_21;
    io_A_Valid_7_delay_19_19 <= io_A_Valid_7_delay_18_20;
    io_A_Valid_7_delay_20_18 <= io_A_Valid_7_delay_19_19;
    io_A_Valid_7_delay_21_17 <= io_A_Valid_7_delay_20_18;
    io_A_Valid_7_delay_22_16 <= io_A_Valid_7_delay_21_17;
    io_A_Valid_7_delay_23_15 <= io_A_Valid_7_delay_22_16;
    io_A_Valid_7_delay_24_14 <= io_A_Valid_7_delay_23_15;
    io_A_Valid_7_delay_25_13 <= io_A_Valid_7_delay_24_14;
    io_A_Valid_7_delay_26_12 <= io_A_Valid_7_delay_25_13;
    io_A_Valid_7_delay_27_11 <= io_A_Valid_7_delay_26_12;
    io_A_Valid_7_delay_28_10 <= io_A_Valid_7_delay_27_11;
    io_A_Valid_7_delay_29_9 <= io_A_Valid_7_delay_28_10;
    io_A_Valid_7_delay_30_8 <= io_A_Valid_7_delay_29_9;
    io_A_Valid_7_delay_31_7 <= io_A_Valid_7_delay_30_8;
    io_A_Valid_7_delay_32_6 <= io_A_Valid_7_delay_31_7;
    io_A_Valid_7_delay_33_5 <= io_A_Valid_7_delay_32_6;
    io_A_Valid_7_delay_34_4 <= io_A_Valid_7_delay_33_5;
    io_A_Valid_7_delay_35_3 <= io_A_Valid_7_delay_34_4;
    io_A_Valid_7_delay_36_2 <= io_A_Valid_7_delay_35_3;
    io_A_Valid_7_delay_37_1 <= io_A_Valid_7_delay_36_2;
    io_A_Valid_7_delay_38 <= io_A_Valid_7_delay_37_1;
    io_B_Valid_38_delay_1_6 <= io_B_Valid_38;
    io_B_Valid_38_delay_2_5 <= io_B_Valid_38_delay_1_6;
    io_B_Valid_38_delay_3_4 <= io_B_Valid_38_delay_2_5;
    io_B_Valid_38_delay_4_3 <= io_B_Valid_38_delay_3_4;
    io_B_Valid_38_delay_5_2 <= io_B_Valid_38_delay_4_3;
    io_B_Valid_38_delay_6_1 <= io_B_Valid_38_delay_5_2;
    io_B_Valid_38_delay_7 <= io_B_Valid_38_delay_6_1;
    io_A_Valid_7_delay_1_38 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_37 <= io_A_Valid_7_delay_1_38;
    io_A_Valid_7_delay_3_36 <= io_A_Valid_7_delay_2_37;
    io_A_Valid_7_delay_4_35 <= io_A_Valid_7_delay_3_36;
    io_A_Valid_7_delay_5_34 <= io_A_Valid_7_delay_4_35;
    io_A_Valid_7_delay_6_33 <= io_A_Valid_7_delay_5_34;
    io_A_Valid_7_delay_7_32 <= io_A_Valid_7_delay_6_33;
    io_A_Valid_7_delay_8_31 <= io_A_Valid_7_delay_7_32;
    io_A_Valid_7_delay_9_30 <= io_A_Valid_7_delay_8_31;
    io_A_Valid_7_delay_10_29 <= io_A_Valid_7_delay_9_30;
    io_A_Valid_7_delay_11_28 <= io_A_Valid_7_delay_10_29;
    io_A_Valid_7_delay_12_27 <= io_A_Valid_7_delay_11_28;
    io_A_Valid_7_delay_13_26 <= io_A_Valid_7_delay_12_27;
    io_A_Valid_7_delay_14_25 <= io_A_Valid_7_delay_13_26;
    io_A_Valid_7_delay_15_24 <= io_A_Valid_7_delay_14_25;
    io_A_Valid_7_delay_16_23 <= io_A_Valid_7_delay_15_24;
    io_A_Valid_7_delay_17_22 <= io_A_Valid_7_delay_16_23;
    io_A_Valid_7_delay_18_21 <= io_A_Valid_7_delay_17_22;
    io_A_Valid_7_delay_19_20 <= io_A_Valid_7_delay_18_21;
    io_A_Valid_7_delay_20_19 <= io_A_Valid_7_delay_19_20;
    io_A_Valid_7_delay_21_18 <= io_A_Valid_7_delay_20_19;
    io_A_Valid_7_delay_22_17 <= io_A_Valid_7_delay_21_18;
    io_A_Valid_7_delay_23_16 <= io_A_Valid_7_delay_22_17;
    io_A_Valid_7_delay_24_15 <= io_A_Valid_7_delay_23_16;
    io_A_Valid_7_delay_25_14 <= io_A_Valid_7_delay_24_15;
    io_A_Valid_7_delay_26_13 <= io_A_Valid_7_delay_25_14;
    io_A_Valid_7_delay_27_12 <= io_A_Valid_7_delay_26_13;
    io_A_Valid_7_delay_28_11 <= io_A_Valid_7_delay_27_12;
    io_A_Valid_7_delay_29_10 <= io_A_Valid_7_delay_28_11;
    io_A_Valid_7_delay_30_9 <= io_A_Valid_7_delay_29_10;
    io_A_Valid_7_delay_31_8 <= io_A_Valid_7_delay_30_9;
    io_A_Valid_7_delay_32_7 <= io_A_Valid_7_delay_31_8;
    io_A_Valid_7_delay_33_6 <= io_A_Valid_7_delay_32_7;
    io_A_Valid_7_delay_34_5 <= io_A_Valid_7_delay_33_6;
    io_A_Valid_7_delay_35_4 <= io_A_Valid_7_delay_34_5;
    io_A_Valid_7_delay_36_3 <= io_A_Valid_7_delay_35_4;
    io_A_Valid_7_delay_37_2 <= io_A_Valid_7_delay_36_3;
    io_A_Valid_7_delay_38_1 <= io_A_Valid_7_delay_37_2;
    io_A_Valid_7_delay_39 <= io_A_Valid_7_delay_38_1;
    io_B_Valid_39_delay_1_6 <= io_B_Valid_39;
    io_B_Valid_39_delay_2_5 <= io_B_Valid_39_delay_1_6;
    io_B_Valid_39_delay_3_4 <= io_B_Valid_39_delay_2_5;
    io_B_Valid_39_delay_4_3 <= io_B_Valid_39_delay_3_4;
    io_B_Valid_39_delay_5_2 <= io_B_Valid_39_delay_4_3;
    io_B_Valid_39_delay_6_1 <= io_B_Valid_39_delay_5_2;
    io_B_Valid_39_delay_7 <= io_B_Valid_39_delay_6_1;
    io_A_Valid_7_delay_1_39 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_38 <= io_A_Valid_7_delay_1_39;
    io_A_Valid_7_delay_3_37 <= io_A_Valid_7_delay_2_38;
    io_A_Valid_7_delay_4_36 <= io_A_Valid_7_delay_3_37;
    io_A_Valid_7_delay_5_35 <= io_A_Valid_7_delay_4_36;
    io_A_Valid_7_delay_6_34 <= io_A_Valid_7_delay_5_35;
    io_A_Valid_7_delay_7_33 <= io_A_Valid_7_delay_6_34;
    io_A_Valid_7_delay_8_32 <= io_A_Valid_7_delay_7_33;
    io_A_Valid_7_delay_9_31 <= io_A_Valid_7_delay_8_32;
    io_A_Valid_7_delay_10_30 <= io_A_Valid_7_delay_9_31;
    io_A_Valid_7_delay_11_29 <= io_A_Valid_7_delay_10_30;
    io_A_Valid_7_delay_12_28 <= io_A_Valid_7_delay_11_29;
    io_A_Valid_7_delay_13_27 <= io_A_Valid_7_delay_12_28;
    io_A_Valid_7_delay_14_26 <= io_A_Valid_7_delay_13_27;
    io_A_Valid_7_delay_15_25 <= io_A_Valid_7_delay_14_26;
    io_A_Valid_7_delay_16_24 <= io_A_Valid_7_delay_15_25;
    io_A_Valid_7_delay_17_23 <= io_A_Valid_7_delay_16_24;
    io_A_Valid_7_delay_18_22 <= io_A_Valid_7_delay_17_23;
    io_A_Valid_7_delay_19_21 <= io_A_Valid_7_delay_18_22;
    io_A_Valid_7_delay_20_20 <= io_A_Valid_7_delay_19_21;
    io_A_Valid_7_delay_21_19 <= io_A_Valid_7_delay_20_20;
    io_A_Valid_7_delay_22_18 <= io_A_Valid_7_delay_21_19;
    io_A_Valid_7_delay_23_17 <= io_A_Valid_7_delay_22_18;
    io_A_Valid_7_delay_24_16 <= io_A_Valid_7_delay_23_17;
    io_A_Valid_7_delay_25_15 <= io_A_Valid_7_delay_24_16;
    io_A_Valid_7_delay_26_14 <= io_A_Valid_7_delay_25_15;
    io_A_Valid_7_delay_27_13 <= io_A_Valid_7_delay_26_14;
    io_A_Valid_7_delay_28_12 <= io_A_Valid_7_delay_27_13;
    io_A_Valid_7_delay_29_11 <= io_A_Valid_7_delay_28_12;
    io_A_Valid_7_delay_30_10 <= io_A_Valid_7_delay_29_11;
    io_A_Valid_7_delay_31_9 <= io_A_Valid_7_delay_30_10;
    io_A_Valid_7_delay_32_8 <= io_A_Valid_7_delay_31_9;
    io_A_Valid_7_delay_33_7 <= io_A_Valid_7_delay_32_8;
    io_A_Valid_7_delay_34_6 <= io_A_Valid_7_delay_33_7;
    io_A_Valid_7_delay_35_5 <= io_A_Valid_7_delay_34_6;
    io_A_Valid_7_delay_36_4 <= io_A_Valid_7_delay_35_5;
    io_A_Valid_7_delay_37_3 <= io_A_Valid_7_delay_36_4;
    io_A_Valid_7_delay_38_2 <= io_A_Valid_7_delay_37_3;
    io_A_Valid_7_delay_39_1 <= io_A_Valid_7_delay_38_2;
    io_A_Valid_7_delay_40 <= io_A_Valid_7_delay_39_1;
    io_B_Valid_40_delay_1_6 <= io_B_Valid_40;
    io_B_Valid_40_delay_2_5 <= io_B_Valid_40_delay_1_6;
    io_B_Valid_40_delay_3_4 <= io_B_Valid_40_delay_2_5;
    io_B_Valid_40_delay_4_3 <= io_B_Valid_40_delay_3_4;
    io_B_Valid_40_delay_5_2 <= io_B_Valid_40_delay_4_3;
    io_B_Valid_40_delay_6_1 <= io_B_Valid_40_delay_5_2;
    io_B_Valid_40_delay_7 <= io_B_Valid_40_delay_6_1;
    io_A_Valid_7_delay_1_40 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_39 <= io_A_Valid_7_delay_1_40;
    io_A_Valid_7_delay_3_38 <= io_A_Valid_7_delay_2_39;
    io_A_Valid_7_delay_4_37 <= io_A_Valid_7_delay_3_38;
    io_A_Valid_7_delay_5_36 <= io_A_Valid_7_delay_4_37;
    io_A_Valid_7_delay_6_35 <= io_A_Valid_7_delay_5_36;
    io_A_Valid_7_delay_7_34 <= io_A_Valid_7_delay_6_35;
    io_A_Valid_7_delay_8_33 <= io_A_Valid_7_delay_7_34;
    io_A_Valid_7_delay_9_32 <= io_A_Valid_7_delay_8_33;
    io_A_Valid_7_delay_10_31 <= io_A_Valid_7_delay_9_32;
    io_A_Valid_7_delay_11_30 <= io_A_Valid_7_delay_10_31;
    io_A_Valid_7_delay_12_29 <= io_A_Valid_7_delay_11_30;
    io_A_Valid_7_delay_13_28 <= io_A_Valid_7_delay_12_29;
    io_A_Valid_7_delay_14_27 <= io_A_Valid_7_delay_13_28;
    io_A_Valid_7_delay_15_26 <= io_A_Valid_7_delay_14_27;
    io_A_Valid_7_delay_16_25 <= io_A_Valid_7_delay_15_26;
    io_A_Valid_7_delay_17_24 <= io_A_Valid_7_delay_16_25;
    io_A_Valid_7_delay_18_23 <= io_A_Valid_7_delay_17_24;
    io_A_Valid_7_delay_19_22 <= io_A_Valid_7_delay_18_23;
    io_A_Valid_7_delay_20_21 <= io_A_Valid_7_delay_19_22;
    io_A_Valid_7_delay_21_20 <= io_A_Valid_7_delay_20_21;
    io_A_Valid_7_delay_22_19 <= io_A_Valid_7_delay_21_20;
    io_A_Valid_7_delay_23_18 <= io_A_Valid_7_delay_22_19;
    io_A_Valid_7_delay_24_17 <= io_A_Valid_7_delay_23_18;
    io_A_Valid_7_delay_25_16 <= io_A_Valid_7_delay_24_17;
    io_A_Valid_7_delay_26_15 <= io_A_Valid_7_delay_25_16;
    io_A_Valid_7_delay_27_14 <= io_A_Valid_7_delay_26_15;
    io_A_Valid_7_delay_28_13 <= io_A_Valid_7_delay_27_14;
    io_A_Valid_7_delay_29_12 <= io_A_Valid_7_delay_28_13;
    io_A_Valid_7_delay_30_11 <= io_A_Valid_7_delay_29_12;
    io_A_Valid_7_delay_31_10 <= io_A_Valid_7_delay_30_11;
    io_A_Valid_7_delay_32_9 <= io_A_Valid_7_delay_31_10;
    io_A_Valid_7_delay_33_8 <= io_A_Valid_7_delay_32_9;
    io_A_Valid_7_delay_34_7 <= io_A_Valid_7_delay_33_8;
    io_A_Valid_7_delay_35_6 <= io_A_Valid_7_delay_34_7;
    io_A_Valid_7_delay_36_5 <= io_A_Valid_7_delay_35_6;
    io_A_Valid_7_delay_37_4 <= io_A_Valid_7_delay_36_5;
    io_A_Valid_7_delay_38_3 <= io_A_Valid_7_delay_37_4;
    io_A_Valid_7_delay_39_2 <= io_A_Valid_7_delay_38_3;
    io_A_Valid_7_delay_40_1 <= io_A_Valid_7_delay_39_2;
    io_A_Valid_7_delay_41 <= io_A_Valid_7_delay_40_1;
    io_B_Valid_41_delay_1_6 <= io_B_Valid_41;
    io_B_Valid_41_delay_2_5 <= io_B_Valid_41_delay_1_6;
    io_B_Valid_41_delay_3_4 <= io_B_Valid_41_delay_2_5;
    io_B_Valid_41_delay_4_3 <= io_B_Valid_41_delay_3_4;
    io_B_Valid_41_delay_5_2 <= io_B_Valid_41_delay_4_3;
    io_B_Valid_41_delay_6_1 <= io_B_Valid_41_delay_5_2;
    io_B_Valid_41_delay_7 <= io_B_Valid_41_delay_6_1;
    io_A_Valid_7_delay_1_41 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_40 <= io_A_Valid_7_delay_1_41;
    io_A_Valid_7_delay_3_39 <= io_A_Valid_7_delay_2_40;
    io_A_Valid_7_delay_4_38 <= io_A_Valid_7_delay_3_39;
    io_A_Valid_7_delay_5_37 <= io_A_Valid_7_delay_4_38;
    io_A_Valid_7_delay_6_36 <= io_A_Valid_7_delay_5_37;
    io_A_Valid_7_delay_7_35 <= io_A_Valid_7_delay_6_36;
    io_A_Valid_7_delay_8_34 <= io_A_Valid_7_delay_7_35;
    io_A_Valid_7_delay_9_33 <= io_A_Valid_7_delay_8_34;
    io_A_Valid_7_delay_10_32 <= io_A_Valid_7_delay_9_33;
    io_A_Valid_7_delay_11_31 <= io_A_Valid_7_delay_10_32;
    io_A_Valid_7_delay_12_30 <= io_A_Valid_7_delay_11_31;
    io_A_Valid_7_delay_13_29 <= io_A_Valid_7_delay_12_30;
    io_A_Valid_7_delay_14_28 <= io_A_Valid_7_delay_13_29;
    io_A_Valid_7_delay_15_27 <= io_A_Valid_7_delay_14_28;
    io_A_Valid_7_delay_16_26 <= io_A_Valid_7_delay_15_27;
    io_A_Valid_7_delay_17_25 <= io_A_Valid_7_delay_16_26;
    io_A_Valid_7_delay_18_24 <= io_A_Valid_7_delay_17_25;
    io_A_Valid_7_delay_19_23 <= io_A_Valid_7_delay_18_24;
    io_A_Valid_7_delay_20_22 <= io_A_Valid_7_delay_19_23;
    io_A_Valid_7_delay_21_21 <= io_A_Valid_7_delay_20_22;
    io_A_Valid_7_delay_22_20 <= io_A_Valid_7_delay_21_21;
    io_A_Valid_7_delay_23_19 <= io_A_Valid_7_delay_22_20;
    io_A_Valid_7_delay_24_18 <= io_A_Valid_7_delay_23_19;
    io_A_Valid_7_delay_25_17 <= io_A_Valid_7_delay_24_18;
    io_A_Valid_7_delay_26_16 <= io_A_Valid_7_delay_25_17;
    io_A_Valid_7_delay_27_15 <= io_A_Valid_7_delay_26_16;
    io_A_Valid_7_delay_28_14 <= io_A_Valid_7_delay_27_15;
    io_A_Valid_7_delay_29_13 <= io_A_Valid_7_delay_28_14;
    io_A_Valid_7_delay_30_12 <= io_A_Valid_7_delay_29_13;
    io_A_Valid_7_delay_31_11 <= io_A_Valid_7_delay_30_12;
    io_A_Valid_7_delay_32_10 <= io_A_Valid_7_delay_31_11;
    io_A_Valid_7_delay_33_9 <= io_A_Valid_7_delay_32_10;
    io_A_Valid_7_delay_34_8 <= io_A_Valid_7_delay_33_9;
    io_A_Valid_7_delay_35_7 <= io_A_Valid_7_delay_34_8;
    io_A_Valid_7_delay_36_6 <= io_A_Valid_7_delay_35_7;
    io_A_Valid_7_delay_37_5 <= io_A_Valid_7_delay_36_6;
    io_A_Valid_7_delay_38_4 <= io_A_Valid_7_delay_37_5;
    io_A_Valid_7_delay_39_3 <= io_A_Valid_7_delay_38_4;
    io_A_Valid_7_delay_40_2 <= io_A_Valid_7_delay_39_3;
    io_A_Valid_7_delay_41_1 <= io_A_Valid_7_delay_40_2;
    io_A_Valid_7_delay_42 <= io_A_Valid_7_delay_41_1;
    io_B_Valid_42_delay_1_6 <= io_B_Valid_42;
    io_B_Valid_42_delay_2_5 <= io_B_Valid_42_delay_1_6;
    io_B_Valid_42_delay_3_4 <= io_B_Valid_42_delay_2_5;
    io_B_Valid_42_delay_4_3 <= io_B_Valid_42_delay_3_4;
    io_B_Valid_42_delay_5_2 <= io_B_Valid_42_delay_4_3;
    io_B_Valid_42_delay_6_1 <= io_B_Valid_42_delay_5_2;
    io_B_Valid_42_delay_7 <= io_B_Valid_42_delay_6_1;
    io_A_Valid_7_delay_1_42 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_41 <= io_A_Valid_7_delay_1_42;
    io_A_Valid_7_delay_3_40 <= io_A_Valid_7_delay_2_41;
    io_A_Valid_7_delay_4_39 <= io_A_Valid_7_delay_3_40;
    io_A_Valid_7_delay_5_38 <= io_A_Valid_7_delay_4_39;
    io_A_Valid_7_delay_6_37 <= io_A_Valid_7_delay_5_38;
    io_A_Valid_7_delay_7_36 <= io_A_Valid_7_delay_6_37;
    io_A_Valid_7_delay_8_35 <= io_A_Valid_7_delay_7_36;
    io_A_Valid_7_delay_9_34 <= io_A_Valid_7_delay_8_35;
    io_A_Valid_7_delay_10_33 <= io_A_Valid_7_delay_9_34;
    io_A_Valid_7_delay_11_32 <= io_A_Valid_7_delay_10_33;
    io_A_Valid_7_delay_12_31 <= io_A_Valid_7_delay_11_32;
    io_A_Valid_7_delay_13_30 <= io_A_Valid_7_delay_12_31;
    io_A_Valid_7_delay_14_29 <= io_A_Valid_7_delay_13_30;
    io_A_Valid_7_delay_15_28 <= io_A_Valid_7_delay_14_29;
    io_A_Valid_7_delay_16_27 <= io_A_Valid_7_delay_15_28;
    io_A_Valid_7_delay_17_26 <= io_A_Valid_7_delay_16_27;
    io_A_Valid_7_delay_18_25 <= io_A_Valid_7_delay_17_26;
    io_A_Valid_7_delay_19_24 <= io_A_Valid_7_delay_18_25;
    io_A_Valid_7_delay_20_23 <= io_A_Valid_7_delay_19_24;
    io_A_Valid_7_delay_21_22 <= io_A_Valid_7_delay_20_23;
    io_A_Valid_7_delay_22_21 <= io_A_Valid_7_delay_21_22;
    io_A_Valid_7_delay_23_20 <= io_A_Valid_7_delay_22_21;
    io_A_Valid_7_delay_24_19 <= io_A_Valid_7_delay_23_20;
    io_A_Valid_7_delay_25_18 <= io_A_Valid_7_delay_24_19;
    io_A_Valid_7_delay_26_17 <= io_A_Valid_7_delay_25_18;
    io_A_Valid_7_delay_27_16 <= io_A_Valid_7_delay_26_17;
    io_A_Valid_7_delay_28_15 <= io_A_Valid_7_delay_27_16;
    io_A_Valid_7_delay_29_14 <= io_A_Valid_7_delay_28_15;
    io_A_Valid_7_delay_30_13 <= io_A_Valid_7_delay_29_14;
    io_A_Valid_7_delay_31_12 <= io_A_Valid_7_delay_30_13;
    io_A_Valid_7_delay_32_11 <= io_A_Valid_7_delay_31_12;
    io_A_Valid_7_delay_33_10 <= io_A_Valid_7_delay_32_11;
    io_A_Valid_7_delay_34_9 <= io_A_Valid_7_delay_33_10;
    io_A_Valid_7_delay_35_8 <= io_A_Valid_7_delay_34_9;
    io_A_Valid_7_delay_36_7 <= io_A_Valid_7_delay_35_8;
    io_A_Valid_7_delay_37_6 <= io_A_Valid_7_delay_36_7;
    io_A_Valid_7_delay_38_5 <= io_A_Valid_7_delay_37_6;
    io_A_Valid_7_delay_39_4 <= io_A_Valid_7_delay_38_5;
    io_A_Valid_7_delay_40_3 <= io_A_Valid_7_delay_39_4;
    io_A_Valid_7_delay_41_2 <= io_A_Valid_7_delay_40_3;
    io_A_Valid_7_delay_42_1 <= io_A_Valid_7_delay_41_2;
    io_A_Valid_7_delay_43 <= io_A_Valid_7_delay_42_1;
    io_B_Valid_43_delay_1_6 <= io_B_Valid_43;
    io_B_Valid_43_delay_2_5 <= io_B_Valid_43_delay_1_6;
    io_B_Valid_43_delay_3_4 <= io_B_Valid_43_delay_2_5;
    io_B_Valid_43_delay_4_3 <= io_B_Valid_43_delay_3_4;
    io_B_Valid_43_delay_5_2 <= io_B_Valid_43_delay_4_3;
    io_B_Valid_43_delay_6_1 <= io_B_Valid_43_delay_5_2;
    io_B_Valid_43_delay_7 <= io_B_Valid_43_delay_6_1;
    io_A_Valid_7_delay_1_43 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_42 <= io_A_Valid_7_delay_1_43;
    io_A_Valid_7_delay_3_41 <= io_A_Valid_7_delay_2_42;
    io_A_Valid_7_delay_4_40 <= io_A_Valid_7_delay_3_41;
    io_A_Valid_7_delay_5_39 <= io_A_Valid_7_delay_4_40;
    io_A_Valid_7_delay_6_38 <= io_A_Valid_7_delay_5_39;
    io_A_Valid_7_delay_7_37 <= io_A_Valid_7_delay_6_38;
    io_A_Valid_7_delay_8_36 <= io_A_Valid_7_delay_7_37;
    io_A_Valid_7_delay_9_35 <= io_A_Valid_7_delay_8_36;
    io_A_Valid_7_delay_10_34 <= io_A_Valid_7_delay_9_35;
    io_A_Valid_7_delay_11_33 <= io_A_Valid_7_delay_10_34;
    io_A_Valid_7_delay_12_32 <= io_A_Valid_7_delay_11_33;
    io_A_Valid_7_delay_13_31 <= io_A_Valid_7_delay_12_32;
    io_A_Valid_7_delay_14_30 <= io_A_Valid_7_delay_13_31;
    io_A_Valid_7_delay_15_29 <= io_A_Valid_7_delay_14_30;
    io_A_Valid_7_delay_16_28 <= io_A_Valid_7_delay_15_29;
    io_A_Valid_7_delay_17_27 <= io_A_Valid_7_delay_16_28;
    io_A_Valid_7_delay_18_26 <= io_A_Valid_7_delay_17_27;
    io_A_Valid_7_delay_19_25 <= io_A_Valid_7_delay_18_26;
    io_A_Valid_7_delay_20_24 <= io_A_Valid_7_delay_19_25;
    io_A_Valid_7_delay_21_23 <= io_A_Valid_7_delay_20_24;
    io_A_Valid_7_delay_22_22 <= io_A_Valid_7_delay_21_23;
    io_A_Valid_7_delay_23_21 <= io_A_Valid_7_delay_22_22;
    io_A_Valid_7_delay_24_20 <= io_A_Valid_7_delay_23_21;
    io_A_Valid_7_delay_25_19 <= io_A_Valid_7_delay_24_20;
    io_A_Valid_7_delay_26_18 <= io_A_Valid_7_delay_25_19;
    io_A_Valid_7_delay_27_17 <= io_A_Valid_7_delay_26_18;
    io_A_Valid_7_delay_28_16 <= io_A_Valid_7_delay_27_17;
    io_A_Valid_7_delay_29_15 <= io_A_Valid_7_delay_28_16;
    io_A_Valid_7_delay_30_14 <= io_A_Valid_7_delay_29_15;
    io_A_Valid_7_delay_31_13 <= io_A_Valid_7_delay_30_14;
    io_A_Valid_7_delay_32_12 <= io_A_Valid_7_delay_31_13;
    io_A_Valid_7_delay_33_11 <= io_A_Valid_7_delay_32_12;
    io_A_Valid_7_delay_34_10 <= io_A_Valid_7_delay_33_11;
    io_A_Valid_7_delay_35_9 <= io_A_Valid_7_delay_34_10;
    io_A_Valid_7_delay_36_8 <= io_A_Valid_7_delay_35_9;
    io_A_Valid_7_delay_37_7 <= io_A_Valid_7_delay_36_8;
    io_A_Valid_7_delay_38_6 <= io_A_Valid_7_delay_37_7;
    io_A_Valid_7_delay_39_5 <= io_A_Valid_7_delay_38_6;
    io_A_Valid_7_delay_40_4 <= io_A_Valid_7_delay_39_5;
    io_A_Valid_7_delay_41_3 <= io_A_Valid_7_delay_40_4;
    io_A_Valid_7_delay_42_2 <= io_A_Valid_7_delay_41_3;
    io_A_Valid_7_delay_43_1 <= io_A_Valid_7_delay_42_2;
    io_A_Valid_7_delay_44 <= io_A_Valid_7_delay_43_1;
    io_B_Valid_44_delay_1_6 <= io_B_Valid_44;
    io_B_Valid_44_delay_2_5 <= io_B_Valid_44_delay_1_6;
    io_B_Valid_44_delay_3_4 <= io_B_Valid_44_delay_2_5;
    io_B_Valid_44_delay_4_3 <= io_B_Valid_44_delay_3_4;
    io_B_Valid_44_delay_5_2 <= io_B_Valid_44_delay_4_3;
    io_B_Valid_44_delay_6_1 <= io_B_Valid_44_delay_5_2;
    io_B_Valid_44_delay_7 <= io_B_Valid_44_delay_6_1;
    io_A_Valid_7_delay_1_44 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_43 <= io_A_Valid_7_delay_1_44;
    io_A_Valid_7_delay_3_42 <= io_A_Valid_7_delay_2_43;
    io_A_Valid_7_delay_4_41 <= io_A_Valid_7_delay_3_42;
    io_A_Valid_7_delay_5_40 <= io_A_Valid_7_delay_4_41;
    io_A_Valid_7_delay_6_39 <= io_A_Valid_7_delay_5_40;
    io_A_Valid_7_delay_7_38 <= io_A_Valid_7_delay_6_39;
    io_A_Valid_7_delay_8_37 <= io_A_Valid_7_delay_7_38;
    io_A_Valid_7_delay_9_36 <= io_A_Valid_7_delay_8_37;
    io_A_Valid_7_delay_10_35 <= io_A_Valid_7_delay_9_36;
    io_A_Valid_7_delay_11_34 <= io_A_Valid_7_delay_10_35;
    io_A_Valid_7_delay_12_33 <= io_A_Valid_7_delay_11_34;
    io_A_Valid_7_delay_13_32 <= io_A_Valid_7_delay_12_33;
    io_A_Valid_7_delay_14_31 <= io_A_Valid_7_delay_13_32;
    io_A_Valid_7_delay_15_30 <= io_A_Valid_7_delay_14_31;
    io_A_Valid_7_delay_16_29 <= io_A_Valid_7_delay_15_30;
    io_A_Valid_7_delay_17_28 <= io_A_Valid_7_delay_16_29;
    io_A_Valid_7_delay_18_27 <= io_A_Valid_7_delay_17_28;
    io_A_Valid_7_delay_19_26 <= io_A_Valid_7_delay_18_27;
    io_A_Valid_7_delay_20_25 <= io_A_Valid_7_delay_19_26;
    io_A_Valid_7_delay_21_24 <= io_A_Valid_7_delay_20_25;
    io_A_Valid_7_delay_22_23 <= io_A_Valid_7_delay_21_24;
    io_A_Valid_7_delay_23_22 <= io_A_Valid_7_delay_22_23;
    io_A_Valid_7_delay_24_21 <= io_A_Valid_7_delay_23_22;
    io_A_Valid_7_delay_25_20 <= io_A_Valid_7_delay_24_21;
    io_A_Valid_7_delay_26_19 <= io_A_Valid_7_delay_25_20;
    io_A_Valid_7_delay_27_18 <= io_A_Valid_7_delay_26_19;
    io_A_Valid_7_delay_28_17 <= io_A_Valid_7_delay_27_18;
    io_A_Valid_7_delay_29_16 <= io_A_Valid_7_delay_28_17;
    io_A_Valid_7_delay_30_15 <= io_A_Valid_7_delay_29_16;
    io_A_Valid_7_delay_31_14 <= io_A_Valid_7_delay_30_15;
    io_A_Valid_7_delay_32_13 <= io_A_Valid_7_delay_31_14;
    io_A_Valid_7_delay_33_12 <= io_A_Valid_7_delay_32_13;
    io_A_Valid_7_delay_34_11 <= io_A_Valid_7_delay_33_12;
    io_A_Valid_7_delay_35_10 <= io_A_Valid_7_delay_34_11;
    io_A_Valid_7_delay_36_9 <= io_A_Valid_7_delay_35_10;
    io_A_Valid_7_delay_37_8 <= io_A_Valid_7_delay_36_9;
    io_A_Valid_7_delay_38_7 <= io_A_Valid_7_delay_37_8;
    io_A_Valid_7_delay_39_6 <= io_A_Valid_7_delay_38_7;
    io_A_Valid_7_delay_40_5 <= io_A_Valid_7_delay_39_6;
    io_A_Valid_7_delay_41_4 <= io_A_Valid_7_delay_40_5;
    io_A_Valid_7_delay_42_3 <= io_A_Valid_7_delay_41_4;
    io_A_Valid_7_delay_43_2 <= io_A_Valid_7_delay_42_3;
    io_A_Valid_7_delay_44_1 <= io_A_Valid_7_delay_43_2;
    io_A_Valid_7_delay_45 <= io_A_Valid_7_delay_44_1;
    io_B_Valid_45_delay_1_6 <= io_B_Valid_45;
    io_B_Valid_45_delay_2_5 <= io_B_Valid_45_delay_1_6;
    io_B_Valid_45_delay_3_4 <= io_B_Valid_45_delay_2_5;
    io_B_Valid_45_delay_4_3 <= io_B_Valid_45_delay_3_4;
    io_B_Valid_45_delay_5_2 <= io_B_Valid_45_delay_4_3;
    io_B_Valid_45_delay_6_1 <= io_B_Valid_45_delay_5_2;
    io_B_Valid_45_delay_7 <= io_B_Valid_45_delay_6_1;
    io_A_Valid_7_delay_1_45 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_44 <= io_A_Valid_7_delay_1_45;
    io_A_Valid_7_delay_3_43 <= io_A_Valid_7_delay_2_44;
    io_A_Valid_7_delay_4_42 <= io_A_Valid_7_delay_3_43;
    io_A_Valid_7_delay_5_41 <= io_A_Valid_7_delay_4_42;
    io_A_Valid_7_delay_6_40 <= io_A_Valid_7_delay_5_41;
    io_A_Valid_7_delay_7_39 <= io_A_Valid_7_delay_6_40;
    io_A_Valid_7_delay_8_38 <= io_A_Valid_7_delay_7_39;
    io_A_Valid_7_delay_9_37 <= io_A_Valid_7_delay_8_38;
    io_A_Valid_7_delay_10_36 <= io_A_Valid_7_delay_9_37;
    io_A_Valid_7_delay_11_35 <= io_A_Valid_7_delay_10_36;
    io_A_Valid_7_delay_12_34 <= io_A_Valid_7_delay_11_35;
    io_A_Valid_7_delay_13_33 <= io_A_Valid_7_delay_12_34;
    io_A_Valid_7_delay_14_32 <= io_A_Valid_7_delay_13_33;
    io_A_Valid_7_delay_15_31 <= io_A_Valid_7_delay_14_32;
    io_A_Valid_7_delay_16_30 <= io_A_Valid_7_delay_15_31;
    io_A_Valid_7_delay_17_29 <= io_A_Valid_7_delay_16_30;
    io_A_Valid_7_delay_18_28 <= io_A_Valid_7_delay_17_29;
    io_A_Valid_7_delay_19_27 <= io_A_Valid_7_delay_18_28;
    io_A_Valid_7_delay_20_26 <= io_A_Valid_7_delay_19_27;
    io_A_Valid_7_delay_21_25 <= io_A_Valid_7_delay_20_26;
    io_A_Valid_7_delay_22_24 <= io_A_Valid_7_delay_21_25;
    io_A_Valid_7_delay_23_23 <= io_A_Valid_7_delay_22_24;
    io_A_Valid_7_delay_24_22 <= io_A_Valid_7_delay_23_23;
    io_A_Valid_7_delay_25_21 <= io_A_Valid_7_delay_24_22;
    io_A_Valid_7_delay_26_20 <= io_A_Valid_7_delay_25_21;
    io_A_Valid_7_delay_27_19 <= io_A_Valid_7_delay_26_20;
    io_A_Valid_7_delay_28_18 <= io_A_Valid_7_delay_27_19;
    io_A_Valid_7_delay_29_17 <= io_A_Valid_7_delay_28_18;
    io_A_Valid_7_delay_30_16 <= io_A_Valid_7_delay_29_17;
    io_A_Valid_7_delay_31_15 <= io_A_Valid_7_delay_30_16;
    io_A_Valid_7_delay_32_14 <= io_A_Valid_7_delay_31_15;
    io_A_Valid_7_delay_33_13 <= io_A_Valid_7_delay_32_14;
    io_A_Valid_7_delay_34_12 <= io_A_Valid_7_delay_33_13;
    io_A_Valid_7_delay_35_11 <= io_A_Valid_7_delay_34_12;
    io_A_Valid_7_delay_36_10 <= io_A_Valid_7_delay_35_11;
    io_A_Valid_7_delay_37_9 <= io_A_Valid_7_delay_36_10;
    io_A_Valid_7_delay_38_8 <= io_A_Valid_7_delay_37_9;
    io_A_Valid_7_delay_39_7 <= io_A_Valid_7_delay_38_8;
    io_A_Valid_7_delay_40_6 <= io_A_Valid_7_delay_39_7;
    io_A_Valid_7_delay_41_5 <= io_A_Valid_7_delay_40_6;
    io_A_Valid_7_delay_42_4 <= io_A_Valid_7_delay_41_5;
    io_A_Valid_7_delay_43_3 <= io_A_Valid_7_delay_42_4;
    io_A_Valid_7_delay_44_2 <= io_A_Valid_7_delay_43_3;
    io_A_Valid_7_delay_45_1 <= io_A_Valid_7_delay_44_2;
    io_A_Valid_7_delay_46 <= io_A_Valid_7_delay_45_1;
    io_B_Valid_46_delay_1_6 <= io_B_Valid_46;
    io_B_Valid_46_delay_2_5 <= io_B_Valid_46_delay_1_6;
    io_B_Valid_46_delay_3_4 <= io_B_Valid_46_delay_2_5;
    io_B_Valid_46_delay_4_3 <= io_B_Valid_46_delay_3_4;
    io_B_Valid_46_delay_5_2 <= io_B_Valid_46_delay_4_3;
    io_B_Valid_46_delay_6_1 <= io_B_Valid_46_delay_5_2;
    io_B_Valid_46_delay_7 <= io_B_Valid_46_delay_6_1;
    io_A_Valid_7_delay_1_46 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_45 <= io_A_Valid_7_delay_1_46;
    io_A_Valid_7_delay_3_44 <= io_A_Valid_7_delay_2_45;
    io_A_Valid_7_delay_4_43 <= io_A_Valid_7_delay_3_44;
    io_A_Valid_7_delay_5_42 <= io_A_Valid_7_delay_4_43;
    io_A_Valid_7_delay_6_41 <= io_A_Valid_7_delay_5_42;
    io_A_Valid_7_delay_7_40 <= io_A_Valid_7_delay_6_41;
    io_A_Valid_7_delay_8_39 <= io_A_Valid_7_delay_7_40;
    io_A_Valid_7_delay_9_38 <= io_A_Valid_7_delay_8_39;
    io_A_Valid_7_delay_10_37 <= io_A_Valid_7_delay_9_38;
    io_A_Valid_7_delay_11_36 <= io_A_Valid_7_delay_10_37;
    io_A_Valid_7_delay_12_35 <= io_A_Valid_7_delay_11_36;
    io_A_Valid_7_delay_13_34 <= io_A_Valid_7_delay_12_35;
    io_A_Valid_7_delay_14_33 <= io_A_Valid_7_delay_13_34;
    io_A_Valid_7_delay_15_32 <= io_A_Valid_7_delay_14_33;
    io_A_Valid_7_delay_16_31 <= io_A_Valid_7_delay_15_32;
    io_A_Valid_7_delay_17_30 <= io_A_Valid_7_delay_16_31;
    io_A_Valid_7_delay_18_29 <= io_A_Valid_7_delay_17_30;
    io_A_Valid_7_delay_19_28 <= io_A_Valid_7_delay_18_29;
    io_A_Valid_7_delay_20_27 <= io_A_Valid_7_delay_19_28;
    io_A_Valid_7_delay_21_26 <= io_A_Valid_7_delay_20_27;
    io_A_Valid_7_delay_22_25 <= io_A_Valid_7_delay_21_26;
    io_A_Valid_7_delay_23_24 <= io_A_Valid_7_delay_22_25;
    io_A_Valid_7_delay_24_23 <= io_A_Valid_7_delay_23_24;
    io_A_Valid_7_delay_25_22 <= io_A_Valid_7_delay_24_23;
    io_A_Valid_7_delay_26_21 <= io_A_Valid_7_delay_25_22;
    io_A_Valid_7_delay_27_20 <= io_A_Valid_7_delay_26_21;
    io_A_Valid_7_delay_28_19 <= io_A_Valid_7_delay_27_20;
    io_A_Valid_7_delay_29_18 <= io_A_Valid_7_delay_28_19;
    io_A_Valid_7_delay_30_17 <= io_A_Valid_7_delay_29_18;
    io_A_Valid_7_delay_31_16 <= io_A_Valid_7_delay_30_17;
    io_A_Valid_7_delay_32_15 <= io_A_Valid_7_delay_31_16;
    io_A_Valid_7_delay_33_14 <= io_A_Valid_7_delay_32_15;
    io_A_Valid_7_delay_34_13 <= io_A_Valid_7_delay_33_14;
    io_A_Valid_7_delay_35_12 <= io_A_Valid_7_delay_34_13;
    io_A_Valid_7_delay_36_11 <= io_A_Valid_7_delay_35_12;
    io_A_Valid_7_delay_37_10 <= io_A_Valid_7_delay_36_11;
    io_A_Valid_7_delay_38_9 <= io_A_Valid_7_delay_37_10;
    io_A_Valid_7_delay_39_8 <= io_A_Valid_7_delay_38_9;
    io_A_Valid_7_delay_40_7 <= io_A_Valid_7_delay_39_8;
    io_A_Valid_7_delay_41_6 <= io_A_Valid_7_delay_40_7;
    io_A_Valid_7_delay_42_5 <= io_A_Valid_7_delay_41_6;
    io_A_Valid_7_delay_43_4 <= io_A_Valid_7_delay_42_5;
    io_A_Valid_7_delay_44_3 <= io_A_Valid_7_delay_43_4;
    io_A_Valid_7_delay_45_2 <= io_A_Valid_7_delay_44_3;
    io_A_Valid_7_delay_46_1 <= io_A_Valid_7_delay_45_2;
    io_A_Valid_7_delay_47 <= io_A_Valid_7_delay_46_1;
    io_B_Valid_47_delay_1_6 <= io_B_Valid_47;
    io_B_Valid_47_delay_2_5 <= io_B_Valid_47_delay_1_6;
    io_B_Valid_47_delay_3_4 <= io_B_Valid_47_delay_2_5;
    io_B_Valid_47_delay_4_3 <= io_B_Valid_47_delay_3_4;
    io_B_Valid_47_delay_5_2 <= io_B_Valid_47_delay_4_3;
    io_B_Valid_47_delay_6_1 <= io_B_Valid_47_delay_5_2;
    io_B_Valid_47_delay_7 <= io_B_Valid_47_delay_6_1;
    io_A_Valid_7_delay_1_47 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_46 <= io_A_Valid_7_delay_1_47;
    io_A_Valid_7_delay_3_45 <= io_A_Valid_7_delay_2_46;
    io_A_Valid_7_delay_4_44 <= io_A_Valid_7_delay_3_45;
    io_A_Valid_7_delay_5_43 <= io_A_Valid_7_delay_4_44;
    io_A_Valid_7_delay_6_42 <= io_A_Valid_7_delay_5_43;
    io_A_Valid_7_delay_7_41 <= io_A_Valid_7_delay_6_42;
    io_A_Valid_7_delay_8_40 <= io_A_Valid_7_delay_7_41;
    io_A_Valid_7_delay_9_39 <= io_A_Valid_7_delay_8_40;
    io_A_Valid_7_delay_10_38 <= io_A_Valid_7_delay_9_39;
    io_A_Valid_7_delay_11_37 <= io_A_Valid_7_delay_10_38;
    io_A_Valid_7_delay_12_36 <= io_A_Valid_7_delay_11_37;
    io_A_Valid_7_delay_13_35 <= io_A_Valid_7_delay_12_36;
    io_A_Valid_7_delay_14_34 <= io_A_Valid_7_delay_13_35;
    io_A_Valid_7_delay_15_33 <= io_A_Valid_7_delay_14_34;
    io_A_Valid_7_delay_16_32 <= io_A_Valid_7_delay_15_33;
    io_A_Valid_7_delay_17_31 <= io_A_Valid_7_delay_16_32;
    io_A_Valid_7_delay_18_30 <= io_A_Valid_7_delay_17_31;
    io_A_Valid_7_delay_19_29 <= io_A_Valid_7_delay_18_30;
    io_A_Valid_7_delay_20_28 <= io_A_Valid_7_delay_19_29;
    io_A_Valid_7_delay_21_27 <= io_A_Valid_7_delay_20_28;
    io_A_Valid_7_delay_22_26 <= io_A_Valid_7_delay_21_27;
    io_A_Valid_7_delay_23_25 <= io_A_Valid_7_delay_22_26;
    io_A_Valid_7_delay_24_24 <= io_A_Valid_7_delay_23_25;
    io_A_Valid_7_delay_25_23 <= io_A_Valid_7_delay_24_24;
    io_A_Valid_7_delay_26_22 <= io_A_Valid_7_delay_25_23;
    io_A_Valid_7_delay_27_21 <= io_A_Valid_7_delay_26_22;
    io_A_Valid_7_delay_28_20 <= io_A_Valid_7_delay_27_21;
    io_A_Valid_7_delay_29_19 <= io_A_Valid_7_delay_28_20;
    io_A_Valid_7_delay_30_18 <= io_A_Valid_7_delay_29_19;
    io_A_Valid_7_delay_31_17 <= io_A_Valid_7_delay_30_18;
    io_A_Valid_7_delay_32_16 <= io_A_Valid_7_delay_31_17;
    io_A_Valid_7_delay_33_15 <= io_A_Valid_7_delay_32_16;
    io_A_Valid_7_delay_34_14 <= io_A_Valid_7_delay_33_15;
    io_A_Valid_7_delay_35_13 <= io_A_Valid_7_delay_34_14;
    io_A_Valid_7_delay_36_12 <= io_A_Valid_7_delay_35_13;
    io_A_Valid_7_delay_37_11 <= io_A_Valid_7_delay_36_12;
    io_A_Valid_7_delay_38_10 <= io_A_Valid_7_delay_37_11;
    io_A_Valid_7_delay_39_9 <= io_A_Valid_7_delay_38_10;
    io_A_Valid_7_delay_40_8 <= io_A_Valid_7_delay_39_9;
    io_A_Valid_7_delay_41_7 <= io_A_Valid_7_delay_40_8;
    io_A_Valid_7_delay_42_6 <= io_A_Valid_7_delay_41_7;
    io_A_Valid_7_delay_43_5 <= io_A_Valid_7_delay_42_6;
    io_A_Valid_7_delay_44_4 <= io_A_Valid_7_delay_43_5;
    io_A_Valid_7_delay_45_3 <= io_A_Valid_7_delay_44_4;
    io_A_Valid_7_delay_46_2 <= io_A_Valid_7_delay_45_3;
    io_A_Valid_7_delay_47_1 <= io_A_Valid_7_delay_46_2;
    io_A_Valid_7_delay_48 <= io_A_Valid_7_delay_47_1;
    io_B_Valid_48_delay_1_6 <= io_B_Valid_48;
    io_B_Valid_48_delay_2_5 <= io_B_Valid_48_delay_1_6;
    io_B_Valid_48_delay_3_4 <= io_B_Valid_48_delay_2_5;
    io_B_Valid_48_delay_4_3 <= io_B_Valid_48_delay_3_4;
    io_B_Valid_48_delay_5_2 <= io_B_Valid_48_delay_4_3;
    io_B_Valid_48_delay_6_1 <= io_B_Valid_48_delay_5_2;
    io_B_Valid_48_delay_7 <= io_B_Valid_48_delay_6_1;
    io_A_Valid_7_delay_1_48 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_47 <= io_A_Valid_7_delay_1_48;
    io_A_Valid_7_delay_3_46 <= io_A_Valid_7_delay_2_47;
    io_A_Valid_7_delay_4_45 <= io_A_Valid_7_delay_3_46;
    io_A_Valid_7_delay_5_44 <= io_A_Valid_7_delay_4_45;
    io_A_Valid_7_delay_6_43 <= io_A_Valid_7_delay_5_44;
    io_A_Valid_7_delay_7_42 <= io_A_Valid_7_delay_6_43;
    io_A_Valid_7_delay_8_41 <= io_A_Valid_7_delay_7_42;
    io_A_Valid_7_delay_9_40 <= io_A_Valid_7_delay_8_41;
    io_A_Valid_7_delay_10_39 <= io_A_Valid_7_delay_9_40;
    io_A_Valid_7_delay_11_38 <= io_A_Valid_7_delay_10_39;
    io_A_Valid_7_delay_12_37 <= io_A_Valid_7_delay_11_38;
    io_A_Valid_7_delay_13_36 <= io_A_Valid_7_delay_12_37;
    io_A_Valid_7_delay_14_35 <= io_A_Valid_7_delay_13_36;
    io_A_Valid_7_delay_15_34 <= io_A_Valid_7_delay_14_35;
    io_A_Valid_7_delay_16_33 <= io_A_Valid_7_delay_15_34;
    io_A_Valid_7_delay_17_32 <= io_A_Valid_7_delay_16_33;
    io_A_Valid_7_delay_18_31 <= io_A_Valid_7_delay_17_32;
    io_A_Valid_7_delay_19_30 <= io_A_Valid_7_delay_18_31;
    io_A_Valid_7_delay_20_29 <= io_A_Valid_7_delay_19_30;
    io_A_Valid_7_delay_21_28 <= io_A_Valid_7_delay_20_29;
    io_A_Valid_7_delay_22_27 <= io_A_Valid_7_delay_21_28;
    io_A_Valid_7_delay_23_26 <= io_A_Valid_7_delay_22_27;
    io_A_Valid_7_delay_24_25 <= io_A_Valid_7_delay_23_26;
    io_A_Valid_7_delay_25_24 <= io_A_Valid_7_delay_24_25;
    io_A_Valid_7_delay_26_23 <= io_A_Valid_7_delay_25_24;
    io_A_Valid_7_delay_27_22 <= io_A_Valid_7_delay_26_23;
    io_A_Valid_7_delay_28_21 <= io_A_Valid_7_delay_27_22;
    io_A_Valid_7_delay_29_20 <= io_A_Valid_7_delay_28_21;
    io_A_Valid_7_delay_30_19 <= io_A_Valid_7_delay_29_20;
    io_A_Valid_7_delay_31_18 <= io_A_Valid_7_delay_30_19;
    io_A_Valid_7_delay_32_17 <= io_A_Valid_7_delay_31_18;
    io_A_Valid_7_delay_33_16 <= io_A_Valid_7_delay_32_17;
    io_A_Valid_7_delay_34_15 <= io_A_Valid_7_delay_33_16;
    io_A_Valid_7_delay_35_14 <= io_A_Valid_7_delay_34_15;
    io_A_Valid_7_delay_36_13 <= io_A_Valid_7_delay_35_14;
    io_A_Valid_7_delay_37_12 <= io_A_Valid_7_delay_36_13;
    io_A_Valid_7_delay_38_11 <= io_A_Valid_7_delay_37_12;
    io_A_Valid_7_delay_39_10 <= io_A_Valid_7_delay_38_11;
    io_A_Valid_7_delay_40_9 <= io_A_Valid_7_delay_39_10;
    io_A_Valid_7_delay_41_8 <= io_A_Valid_7_delay_40_9;
    io_A_Valid_7_delay_42_7 <= io_A_Valid_7_delay_41_8;
    io_A_Valid_7_delay_43_6 <= io_A_Valid_7_delay_42_7;
    io_A_Valid_7_delay_44_5 <= io_A_Valid_7_delay_43_6;
    io_A_Valid_7_delay_45_4 <= io_A_Valid_7_delay_44_5;
    io_A_Valid_7_delay_46_3 <= io_A_Valid_7_delay_45_4;
    io_A_Valid_7_delay_47_2 <= io_A_Valid_7_delay_46_3;
    io_A_Valid_7_delay_48_1 <= io_A_Valid_7_delay_47_2;
    io_A_Valid_7_delay_49 <= io_A_Valid_7_delay_48_1;
    io_B_Valid_49_delay_1_6 <= io_B_Valid_49;
    io_B_Valid_49_delay_2_5 <= io_B_Valid_49_delay_1_6;
    io_B_Valid_49_delay_3_4 <= io_B_Valid_49_delay_2_5;
    io_B_Valid_49_delay_4_3 <= io_B_Valid_49_delay_3_4;
    io_B_Valid_49_delay_5_2 <= io_B_Valid_49_delay_4_3;
    io_B_Valid_49_delay_6_1 <= io_B_Valid_49_delay_5_2;
    io_B_Valid_49_delay_7 <= io_B_Valid_49_delay_6_1;
    io_A_Valid_7_delay_1_49 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_48 <= io_A_Valid_7_delay_1_49;
    io_A_Valid_7_delay_3_47 <= io_A_Valid_7_delay_2_48;
    io_A_Valid_7_delay_4_46 <= io_A_Valid_7_delay_3_47;
    io_A_Valid_7_delay_5_45 <= io_A_Valid_7_delay_4_46;
    io_A_Valid_7_delay_6_44 <= io_A_Valid_7_delay_5_45;
    io_A_Valid_7_delay_7_43 <= io_A_Valid_7_delay_6_44;
    io_A_Valid_7_delay_8_42 <= io_A_Valid_7_delay_7_43;
    io_A_Valid_7_delay_9_41 <= io_A_Valid_7_delay_8_42;
    io_A_Valid_7_delay_10_40 <= io_A_Valid_7_delay_9_41;
    io_A_Valid_7_delay_11_39 <= io_A_Valid_7_delay_10_40;
    io_A_Valid_7_delay_12_38 <= io_A_Valid_7_delay_11_39;
    io_A_Valid_7_delay_13_37 <= io_A_Valid_7_delay_12_38;
    io_A_Valid_7_delay_14_36 <= io_A_Valid_7_delay_13_37;
    io_A_Valid_7_delay_15_35 <= io_A_Valid_7_delay_14_36;
    io_A_Valid_7_delay_16_34 <= io_A_Valid_7_delay_15_35;
    io_A_Valid_7_delay_17_33 <= io_A_Valid_7_delay_16_34;
    io_A_Valid_7_delay_18_32 <= io_A_Valid_7_delay_17_33;
    io_A_Valid_7_delay_19_31 <= io_A_Valid_7_delay_18_32;
    io_A_Valid_7_delay_20_30 <= io_A_Valid_7_delay_19_31;
    io_A_Valid_7_delay_21_29 <= io_A_Valid_7_delay_20_30;
    io_A_Valid_7_delay_22_28 <= io_A_Valid_7_delay_21_29;
    io_A_Valid_7_delay_23_27 <= io_A_Valid_7_delay_22_28;
    io_A_Valid_7_delay_24_26 <= io_A_Valid_7_delay_23_27;
    io_A_Valid_7_delay_25_25 <= io_A_Valid_7_delay_24_26;
    io_A_Valid_7_delay_26_24 <= io_A_Valid_7_delay_25_25;
    io_A_Valid_7_delay_27_23 <= io_A_Valid_7_delay_26_24;
    io_A_Valid_7_delay_28_22 <= io_A_Valid_7_delay_27_23;
    io_A_Valid_7_delay_29_21 <= io_A_Valid_7_delay_28_22;
    io_A_Valid_7_delay_30_20 <= io_A_Valid_7_delay_29_21;
    io_A_Valid_7_delay_31_19 <= io_A_Valid_7_delay_30_20;
    io_A_Valid_7_delay_32_18 <= io_A_Valid_7_delay_31_19;
    io_A_Valid_7_delay_33_17 <= io_A_Valid_7_delay_32_18;
    io_A_Valid_7_delay_34_16 <= io_A_Valid_7_delay_33_17;
    io_A_Valid_7_delay_35_15 <= io_A_Valid_7_delay_34_16;
    io_A_Valid_7_delay_36_14 <= io_A_Valid_7_delay_35_15;
    io_A_Valid_7_delay_37_13 <= io_A_Valid_7_delay_36_14;
    io_A_Valid_7_delay_38_12 <= io_A_Valid_7_delay_37_13;
    io_A_Valid_7_delay_39_11 <= io_A_Valid_7_delay_38_12;
    io_A_Valid_7_delay_40_10 <= io_A_Valid_7_delay_39_11;
    io_A_Valid_7_delay_41_9 <= io_A_Valid_7_delay_40_10;
    io_A_Valid_7_delay_42_8 <= io_A_Valid_7_delay_41_9;
    io_A_Valid_7_delay_43_7 <= io_A_Valid_7_delay_42_8;
    io_A_Valid_7_delay_44_6 <= io_A_Valid_7_delay_43_7;
    io_A_Valid_7_delay_45_5 <= io_A_Valid_7_delay_44_6;
    io_A_Valid_7_delay_46_4 <= io_A_Valid_7_delay_45_5;
    io_A_Valid_7_delay_47_3 <= io_A_Valid_7_delay_46_4;
    io_A_Valid_7_delay_48_2 <= io_A_Valid_7_delay_47_3;
    io_A_Valid_7_delay_49_1 <= io_A_Valid_7_delay_48_2;
    io_A_Valid_7_delay_50 <= io_A_Valid_7_delay_49_1;
    io_B_Valid_50_delay_1_6 <= io_B_Valid_50;
    io_B_Valid_50_delay_2_5 <= io_B_Valid_50_delay_1_6;
    io_B_Valid_50_delay_3_4 <= io_B_Valid_50_delay_2_5;
    io_B_Valid_50_delay_4_3 <= io_B_Valid_50_delay_3_4;
    io_B_Valid_50_delay_5_2 <= io_B_Valid_50_delay_4_3;
    io_B_Valid_50_delay_6_1 <= io_B_Valid_50_delay_5_2;
    io_B_Valid_50_delay_7 <= io_B_Valid_50_delay_6_1;
    io_A_Valid_7_delay_1_50 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_49 <= io_A_Valid_7_delay_1_50;
    io_A_Valid_7_delay_3_48 <= io_A_Valid_7_delay_2_49;
    io_A_Valid_7_delay_4_47 <= io_A_Valid_7_delay_3_48;
    io_A_Valid_7_delay_5_46 <= io_A_Valid_7_delay_4_47;
    io_A_Valid_7_delay_6_45 <= io_A_Valid_7_delay_5_46;
    io_A_Valid_7_delay_7_44 <= io_A_Valid_7_delay_6_45;
    io_A_Valid_7_delay_8_43 <= io_A_Valid_7_delay_7_44;
    io_A_Valid_7_delay_9_42 <= io_A_Valid_7_delay_8_43;
    io_A_Valid_7_delay_10_41 <= io_A_Valid_7_delay_9_42;
    io_A_Valid_7_delay_11_40 <= io_A_Valid_7_delay_10_41;
    io_A_Valid_7_delay_12_39 <= io_A_Valid_7_delay_11_40;
    io_A_Valid_7_delay_13_38 <= io_A_Valid_7_delay_12_39;
    io_A_Valid_7_delay_14_37 <= io_A_Valid_7_delay_13_38;
    io_A_Valid_7_delay_15_36 <= io_A_Valid_7_delay_14_37;
    io_A_Valid_7_delay_16_35 <= io_A_Valid_7_delay_15_36;
    io_A_Valid_7_delay_17_34 <= io_A_Valid_7_delay_16_35;
    io_A_Valid_7_delay_18_33 <= io_A_Valid_7_delay_17_34;
    io_A_Valid_7_delay_19_32 <= io_A_Valid_7_delay_18_33;
    io_A_Valid_7_delay_20_31 <= io_A_Valid_7_delay_19_32;
    io_A_Valid_7_delay_21_30 <= io_A_Valid_7_delay_20_31;
    io_A_Valid_7_delay_22_29 <= io_A_Valid_7_delay_21_30;
    io_A_Valid_7_delay_23_28 <= io_A_Valid_7_delay_22_29;
    io_A_Valid_7_delay_24_27 <= io_A_Valid_7_delay_23_28;
    io_A_Valid_7_delay_25_26 <= io_A_Valid_7_delay_24_27;
    io_A_Valid_7_delay_26_25 <= io_A_Valid_7_delay_25_26;
    io_A_Valid_7_delay_27_24 <= io_A_Valid_7_delay_26_25;
    io_A_Valid_7_delay_28_23 <= io_A_Valid_7_delay_27_24;
    io_A_Valid_7_delay_29_22 <= io_A_Valid_7_delay_28_23;
    io_A_Valid_7_delay_30_21 <= io_A_Valid_7_delay_29_22;
    io_A_Valid_7_delay_31_20 <= io_A_Valid_7_delay_30_21;
    io_A_Valid_7_delay_32_19 <= io_A_Valid_7_delay_31_20;
    io_A_Valid_7_delay_33_18 <= io_A_Valid_7_delay_32_19;
    io_A_Valid_7_delay_34_17 <= io_A_Valid_7_delay_33_18;
    io_A_Valid_7_delay_35_16 <= io_A_Valid_7_delay_34_17;
    io_A_Valid_7_delay_36_15 <= io_A_Valid_7_delay_35_16;
    io_A_Valid_7_delay_37_14 <= io_A_Valid_7_delay_36_15;
    io_A_Valid_7_delay_38_13 <= io_A_Valid_7_delay_37_14;
    io_A_Valid_7_delay_39_12 <= io_A_Valid_7_delay_38_13;
    io_A_Valid_7_delay_40_11 <= io_A_Valid_7_delay_39_12;
    io_A_Valid_7_delay_41_10 <= io_A_Valid_7_delay_40_11;
    io_A_Valid_7_delay_42_9 <= io_A_Valid_7_delay_41_10;
    io_A_Valid_7_delay_43_8 <= io_A_Valid_7_delay_42_9;
    io_A_Valid_7_delay_44_7 <= io_A_Valid_7_delay_43_8;
    io_A_Valid_7_delay_45_6 <= io_A_Valid_7_delay_44_7;
    io_A_Valid_7_delay_46_5 <= io_A_Valid_7_delay_45_6;
    io_A_Valid_7_delay_47_4 <= io_A_Valid_7_delay_46_5;
    io_A_Valid_7_delay_48_3 <= io_A_Valid_7_delay_47_4;
    io_A_Valid_7_delay_49_2 <= io_A_Valid_7_delay_48_3;
    io_A_Valid_7_delay_50_1 <= io_A_Valid_7_delay_49_2;
    io_A_Valid_7_delay_51 <= io_A_Valid_7_delay_50_1;
    io_B_Valid_51_delay_1_6 <= io_B_Valid_51;
    io_B_Valid_51_delay_2_5 <= io_B_Valid_51_delay_1_6;
    io_B_Valid_51_delay_3_4 <= io_B_Valid_51_delay_2_5;
    io_B_Valid_51_delay_4_3 <= io_B_Valid_51_delay_3_4;
    io_B_Valid_51_delay_5_2 <= io_B_Valid_51_delay_4_3;
    io_B_Valid_51_delay_6_1 <= io_B_Valid_51_delay_5_2;
    io_B_Valid_51_delay_7 <= io_B_Valid_51_delay_6_1;
    io_A_Valid_7_delay_1_51 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_50 <= io_A_Valid_7_delay_1_51;
    io_A_Valid_7_delay_3_49 <= io_A_Valid_7_delay_2_50;
    io_A_Valid_7_delay_4_48 <= io_A_Valid_7_delay_3_49;
    io_A_Valid_7_delay_5_47 <= io_A_Valid_7_delay_4_48;
    io_A_Valid_7_delay_6_46 <= io_A_Valid_7_delay_5_47;
    io_A_Valid_7_delay_7_45 <= io_A_Valid_7_delay_6_46;
    io_A_Valid_7_delay_8_44 <= io_A_Valid_7_delay_7_45;
    io_A_Valid_7_delay_9_43 <= io_A_Valid_7_delay_8_44;
    io_A_Valid_7_delay_10_42 <= io_A_Valid_7_delay_9_43;
    io_A_Valid_7_delay_11_41 <= io_A_Valid_7_delay_10_42;
    io_A_Valid_7_delay_12_40 <= io_A_Valid_7_delay_11_41;
    io_A_Valid_7_delay_13_39 <= io_A_Valid_7_delay_12_40;
    io_A_Valid_7_delay_14_38 <= io_A_Valid_7_delay_13_39;
    io_A_Valid_7_delay_15_37 <= io_A_Valid_7_delay_14_38;
    io_A_Valid_7_delay_16_36 <= io_A_Valid_7_delay_15_37;
    io_A_Valid_7_delay_17_35 <= io_A_Valid_7_delay_16_36;
    io_A_Valid_7_delay_18_34 <= io_A_Valid_7_delay_17_35;
    io_A_Valid_7_delay_19_33 <= io_A_Valid_7_delay_18_34;
    io_A_Valid_7_delay_20_32 <= io_A_Valid_7_delay_19_33;
    io_A_Valid_7_delay_21_31 <= io_A_Valid_7_delay_20_32;
    io_A_Valid_7_delay_22_30 <= io_A_Valid_7_delay_21_31;
    io_A_Valid_7_delay_23_29 <= io_A_Valid_7_delay_22_30;
    io_A_Valid_7_delay_24_28 <= io_A_Valid_7_delay_23_29;
    io_A_Valid_7_delay_25_27 <= io_A_Valid_7_delay_24_28;
    io_A_Valid_7_delay_26_26 <= io_A_Valid_7_delay_25_27;
    io_A_Valid_7_delay_27_25 <= io_A_Valid_7_delay_26_26;
    io_A_Valid_7_delay_28_24 <= io_A_Valid_7_delay_27_25;
    io_A_Valid_7_delay_29_23 <= io_A_Valid_7_delay_28_24;
    io_A_Valid_7_delay_30_22 <= io_A_Valid_7_delay_29_23;
    io_A_Valid_7_delay_31_21 <= io_A_Valid_7_delay_30_22;
    io_A_Valid_7_delay_32_20 <= io_A_Valid_7_delay_31_21;
    io_A_Valid_7_delay_33_19 <= io_A_Valid_7_delay_32_20;
    io_A_Valid_7_delay_34_18 <= io_A_Valid_7_delay_33_19;
    io_A_Valid_7_delay_35_17 <= io_A_Valid_7_delay_34_18;
    io_A_Valid_7_delay_36_16 <= io_A_Valid_7_delay_35_17;
    io_A_Valid_7_delay_37_15 <= io_A_Valid_7_delay_36_16;
    io_A_Valid_7_delay_38_14 <= io_A_Valid_7_delay_37_15;
    io_A_Valid_7_delay_39_13 <= io_A_Valid_7_delay_38_14;
    io_A_Valid_7_delay_40_12 <= io_A_Valid_7_delay_39_13;
    io_A_Valid_7_delay_41_11 <= io_A_Valid_7_delay_40_12;
    io_A_Valid_7_delay_42_10 <= io_A_Valid_7_delay_41_11;
    io_A_Valid_7_delay_43_9 <= io_A_Valid_7_delay_42_10;
    io_A_Valid_7_delay_44_8 <= io_A_Valid_7_delay_43_9;
    io_A_Valid_7_delay_45_7 <= io_A_Valid_7_delay_44_8;
    io_A_Valid_7_delay_46_6 <= io_A_Valid_7_delay_45_7;
    io_A_Valid_7_delay_47_5 <= io_A_Valid_7_delay_46_6;
    io_A_Valid_7_delay_48_4 <= io_A_Valid_7_delay_47_5;
    io_A_Valid_7_delay_49_3 <= io_A_Valid_7_delay_48_4;
    io_A_Valid_7_delay_50_2 <= io_A_Valid_7_delay_49_3;
    io_A_Valid_7_delay_51_1 <= io_A_Valid_7_delay_50_2;
    io_A_Valid_7_delay_52 <= io_A_Valid_7_delay_51_1;
    io_B_Valid_52_delay_1_6 <= io_B_Valid_52;
    io_B_Valid_52_delay_2_5 <= io_B_Valid_52_delay_1_6;
    io_B_Valid_52_delay_3_4 <= io_B_Valid_52_delay_2_5;
    io_B_Valid_52_delay_4_3 <= io_B_Valid_52_delay_3_4;
    io_B_Valid_52_delay_5_2 <= io_B_Valid_52_delay_4_3;
    io_B_Valid_52_delay_6_1 <= io_B_Valid_52_delay_5_2;
    io_B_Valid_52_delay_7 <= io_B_Valid_52_delay_6_1;
    io_A_Valid_7_delay_1_52 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_51 <= io_A_Valid_7_delay_1_52;
    io_A_Valid_7_delay_3_50 <= io_A_Valid_7_delay_2_51;
    io_A_Valid_7_delay_4_49 <= io_A_Valid_7_delay_3_50;
    io_A_Valid_7_delay_5_48 <= io_A_Valid_7_delay_4_49;
    io_A_Valid_7_delay_6_47 <= io_A_Valid_7_delay_5_48;
    io_A_Valid_7_delay_7_46 <= io_A_Valid_7_delay_6_47;
    io_A_Valid_7_delay_8_45 <= io_A_Valid_7_delay_7_46;
    io_A_Valid_7_delay_9_44 <= io_A_Valid_7_delay_8_45;
    io_A_Valid_7_delay_10_43 <= io_A_Valid_7_delay_9_44;
    io_A_Valid_7_delay_11_42 <= io_A_Valid_7_delay_10_43;
    io_A_Valid_7_delay_12_41 <= io_A_Valid_7_delay_11_42;
    io_A_Valid_7_delay_13_40 <= io_A_Valid_7_delay_12_41;
    io_A_Valid_7_delay_14_39 <= io_A_Valid_7_delay_13_40;
    io_A_Valid_7_delay_15_38 <= io_A_Valid_7_delay_14_39;
    io_A_Valid_7_delay_16_37 <= io_A_Valid_7_delay_15_38;
    io_A_Valid_7_delay_17_36 <= io_A_Valid_7_delay_16_37;
    io_A_Valid_7_delay_18_35 <= io_A_Valid_7_delay_17_36;
    io_A_Valid_7_delay_19_34 <= io_A_Valid_7_delay_18_35;
    io_A_Valid_7_delay_20_33 <= io_A_Valid_7_delay_19_34;
    io_A_Valid_7_delay_21_32 <= io_A_Valid_7_delay_20_33;
    io_A_Valid_7_delay_22_31 <= io_A_Valid_7_delay_21_32;
    io_A_Valid_7_delay_23_30 <= io_A_Valid_7_delay_22_31;
    io_A_Valid_7_delay_24_29 <= io_A_Valid_7_delay_23_30;
    io_A_Valid_7_delay_25_28 <= io_A_Valid_7_delay_24_29;
    io_A_Valid_7_delay_26_27 <= io_A_Valid_7_delay_25_28;
    io_A_Valid_7_delay_27_26 <= io_A_Valid_7_delay_26_27;
    io_A_Valid_7_delay_28_25 <= io_A_Valid_7_delay_27_26;
    io_A_Valid_7_delay_29_24 <= io_A_Valid_7_delay_28_25;
    io_A_Valid_7_delay_30_23 <= io_A_Valid_7_delay_29_24;
    io_A_Valid_7_delay_31_22 <= io_A_Valid_7_delay_30_23;
    io_A_Valid_7_delay_32_21 <= io_A_Valid_7_delay_31_22;
    io_A_Valid_7_delay_33_20 <= io_A_Valid_7_delay_32_21;
    io_A_Valid_7_delay_34_19 <= io_A_Valid_7_delay_33_20;
    io_A_Valid_7_delay_35_18 <= io_A_Valid_7_delay_34_19;
    io_A_Valid_7_delay_36_17 <= io_A_Valid_7_delay_35_18;
    io_A_Valid_7_delay_37_16 <= io_A_Valid_7_delay_36_17;
    io_A_Valid_7_delay_38_15 <= io_A_Valid_7_delay_37_16;
    io_A_Valid_7_delay_39_14 <= io_A_Valid_7_delay_38_15;
    io_A_Valid_7_delay_40_13 <= io_A_Valid_7_delay_39_14;
    io_A_Valid_7_delay_41_12 <= io_A_Valid_7_delay_40_13;
    io_A_Valid_7_delay_42_11 <= io_A_Valid_7_delay_41_12;
    io_A_Valid_7_delay_43_10 <= io_A_Valid_7_delay_42_11;
    io_A_Valid_7_delay_44_9 <= io_A_Valid_7_delay_43_10;
    io_A_Valid_7_delay_45_8 <= io_A_Valid_7_delay_44_9;
    io_A_Valid_7_delay_46_7 <= io_A_Valid_7_delay_45_8;
    io_A_Valid_7_delay_47_6 <= io_A_Valid_7_delay_46_7;
    io_A_Valid_7_delay_48_5 <= io_A_Valid_7_delay_47_6;
    io_A_Valid_7_delay_49_4 <= io_A_Valid_7_delay_48_5;
    io_A_Valid_7_delay_50_3 <= io_A_Valid_7_delay_49_4;
    io_A_Valid_7_delay_51_2 <= io_A_Valid_7_delay_50_3;
    io_A_Valid_7_delay_52_1 <= io_A_Valid_7_delay_51_2;
    io_A_Valid_7_delay_53 <= io_A_Valid_7_delay_52_1;
    io_B_Valid_53_delay_1_6 <= io_B_Valid_53;
    io_B_Valid_53_delay_2_5 <= io_B_Valid_53_delay_1_6;
    io_B_Valid_53_delay_3_4 <= io_B_Valid_53_delay_2_5;
    io_B_Valid_53_delay_4_3 <= io_B_Valid_53_delay_3_4;
    io_B_Valid_53_delay_5_2 <= io_B_Valid_53_delay_4_3;
    io_B_Valid_53_delay_6_1 <= io_B_Valid_53_delay_5_2;
    io_B_Valid_53_delay_7 <= io_B_Valid_53_delay_6_1;
    io_A_Valid_7_delay_1_53 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_52 <= io_A_Valid_7_delay_1_53;
    io_A_Valid_7_delay_3_51 <= io_A_Valid_7_delay_2_52;
    io_A_Valid_7_delay_4_50 <= io_A_Valid_7_delay_3_51;
    io_A_Valid_7_delay_5_49 <= io_A_Valid_7_delay_4_50;
    io_A_Valid_7_delay_6_48 <= io_A_Valid_7_delay_5_49;
    io_A_Valid_7_delay_7_47 <= io_A_Valid_7_delay_6_48;
    io_A_Valid_7_delay_8_46 <= io_A_Valid_7_delay_7_47;
    io_A_Valid_7_delay_9_45 <= io_A_Valid_7_delay_8_46;
    io_A_Valid_7_delay_10_44 <= io_A_Valid_7_delay_9_45;
    io_A_Valid_7_delay_11_43 <= io_A_Valid_7_delay_10_44;
    io_A_Valid_7_delay_12_42 <= io_A_Valid_7_delay_11_43;
    io_A_Valid_7_delay_13_41 <= io_A_Valid_7_delay_12_42;
    io_A_Valid_7_delay_14_40 <= io_A_Valid_7_delay_13_41;
    io_A_Valid_7_delay_15_39 <= io_A_Valid_7_delay_14_40;
    io_A_Valid_7_delay_16_38 <= io_A_Valid_7_delay_15_39;
    io_A_Valid_7_delay_17_37 <= io_A_Valid_7_delay_16_38;
    io_A_Valid_7_delay_18_36 <= io_A_Valid_7_delay_17_37;
    io_A_Valid_7_delay_19_35 <= io_A_Valid_7_delay_18_36;
    io_A_Valid_7_delay_20_34 <= io_A_Valid_7_delay_19_35;
    io_A_Valid_7_delay_21_33 <= io_A_Valid_7_delay_20_34;
    io_A_Valid_7_delay_22_32 <= io_A_Valid_7_delay_21_33;
    io_A_Valid_7_delay_23_31 <= io_A_Valid_7_delay_22_32;
    io_A_Valid_7_delay_24_30 <= io_A_Valid_7_delay_23_31;
    io_A_Valid_7_delay_25_29 <= io_A_Valid_7_delay_24_30;
    io_A_Valid_7_delay_26_28 <= io_A_Valid_7_delay_25_29;
    io_A_Valid_7_delay_27_27 <= io_A_Valid_7_delay_26_28;
    io_A_Valid_7_delay_28_26 <= io_A_Valid_7_delay_27_27;
    io_A_Valid_7_delay_29_25 <= io_A_Valid_7_delay_28_26;
    io_A_Valid_7_delay_30_24 <= io_A_Valid_7_delay_29_25;
    io_A_Valid_7_delay_31_23 <= io_A_Valid_7_delay_30_24;
    io_A_Valid_7_delay_32_22 <= io_A_Valid_7_delay_31_23;
    io_A_Valid_7_delay_33_21 <= io_A_Valid_7_delay_32_22;
    io_A_Valid_7_delay_34_20 <= io_A_Valid_7_delay_33_21;
    io_A_Valid_7_delay_35_19 <= io_A_Valid_7_delay_34_20;
    io_A_Valid_7_delay_36_18 <= io_A_Valid_7_delay_35_19;
    io_A_Valid_7_delay_37_17 <= io_A_Valid_7_delay_36_18;
    io_A_Valid_7_delay_38_16 <= io_A_Valid_7_delay_37_17;
    io_A_Valid_7_delay_39_15 <= io_A_Valid_7_delay_38_16;
    io_A_Valid_7_delay_40_14 <= io_A_Valid_7_delay_39_15;
    io_A_Valid_7_delay_41_13 <= io_A_Valid_7_delay_40_14;
    io_A_Valid_7_delay_42_12 <= io_A_Valid_7_delay_41_13;
    io_A_Valid_7_delay_43_11 <= io_A_Valid_7_delay_42_12;
    io_A_Valid_7_delay_44_10 <= io_A_Valid_7_delay_43_11;
    io_A_Valid_7_delay_45_9 <= io_A_Valid_7_delay_44_10;
    io_A_Valid_7_delay_46_8 <= io_A_Valid_7_delay_45_9;
    io_A_Valid_7_delay_47_7 <= io_A_Valid_7_delay_46_8;
    io_A_Valid_7_delay_48_6 <= io_A_Valid_7_delay_47_7;
    io_A_Valid_7_delay_49_5 <= io_A_Valid_7_delay_48_6;
    io_A_Valid_7_delay_50_4 <= io_A_Valid_7_delay_49_5;
    io_A_Valid_7_delay_51_3 <= io_A_Valid_7_delay_50_4;
    io_A_Valid_7_delay_52_2 <= io_A_Valid_7_delay_51_3;
    io_A_Valid_7_delay_53_1 <= io_A_Valid_7_delay_52_2;
    io_A_Valid_7_delay_54 <= io_A_Valid_7_delay_53_1;
    io_B_Valid_54_delay_1_6 <= io_B_Valid_54;
    io_B_Valid_54_delay_2_5 <= io_B_Valid_54_delay_1_6;
    io_B_Valid_54_delay_3_4 <= io_B_Valid_54_delay_2_5;
    io_B_Valid_54_delay_4_3 <= io_B_Valid_54_delay_3_4;
    io_B_Valid_54_delay_5_2 <= io_B_Valid_54_delay_4_3;
    io_B_Valid_54_delay_6_1 <= io_B_Valid_54_delay_5_2;
    io_B_Valid_54_delay_7 <= io_B_Valid_54_delay_6_1;
    io_A_Valid_7_delay_1_54 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_53 <= io_A_Valid_7_delay_1_54;
    io_A_Valid_7_delay_3_52 <= io_A_Valid_7_delay_2_53;
    io_A_Valid_7_delay_4_51 <= io_A_Valid_7_delay_3_52;
    io_A_Valid_7_delay_5_50 <= io_A_Valid_7_delay_4_51;
    io_A_Valid_7_delay_6_49 <= io_A_Valid_7_delay_5_50;
    io_A_Valid_7_delay_7_48 <= io_A_Valid_7_delay_6_49;
    io_A_Valid_7_delay_8_47 <= io_A_Valid_7_delay_7_48;
    io_A_Valid_7_delay_9_46 <= io_A_Valid_7_delay_8_47;
    io_A_Valid_7_delay_10_45 <= io_A_Valid_7_delay_9_46;
    io_A_Valid_7_delay_11_44 <= io_A_Valid_7_delay_10_45;
    io_A_Valid_7_delay_12_43 <= io_A_Valid_7_delay_11_44;
    io_A_Valid_7_delay_13_42 <= io_A_Valid_7_delay_12_43;
    io_A_Valid_7_delay_14_41 <= io_A_Valid_7_delay_13_42;
    io_A_Valid_7_delay_15_40 <= io_A_Valid_7_delay_14_41;
    io_A_Valid_7_delay_16_39 <= io_A_Valid_7_delay_15_40;
    io_A_Valid_7_delay_17_38 <= io_A_Valid_7_delay_16_39;
    io_A_Valid_7_delay_18_37 <= io_A_Valid_7_delay_17_38;
    io_A_Valid_7_delay_19_36 <= io_A_Valid_7_delay_18_37;
    io_A_Valid_7_delay_20_35 <= io_A_Valid_7_delay_19_36;
    io_A_Valid_7_delay_21_34 <= io_A_Valid_7_delay_20_35;
    io_A_Valid_7_delay_22_33 <= io_A_Valid_7_delay_21_34;
    io_A_Valid_7_delay_23_32 <= io_A_Valid_7_delay_22_33;
    io_A_Valid_7_delay_24_31 <= io_A_Valid_7_delay_23_32;
    io_A_Valid_7_delay_25_30 <= io_A_Valid_7_delay_24_31;
    io_A_Valid_7_delay_26_29 <= io_A_Valid_7_delay_25_30;
    io_A_Valid_7_delay_27_28 <= io_A_Valid_7_delay_26_29;
    io_A_Valid_7_delay_28_27 <= io_A_Valid_7_delay_27_28;
    io_A_Valid_7_delay_29_26 <= io_A_Valid_7_delay_28_27;
    io_A_Valid_7_delay_30_25 <= io_A_Valid_7_delay_29_26;
    io_A_Valid_7_delay_31_24 <= io_A_Valid_7_delay_30_25;
    io_A_Valid_7_delay_32_23 <= io_A_Valid_7_delay_31_24;
    io_A_Valid_7_delay_33_22 <= io_A_Valid_7_delay_32_23;
    io_A_Valid_7_delay_34_21 <= io_A_Valid_7_delay_33_22;
    io_A_Valid_7_delay_35_20 <= io_A_Valid_7_delay_34_21;
    io_A_Valid_7_delay_36_19 <= io_A_Valid_7_delay_35_20;
    io_A_Valid_7_delay_37_18 <= io_A_Valid_7_delay_36_19;
    io_A_Valid_7_delay_38_17 <= io_A_Valid_7_delay_37_18;
    io_A_Valid_7_delay_39_16 <= io_A_Valid_7_delay_38_17;
    io_A_Valid_7_delay_40_15 <= io_A_Valid_7_delay_39_16;
    io_A_Valid_7_delay_41_14 <= io_A_Valid_7_delay_40_15;
    io_A_Valid_7_delay_42_13 <= io_A_Valid_7_delay_41_14;
    io_A_Valid_7_delay_43_12 <= io_A_Valid_7_delay_42_13;
    io_A_Valid_7_delay_44_11 <= io_A_Valid_7_delay_43_12;
    io_A_Valid_7_delay_45_10 <= io_A_Valid_7_delay_44_11;
    io_A_Valid_7_delay_46_9 <= io_A_Valid_7_delay_45_10;
    io_A_Valid_7_delay_47_8 <= io_A_Valid_7_delay_46_9;
    io_A_Valid_7_delay_48_7 <= io_A_Valid_7_delay_47_8;
    io_A_Valid_7_delay_49_6 <= io_A_Valid_7_delay_48_7;
    io_A_Valid_7_delay_50_5 <= io_A_Valid_7_delay_49_6;
    io_A_Valid_7_delay_51_4 <= io_A_Valid_7_delay_50_5;
    io_A_Valid_7_delay_52_3 <= io_A_Valid_7_delay_51_4;
    io_A_Valid_7_delay_53_2 <= io_A_Valid_7_delay_52_3;
    io_A_Valid_7_delay_54_1 <= io_A_Valid_7_delay_53_2;
    io_A_Valid_7_delay_55 <= io_A_Valid_7_delay_54_1;
    io_B_Valid_55_delay_1_6 <= io_B_Valid_55;
    io_B_Valid_55_delay_2_5 <= io_B_Valid_55_delay_1_6;
    io_B_Valid_55_delay_3_4 <= io_B_Valid_55_delay_2_5;
    io_B_Valid_55_delay_4_3 <= io_B_Valid_55_delay_3_4;
    io_B_Valid_55_delay_5_2 <= io_B_Valid_55_delay_4_3;
    io_B_Valid_55_delay_6_1 <= io_B_Valid_55_delay_5_2;
    io_B_Valid_55_delay_7 <= io_B_Valid_55_delay_6_1;
    io_A_Valid_7_delay_1_55 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_54 <= io_A_Valid_7_delay_1_55;
    io_A_Valid_7_delay_3_53 <= io_A_Valid_7_delay_2_54;
    io_A_Valid_7_delay_4_52 <= io_A_Valid_7_delay_3_53;
    io_A_Valid_7_delay_5_51 <= io_A_Valid_7_delay_4_52;
    io_A_Valid_7_delay_6_50 <= io_A_Valid_7_delay_5_51;
    io_A_Valid_7_delay_7_49 <= io_A_Valid_7_delay_6_50;
    io_A_Valid_7_delay_8_48 <= io_A_Valid_7_delay_7_49;
    io_A_Valid_7_delay_9_47 <= io_A_Valid_7_delay_8_48;
    io_A_Valid_7_delay_10_46 <= io_A_Valid_7_delay_9_47;
    io_A_Valid_7_delay_11_45 <= io_A_Valid_7_delay_10_46;
    io_A_Valid_7_delay_12_44 <= io_A_Valid_7_delay_11_45;
    io_A_Valid_7_delay_13_43 <= io_A_Valid_7_delay_12_44;
    io_A_Valid_7_delay_14_42 <= io_A_Valid_7_delay_13_43;
    io_A_Valid_7_delay_15_41 <= io_A_Valid_7_delay_14_42;
    io_A_Valid_7_delay_16_40 <= io_A_Valid_7_delay_15_41;
    io_A_Valid_7_delay_17_39 <= io_A_Valid_7_delay_16_40;
    io_A_Valid_7_delay_18_38 <= io_A_Valid_7_delay_17_39;
    io_A_Valid_7_delay_19_37 <= io_A_Valid_7_delay_18_38;
    io_A_Valid_7_delay_20_36 <= io_A_Valid_7_delay_19_37;
    io_A_Valid_7_delay_21_35 <= io_A_Valid_7_delay_20_36;
    io_A_Valid_7_delay_22_34 <= io_A_Valid_7_delay_21_35;
    io_A_Valid_7_delay_23_33 <= io_A_Valid_7_delay_22_34;
    io_A_Valid_7_delay_24_32 <= io_A_Valid_7_delay_23_33;
    io_A_Valid_7_delay_25_31 <= io_A_Valid_7_delay_24_32;
    io_A_Valid_7_delay_26_30 <= io_A_Valid_7_delay_25_31;
    io_A_Valid_7_delay_27_29 <= io_A_Valid_7_delay_26_30;
    io_A_Valid_7_delay_28_28 <= io_A_Valid_7_delay_27_29;
    io_A_Valid_7_delay_29_27 <= io_A_Valid_7_delay_28_28;
    io_A_Valid_7_delay_30_26 <= io_A_Valid_7_delay_29_27;
    io_A_Valid_7_delay_31_25 <= io_A_Valid_7_delay_30_26;
    io_A_Valid_7_delay_32_24 <= io_A_Valid_7_delay_31_25;
    io_A_Valid_7_delay_33_23 <= io_A_Valid_7_delay_32_24;
    io_A_Valid_7_delay_34_22 <= io_A_Valid_7_delay_33_23;
    io_A_Valid_7_delay_35_21 <= io_A_Valid_7_delay_34_22;
    io_A_Valid_7_delay_36_20 <= io_A_Valid_7_delay_35_21;
    io_A_Valid_7_delay_37_19 <= io_A_Valid_7_delay_36_20;
    io_A_Valid_7_delay_38_18 <= io_A_Valid_7_delay_37_19;
    io_A_Valid_7_delay_39_17 <= io_A_Valid_7_delay_38_18;
    io_A_Valid_7_delay_40_16 <= io_A_Valid_7_delay_39_17;
    io_A_Valid_7_delay_41_15 <= io_A_Valid_7_delay_40_16;
    io_A_Valid_7_delay_42_14 <= io_A_Valid_7_delay_41_15;
    io_A_Valid_7_delay_43_13 <= io_A_Valid_7_delay_42_14;
    io_A_Valid_7_delay_44_12 <= io_A_Valid_7_delay_43_13;
    io_A_Valid_7_delay_45_11 <= io_A_Valid_7_delay_44_12;
    io_A_Valid_7_delay_46_10 <= io_A_Valid_7_delay_45_11;
    io_A_Valid_7_delay_47_9 <= io_A_Valid_7_delay_46_10;
    io_A_Valid_7_delay_48_8 <= io_A_Valid_7_delay_47_9;
    io_A_Valid_7_delay_49_7 <= io_A_Valid_7_delay_48_8;
    io_A_Valid_7_delay_50_6 <= io_A_Valid_7_delay_49_7;
    io_A_Valid_7_delay_51_5 <= io_A_Valid_7_delay_50_6;
    io_A_Valid_7_delay_52_4 <= io_A_Valid_7_delay_51_5;
    io_A_Valid_7_delay_53_3 <= io_A_Valid_7_delay_52_4;
    io_A_Valid_7_delay_54_2 <= io_A_Valid_7_delay_53_3;
    io_A_Valid_7_delay_55_1 <= io_A_Valid_7_delay_54_2;
    io_A_Valid_7_delay_56 <= io_A_Valid_7_delay_55_1;
    io_B_Valid_56_delay_1_6 <= io_B_Valid_56;
    io_B_Valid_56_delay_2_5 <= io_B_Valid_56_delay_1_6;
    io_B_Valid_56_delay_3_4 <= io_B_Valid_56_delay_2_5;
    io_B_Valid_56_delay_4_3 <= io_B_Valid_56_delay_3_4;
    io_B_Valid_56_delay_5_2 <= io_B_Valid_56_delay_4_3;
    io_B_Valid_56_delay_6_1 <= io_B_Valid_56_delay_5_2;
    io_B_Valid_56_delay_7 <= io_B_Valid_56_delay_6_1;
    io_A_Valid_7_delay_1_56 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_55 <= io_A_Valid_7_delay_1_56;
    io_A_Valid_7_delay_3_54 <= io_A_Valid_7_delay_2_55;
    io_A_Valid_7_delay_4_53 <= io_A_Valid_7_delay_3_54;
    io_A_Valid_7_delay_5_52 <= io_A_Valid_7_delay_4_53;
    io_A_Valid_7_delay_6_51 <= io_A_Valid_7_delay_5_52;
    io_A_Valid_7_delay_7_50 <= io_A_Valid_7_delay_6_51;
    io_A_Valid_7_delay_8_49 <= io_A_Valid_7_delay_7_50;
    io_A_Valid_7_delay_9_48 <= io_A_Valid_7_delay_8_49;
    io_A_Valid_7_delay_10_47 <= io_A_Valid_7_delay_9_48;
    io_A_Valid_7_delay_11_46 <= io_A_Valid_7_delay_10_47;
    io_A_Valid_7_delay_12_45 <= io_A_Valid_7_delay_11_46;
    io_A_Valid_7_delay_13_44 <= io_A_Valid_7_delay_12_45;
    io_A_Valid_7_delay_14_43 <= io_A_Valid_7_delay_13_44;
    io_A_Valid_7_delay_15_42 <= io_A_Valid_7_delay_14_43;
    io_A_Valid_7_delay_16_41 <= io_A_Valid_7_delay_15_42;
    io_A_Valid_7_delay_17_40 <= io_A_Valid_7_delay_16_41;
    io_A_Valid_7_delay_18_39 <= io_A_Valid_7_delay_17_40;
    io_A_Valid_7_delay_19_38 <= io_A_Valid_7_delay_18_39;
    io_A_Valid_7_delay_20_37 <= io_A_Valid_7_delay_19_38;
    io_A_Valid_7_delay_21_36 <= io_A_Valid_7_delay_20_37;
    io_A_Valid_7_delay_22_35 <= io_A_Valid_7_delay_21_36;
    io_A_Valid_7_delay_23_34 <= io_A_Valid_7_delay_22_35;
    io_A_Valid_7_delay_24_33 <= io_A_Valid_7_delay_23_34;
    io_A_Valid_7_delay_25_32 <= io_A_Valid_7_delay_24_33;
    io_A_Valid_7_delay_26_31 <= io_A_Valid_7_delay_25_32;
    io_A_Valid_7_delay_27_30 <= io_A_Valid_7_delay_26_31;
    io_A_Valid_7_delay_28_29 <= io_A_Valid_7_delay_27_30;
    io_A_Valid_7_delay_29_28 <= io_A_Valid_7_delay_28_29;
    io_A_Valid_7_delay_30_27 <= io_A_Valid_7_delay_29_28;
    io_A_Valid_7_delay_31_26 <= io_A_Valid_7_delay_30_27;
    io_A_Valid_7_delay_32_25 <= io_A_Valid_7_delay_31_26;
    io_A_Valid_7_delay_33_24 <= io_A_Valid_7_delay_32_25;
    io_A_Valid_7_delay_34_23 <= io_A_Valid_7_delay_33_24;
    io_A_Valid_7_delay_35_22 <= io_A_Valid_7_delay_34_23;
    io_A_Valid_7_delay_36_21 <= io_A_Valid_7_delay_35_22;
    io_A_Valid_7_delay_37_20 <= io_A_Valid_7_delay_36_21;
    io_A_Valid_7_delay_38_19 <= io_A_Valid_7_delay_37_20;
    io_A_Valid_7_delay_39_18 <= io_A_Valid_7_delay_38_19;
    io_A_Valid_7_delay_40_17 <= io_A_Valid_7_delay_39_18;
    io_A_Valid_7_delay_41_16 <= io_A_Valid_7_delay_40_17;
    io_A_Valid_7_delay_42_15 <= io_A_Valid_7_delay_41_16;
    io_A_Valid_7_delay_43_14 <= io_A_Valid_7_delay_42_15;
    io_A_Valid_7_delay_44_13 <= io_A_Valid_7_delay_43_14;
    io_A_Valid_7_delay_45_12 <= io_A_Valid_7_delay_44_13;
    io_A_Valid_7_delay_46_11 <= io_A_Valid_7_delay_45_12;
    io_A_Valid_7_delay_47_10 <= io_A_Valid_7_delay_46_11;
    io_A_Valid_7_delay_48_9 <= io_A_Valid_7_delay_47_10;
    io_A_Valid_7_delay_49_8 <= io_A_Valid_7_delay_48_9;
    io_A_Valid_7_delay_50_7 <= io_A_Valid_7_delay_49_8;
    io_A_Valid_7_delay_51_6 <= io_A_Valid_7_delay_50_7;
    io_A_Valid_7_delay_52_5 <= io_A_Valid_7_delay_51_6;
    io_A_Valid_7_delay_53_4 <= io_A_Valid_7_delay_52_5;
    io_A_Valid_7_delay_54_3 <= io_A_Valid_7_delay_53_4;
    io_A_Valid_7_delay_55_2 <= io_A_Valid_7_delay_54_3;
    io_A_Valid_7_delay_56_1 <= io_A_Valid_7_delay_55_2;
    io_A_Valid_7_delay_57 <= io_A_Valid_7_delay_56_1;
    io_B_Valid_57_delay_1_6 <= io_B_Valid_57;
    io_B_Valid_57_delay_2_5 <= io_B_Valid_57_delay_1_6;
    io_B_Valid_57_delay_3_4 <= io_B_Valid_57_delay_2_5;
    io_B_Valid_57_delay_4_3 <= io_B_Valid_57_delay_3_4;
    io_B_Valid_57_delay_5_2 <= io_B_Valid_57_delay_4_3;
    io_B_Valid_57_delay_6_1 <= io_B_Valid_57_delay_5_2;
    io_B_Valid_57_delay_7 <= io_B_Valid_57_delay_6_1;
    io_A_Valid_7_delay_1_57 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_56 <= io_A_Valid_7_delay_1_57;
    io_A_Valid_7_delay_3_55 <= io_A_Valid_7_delay_2_56;
    io_A_Valid_7_delay_4_54 <= io_A_Valid_7_delay_3_55;
    io_A_Valid_7_delay_5_53 <= io_A_Valid_7_delay_4_54;
    io_A_Valid_7_delay_6_52 <= io_A_Valid_7_delay_5_53;
    io_A_Valid_7_delay_7_51 <= io_A_Valid_7_delay_6_52;
    io_A_Valid_7_delay_8_50 <= io_A_Valid_7_delay_7_51;
    io_A_Valid_7_delay_9_49 <= io_A_Valid_7_delay_8_50;
    io_A_Valid_7_delay_10_48 <= io_A_Valid_7_delay_9_49;
    io_A_Valid_7_delay_11_47 <= io_A_Valid_7_delay_10_48;
    io_A_Valid_7_delay_12_46 <= io_A_Valid_7_delay_11_47;
    io_A_Valid_7_delay_13_45 <= io_A_Valid_7_delay_12_46;
    io_A_Valid_7_delay_14_44 <= io_A_Valid_7_delay_13_45;
    io_A_Valid_7_delay_15_43 <= io_A_Valid_7_delay_14_44;
    io_A_Valid_7_delay_16_42 <= io_A_Valid_7_delay_15_43;
    io_A_Valid_7_delay_17_41 <= io_A_Valid_7_delay_16_42;
    io_A_Valid_7_delay_18_40 <= io_A_Valid_7_delay_17_41;
    io_A_Valid_7_delay_19_39 <= io_A_Valid_7_delay_18_40;
    io_A_Valid_7_delay_20_38 <= io_A_Valid_7_delay_19_39;
    io_A_Valid_7_delay_21_37 <= io_A_Valid_7_delay_20_38;
    io_A_Valid_7_delay_22_36 <= io_A_Valid_7_delay_21_37;
    io_A_Valid_7_delay_23_35 <= io_A_Valid_7_delay_22_36;
    io_A_Valid_7_delay_24_34 <= io_A_Valid_7_delay_23_35;
    io_A_Valid_7_delay_25_33 <= io_A_Valid_7_delay_24_34;
    io_A_Valid_7_delay_26_32 <= io_A_Valid_7_delay_25_33;
    io_A_Valid_7_delay_27_31 <= io_A_Valid_7_delay_26_32;
    io_A_Valid_7_delay_28_30 <= io_A_Valid_7_delay_27_31;
    io_A_Valid_7_delay_29_29 <= io_A_Valid_7_delay_28_30;
    io_A_Valid_7_delay_30_28 <= io_A_Valid_7_delay_29_29;
    io_A_Valid_7_delay_31_27 <= io_A_Valid_7_delay_30_28;
    io_A_Valid_7_delay_32_26 <= io_A_Valid_7_delay_31_27;
    io_A_Valid_7_delay_33_25 <= io_A_Valid_7_delay_32_26;
    io_A_Valid_7_delay_34_24 <= io_A_Valid_7_delay_33_25;
    io_A_Valid_7_delay_35_23 <= io_A_Valid_7_delay_34_24;
    io_A_Valid_7_delay_36_22 <= io_A_Valid_7_delay_35_23;
    io_A_Valid_7_delay_37_21 <= io_A_Valid_7_delay_36_22;
    io_A_Valid_7_delay_38_20 <= io_A_Valid_7_delay_37_21;
    io_A_Valid_7_delay_39_19 <= io_A_Valid_7_delay_38_20;
    io_A_Valid_7_delay_40_18 <= io_A_Valid_7_delay_39_19;
    io_A_Valid_7_delay_41_17 <= io_A_Valid_7_delay_40_18;
    io_A_Valid_7_delay_42_16 <= io_A_Valid_7_delay_41_17;
    io_A_Valid_7_delay_43_15 <= io_A_Valid_7_delay_42_16;
    io_A_Valid_7_delay_44_14 <= io_A_Valid_7_delay_43_15;
    io_A_Valid_7_delay_45_13 <= io_A_Valid_7_delay_44_14;
    io_A_Valid_7_delay_46_12 <= io_A_Valid_7_delay_45_13;
    io_A_Valid_7_delay_47_11 <= io_A_Valid_7_delay_46_12;
    io_A_Valid_7_delay_48_10 <= io_A_Valid_7_delay_47_11;
    io_A_Valid_7_delay_49_9 <= io_A_Valid_7_delay_48_10;
    io_A_Valid_7_delay_50_8 <= io_A_Valid_7_delay_49_9;
    io_A_Valid_7_delay_51_7 <= io_A_Valid_7_delay_50_8;
    io_A_Valid_7_delay_52_6 <= io_A_Valid_7_delay_51_7;
    io_A_Valid_7_delay_53_5 <= io_A_Valid_7_delay_52_6;
    io_A_Valid_7_delay_54_4 <= io_A_Valid_7_delay_53_5;
    io_A_Valid_7_delay_55_3 <= io_A_Valid_7_delay_54_4;
    io_A_Valid_7_delay_56_2 <= io_A_Valid_7_delay_55_3;
    io_A_Valid_7_delay_57_1 <= io_A_Valid_7_delay_56_2;
    io_A_Valid_7_delay_58 <= io_A_Valid_7_delay_57_1;
    io_B_Valid_58_delay_1_6 <= io_B_Valid_58;
    io_B_Valid_58_delay_2_5 <= io_B_Valid_58_delay_1_6;
    io_B_Valid_58_delay_3_4 <= io_B_Valid_58_delay_2_5;
    io_B_Valid_58_delay_4_3 <= io_B_Valid_58_delay_3_4;
    io_B_Valid_58_delay_5_2 <= io_B_Valid_58_delay_4_3;
    io_B_Valid_58_delay_6_1 <= io_B_Valid_58_delay_5_2;
    io_B_Valid_58_delay_7 <= io_B_Valid_58_delay_6_1;
    io_A_Valid_7_delay_1_58 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_57 <= io_A_Valid_7_delay_1_58;
    io_A_Valid_7_delay_3_56 <= io_A_Valid_7_delay_2_57;
    io_A_Valid_7_delay_4_55 <= io_A_Valid_7_delay_3_56;
    io_A_Valid_7_delay_5_54 <= io_A_Valid_7_delay_4_55;
    io_A_Valid_7_delay_6_53 <= io_A_Valid_7_delay_5_54;
    io_A_Valid_7_delay_7_52 <= io_A_Valid_7_delay_6_53;
    io_A_Valid_7_delay_8_51 <= io_A_Valid_7_delay_7_52;
    io_A_Valid_7_delay_9_50 <= io_A_Valid_7_delay_8_51;
    io_A_Valid_7_delay_10_49 <= io_A_Valid_7_delay_9_50;
    io_A_Valid_7_delay_11_48 <= io_A_Valid_7_delay_10_49;
    io_A_Valid_7_delay_12_47 <= io_A_Valid_7_delay_11_48;
    io_A_Valid_7_delay_13_46 <= io_A_Valid_7_delay_12_47;
    io_A_Valid_7_delay_14_45 <= io_A_Valid_7_delay_13_46;
    io_A_Valid_7_delay_15_44 <= io_A_Valid_7_delay_14_45;
    io_A_Valid_7_delay_16_43 <= io_A_Valid_7_delay_15_44;
    io_A_Valid_7_delay_17_42 <= io_A_Valid_7_delay_16_43;
    io_A_Valid_7_delay_18_41 <= io_A_Valid_7_delay_17_42;
    io_A_Valid_7_delay_19_40 <= io_A_Valid_7_delay_18_41;
    io_A_Valid_7_delay_20_39 <= io_A_Valid_7_delay_19_40;
    io_A_Valid_7_delay_21_38 <= io_A_Valid_7_delay_20_39;
    io_A_Valid_7_delay_22_37 <= io_A_Valid_7_delay_21_38;
    io_A_Valid_7_delay_23_36 <= io_A_Valid_7_delay_22_37;
    io_A_Valid_7_delay_24_35 <= io_A_Valid_7_delay_23_36;
    io_A_Valid_7_delay_25_34 <= io_A_Valid_7_delay_24_35;
    io_A_Valid_7_delay_26_33 <= io_A_Valid_7_delay_25_34;
    io_A_Valid_7_delay_27_32 <= io_A_Valid_7_delay_26_33;
    io_A_Valid_7_delay_28_31 <= io_A_Valid_7_delay_27_32;
    io_A_Valid_7_delay_29_30 <= io_A_Valid_7_delay_28_31;
    io_A_Valid_7_delay_30_29 <= io_A_Valid_7_delay_29_30;
    io_A_Valid_7_delay_31_28 <= io_A_Valid_7_delay_30_29;
    io_A_Valid_7_delay_32_27 <= io_A_Valid_7_delay_31_28;
    io_A_Valid_7_delay_33_26 <= io_A_Valid_7_delay_32_27;
    io_A_Valid_7_delay_34_25 <= io_A_Valid_7_delay_33_26;
    io_A_Valid_7_delay_35_24 <= io_A_Valid_7_delay_34_25;
    io_A_Valid_7_delay_36_23 <= io_A_Valid_7_delay_35_24;
    io_A_Valid_7_delay_37_22 <= io_A_Valid_7_delay_36_23;
    io_A_Valid_7_delay_38_21 <= io_A_Valid_7_delay_37_22;
    io_A_Valid_7_delay_39_20 <= io_A_Valid_7_delay_38_21;
    io_A_Valid_7_delay_40_19 <= io_A_Valid_7_delay_39_20;
    io_A_Valid_7_delay_41_18 <= io_A_Valid_7_delay_40_19;
    io_A_Valid_7_delay_42_17 <= io_A_Valid_7_delay_41_18;
    io_A_Valid_7_delay_43_16 <= io_A_Valid_7_delay_42_17;
    io_A_Valid_7_delay_44_15 <= io_A_Valid_7_delay_43_16;
    io_A_Valid_7_delay_45_14 <= io_A_Valid_7_delay_44_15;
    io_A_Valid_7_delay_46_13 <= io_A_Valid_7_delay_45_14;
    io_A_Valid_7_delay_47_12 <= io_A_Valid_7_delay_46_13;
    io_A_Valid_7_delay_48_11 <= io_A_Valid_7_delay_47_12;
    io_A_Valid_7_delay_49_10 <= io_A_Valid_7_delay_48_11;
    io_A_Valid_7_delay_50_9 <= io_A_Valid_7_delay_49_10;
    io_A_Valid_7_delay_51_8 <= io_A_Valid_7_delay_50_9;
    io_A_Valid_7_delay_52_7 <= io_A_Valid_7_delay_51_8;
    io_A_Valid_7_delay_53_6 <= io_A_Valid_7_delay_52_7;
    io_A_Valid_7_delay_54_5 <= io_A_Valid_7_delay_53_6;
    io_A_Valid_7_delay_55_4 <= io_A_Valid_7_delay_54_5;
    io_A_Valid_7_delay_56_3 <= io_A_Valid_7_delay_55_4;
    io_A_Valid_7_delay_57_2 <= io_A_Valid_7_delay_56_3;
    io_A_Valid_7_delay_58_1 <= io_A_Valid_7_delay_57_2;
    io_A_Valid_7_delay_59 <= io_A_Valid_7_delay_58_1;
    io_B_Valid_59_delay_1_6 <= io_B_Valid_59;
    io_B_Valid_59_delay_2_5 <= io_B_Valid_59_delay_1_6;
    io_B_Valid_59_delay_3_4 <= io_B_Valid_59_delay_2_5;
    io_B_Valid_59_delay_4_3 <= io_B_Valid_59_delay_3_4;
    io_B_Valid_59_delay_5_2 <= io_B_Valid_59_delay_4_3;
    io_B_Valid_59_delay_6_1 <= io_B_Valid_59_delay_5_2;
    io_B_Valid_59_delay_7 <= io_B_Valid_59_delay_6_1;
    io_A_Valid_7_delay_1_59 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_58 <= io_A_Valid_7_delay_1_59;
    io_A_Valid_7_delay_3_57 <= io_A_Valid_7_delay_2_58;
    io_A_Valid_7_delay_4_56 <= io_A_Valid_7_delay_3_57;
    io_A_Valid_7_delay_5_55 <= io_A_Valid_7_delay_4_56;
    io_A_Valid_7_delay_6_54 <= io_A_Valid_7_delay_5_55;
    io_A_Valid_7_delay_7_53 <= io_A_Valid_7_delay_6_54;
    io_A_Valid_7_delay_8_52 <= io_A_Valid_7_delay_7_53;
    io_A_Valid_7_delay_9_51 <= io_A_Valid_7_delay_8_52;
    io_A_Valid_7_delay_10_50 <= io_A_Valid_7_delay_9_51;
    io_A_Valid_7_delay_11_49 <= io_A_Valid_7_delay_10_50;
    io_A_Valid_7_delay_12_48 <= io_A_Valid_7_delay_11_49;
    io_A_Valid_7_delay_13_47 <= io_A_Valid_7_delay_12_48;
    io_A_Valid_7_delay_14_46 <= io_A_Valid_7_delay_13_47;
    io_A_Valid_7_delay_15_45 <= io_A_Valid_7_delay_14_46;
    io_A_Valid_7_delay_16_44 <= io_A_Valid_7_delay_15_45;
    io_A_Valid_7_delay_17_43 <= io_A_Valid_7_delay_16_44;
    io_A_Valid_7_delay_18_42 <= io_A_Valid_7_delay_17_43;
    io_A_Valid_7_delay_19_41 <= io_A_Valid_7_delay_18_42;
    io_A_Valid_7_delay_20_40 <= io_A_Valid_7_delay_19_41;
    io_A_Valid_7_delay_21_39 <= io_A_Valid_7_delay_20_40;
    io_A_Valid_7_delay_22_38 <= io_A_Valid_7_delay_21_39;
    io_A_Valid_7_delay_23_37 <= io_A_Valid_7_delay_22_38;
    io_A_Valid_7_delay_24_36 <= io_A_Valid_7_delay_23_37;
    io_A_Valid_7_delay_25_35 <= io_A_Valid_7_delay_24_36;
    io_A_Valid_7_delay_26_34 <= io_A_Valid_7_delay_25_35;
    io_A_Valid_7_delay_27_33 <= io_A_Valid_7_delay_26_34;
    io_A_Valid_7_delay_28_32 <= io_A_Valid_7_delay_27_33;
    io_A_Valid_7_delay_29_31 <= io_A_Valid_7_delay_28_32;
    io_A_Valid_7_delay_30_30 <= io_A_Valid_7_delay_29_31;
    io_A_Valid_7_delay_31_29 <= io_A_Valid_7_delay_30_30;
    io_A_Valid_7_delay_32_28 <= io_A_Valid_7_delay_31_29;
    io_A_Valid_7_delay_33_27 <= io_A_Valid_7_delay_32_28;
    io_A_Valid_7_delay_34_26 <= io_A_Valid_7_delay_33_27;
    io_A_Valid_7_delay_35_25 <= io_A_Valid_7_delay_34_26;
    io_A_Valid_7_delay_36_24 <= io_A_Valid_7_delay_35_25;
    io_A_Valid_7_delay_37_23 <= io_A_Valid_7_delay_36_24;
    io_A_Valid_7_delay_38_22 <= io_A_Valid_7_delay_37_23;
    io_A_Valid_7_delay_39_21 <= io_A_Valid_7_delay_38_22;
    io_A_Valid_7_delay_40_20 <= io_A_Valid_7_delay_39_21;
    io_A_Valid_7_delay_41_19 <= io_A_Valid_7_delay_40_20;
    io_A_Valid_7_delay_42_18 <= io_A_Valid_7_delay_41_19;
    io_A_Valid_7_delay_43_17 <= io_A_Valid_7_delay_42_18;
    io_A_Valid_7_delay_44_16 <= io_A_Valid_7_delay_43_17;
    io_A_Valid_7_delay_45_15 <= io_A_Valid_7_delay_44_16;
    io_A_Valid_7_delay_46_14 <= io_A_Valid_7_delay_45_15;
    io_A_Valid_7_delay_47_13 <= io_A_Valid_7_delay_46_14;
    io_A_Valid_7_delay_48_12 <= io_A_Valid_7_delay_47_13;
    io_A_Valid_7_delay_49_11 <= io_A_Valid_7_delay_48_12;
    io_A_Valid_7_delay_50_10 <= io_A_Valid_7_delay_49_11;
    io_A_Valid_7_delay_51_9 <= io_A_Valid_7_delay_50_10;
    io_A_Valid_7_delay_52_8 <= io_A_Valid_7_delay_51_9;
    io_A_Valid_7_delay_53_7 <= io_A_Valid_7_delay_52_8;
    io_A_Valid_7_delay_54_6 <= io_A_Valid_7_delay_53_7;
    io_A_Valid_7_delay_55_5 <= io_A_Valid_7_delay_54_6;
    io_A_Valid_7_delay_56_4 <= io_A_Valid_7_delay_55_5;
    io_A_Valid_7_delay_57_3 <= io_A_Valid_7_delay_56_4;
    io_A_Valid_7_delay_58_2 <= io_A_Valid_7_delay_57_3;
    io_A_Valid_7_delay_59_1 <= io_A_Valid_7_delay_58_2;
    io_A_Valid_7_delay_60 <= io_A_Valid_7_delay_59_1;
    io_B_Valid_60_delay_1_6 <= io_B_Valid_60;
    io_B_Valid_60_delay_2_5 <= io_B_Valid_60_delay_1_6;
    io_B_Valid_60_delay_3_4 <= io_B_Valid_60_delay_2_5;
    io_B_Valid_60_delay_4_3 <= io_B_Valid_60_delay_3_4;
    io_B_Valid_60_delay_5_2 <= io_B_Valid_60_delay_4_3;
    io_B_Valid_60_delay_6_1 <= io_B_Valid_60_delay_5_2;
    io_B_Valid_60_delay_7 <= io_B_Valid_60_delay_6_1;
    io_A_Valid_7_delay_1_60 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_59 <= io_A_Valid_7_delay_1_60;
    io_A_Valid_7_delay_3_58 <= io_A_Valid_7_delay_2_59;
    io_A_Valid_7_delay_4_57 <= io_A_Valid_7_delay_3_58;
    io_A_Valid_7_delay_5_56 <= io_A_Valid_7_delay_4_57;
    io_A_Valid_7_delay_6_55 <= io_A_Valid_7_delay_5_56;
    io_A_Valid_7_delay_7_54 <= io_A_Valid_7_delay_6_55;
    io_A_Valid_7_delay_8_53 <= io_A_Valid_7_delay_7_54;
    io_A_Valid_7_delay_9_52 <= io_A_Valid_7_delay_8_53;
    io_A_Valid_7_delay_10_51 <= io_A_Valid_7_delay_9_52;
    io_A_Valid_7_delay_11_50 <= io_A_Valid_7_delay_10_51;
    io_A_Valid_7_delay_12_49 <= io_A_Valid_7_delay_11_50;
    io_A_Valid_7_delay_13_48 <= io_A_Valid_7_delay_12_49;
    io_A_Valid_7_delay_14_47 <= io_A_Valid_7_delay_13_48;
    io_A_Valid_7_delay_15_46 <= io_A_Valid_7_delay_14_47;
    io_A_Valid_7_delay_16_45 <= io_A_Valid_7_delay_15_46;
    io_A_Valid_7_delay_17_44 <= io_A_Valid_7_delay_16_45;
    io_A_Valid_7_delay_18_43 <= io_A_Valid_7_delay_17_44;
    io_A_Valid_7_delay_19_42 <= io_A_Valid_7_delay_18_43;
    io_A_Valid_7_delay_20_41 <= io_A_Valid_7_delay_19_42;
    io_A_Valid_7_delay_21_40 <= io_A_Valid_7_delay_20_41;
    io_A_Valid_7_delay_22_39 <= io_A_Valid_7_delay_21_40;
    io_A_Valid_7_delay_23_38 <= io_A_Valid_7_delay_22_39;
    io_A_Valid_7_delay_24_37 <= io_A_Valid_7_delay_23_38;
    io_A_Valid_7_delay_25_36 <= io_A_Valid_7_delay_24_37;
    io_A_Valid_7_delay_26_35 <= io_A_Valid_7_delay_25_36;
    io_A_Valid_7_delay_27_34 <= io_A_Valid_7_delay_26_35;
    io_A_Valid_7_delay_28_33 <= io_A_Valid_7_delay_27_34;
    io_A_Valid_7_delay_29_32 <= io_A_Valid_7_delay_28_33;
    io_A_Valid_7_delay_30_31 <= io_A_Valid_7_delay_29_32;
    io_A_Valid_7_delay_31_30 <= io_A_Valid_7_delay_30_31;
    io_A_Valid_7_delay_32_29 <= io_A_Valid_7_delay_31_30;
    io_A_Valid_7_delay_33_28 <= io_A_Valid_7_delay_32_29;
    io_A_Valid_7_delay_34_27 <= io_A_Valid_7_delay_33_28;
    io_A_Valid_7_delay_35_26 <= io_A_Valid_7_delay_34_27;
    io_A_Valid_7_delay_36_25 <= io_A_Valid_7_delay_35_26;
    io_A_Valid_7_delay_37_24 <= io_A_Valid_7_delay_36_25;
    io_A_Valid_7_delay_38_23 <= io_A_Valid_7_delay_37_24;
    io_A_Valid_7_delay_39_22 <= io_A_Valid_7_delay_38_23;
    io_A_Valid_7_delay_40_21 <= io_A_Valid_7_delay_39_22;
    io_A_Valid_7_delay_41_20 <= io_A_Valid_7_delay_40_21;
    io_A_Valid_7_delay_42_19 <= io_A_Valid_7_delay_41_20;
    io_A_Valid_7_delay_43_18 <= io_A_Valid_7_delay_42_19;
    io_A_Valid_7_delay_44_17 <= io_A_Valid_7_delay_43_18;
    io_A_Valid_7_delay_45_16 <= io_A_Valid_7_delay_44_17;
    io_A_Valid_7_delay_46_15 <= io_A_Valid_7_delay_45_16;
    io_A_Valid_7_delay_47_14 <= io_A_Valid_7_delay_46_15;
    io_A_Valid_7_delay_48_13 <= io_A_Valid_7_delay_47_14;
    io_A_Valid_7_delay_49_12 <= io_A_Valid_7_delay_48_13;
    io_A_Valid_7_delay_50_11 <= io_A_Valid_7_delay_49_12;
    io_A_Valid_7_delay_51_10 <= io_A_Valid_7_delay_50_11;
    io_A_Valid_7_delay_52_9 <= io_A_Valid_7_delay_51_10;
    io_A_Valid_7_delay_53_8 <= io_A_Valid_7_delay_52_9;
    io_A_Valid_7_delay_54_7 <= io_A_Valid_7_delay_53_8;
    io_A_Valid_7_delay_55_6 <= io_A_Valid_7_delay_54_7;
    io_A_Valid_7_delay_56_5 <= io_A_Valid_7_delay_55_6;
    io_A_Valid_7_delay_57_4 <= io_A_Valid_7_delay_56_5;
    io_A_Valid_7_delay_58_3 <= io_A_Valid_7_delay_57_4;
    io_A_Valid_7_delay_59_2 <= io_A_Valid_7_delay_58_3;
    io_A_Valid_7_delay_60_1 <= io_A_Valid_7_delay_59_2;
    io_A_Valid_7_delay_61 <= io_A_Valid_7_delay_60_1;
    io_B_Valid_61_delay_1_6 <= io_B_Valid_61;
    io_B_Valid_61_delay_2_5 <= io_B_Valid_61_delay_1_6;
    io_B_Valid_61_delay_3_4 <= io_B_Valid_61_delay_2_5;
    io_B_Valid_61_delay_4_3 <= io_B_Valid_61_delay_3_4;
    io_B_Valid_61_delay_5_2 <= io_B_Valid_61_delay_4_3;
    io_B_Valid_61_delay_6_1 <= io_B_Valid_61_delay_5_2;
    io_B_Valid_61_delay_7 <= io_B_Valid_61_delay_6_1;
    io_A_Valid_7_delay_1_61 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_60 <= io_A_Valid_7_delay_1_61;
    io_A_Valid_7_delay_3_59 <= io_A_Valid_7_delay_2_60;
    io_A_Valid_7_delay_4_58 <= io_A_Valid_7_delay_3_59;
    io_A_Valid_7_delay_5_57 <= io_A_Valid_7_delay_4_58;
    io_A_Valid_7_delay_6_56 <= io_A_Valid_7_delay_5_57;
    io_A_Valid_7_delay_7_55 <= io_A_Valid_7_delay_6_56;
    io_A_Valid_7_delay_8_54 <= io_A_Valid_7_delay_7_55;
    io_A_Valid_7_delay_9_53 <= io_A_Valid_7_delay_8_54;
    io_A_Valid_7_delay_10_52 <= io_A_Valid_7_delay_9_53;
    io_A_Valid_7_delay_11_51 <= io_A_Valid_7_delay_10_52;
    io_A_Valid_7_delay_12_50 <= io_A_Valid_7_delay_11_51;
    io_A_Valid_7_delay_13_49 <= io_A_Valid_7_delay_12_50;
    io_A_Valid_7_delay_14_48 <= io_A_Valid_7_delay_13_49;
    io_A_Valid_7_delay_15_47 <= io_A_Valid_7_delay_14_48;
    io_A_Valid_7_delay_16_46 <= io_A_Valid_7_delay_15_47;
    io_A_Valid_7_delay_17_45 <= io_A_Valid_7_delay_16_46;
    io_A_Valid_7_delay_18_44 <= io_A_Valid_7_delay_17_45;
    io_A_Valid_7_delay_19_43 <= io_A_Valid_7_delay_18_44;
    io_A_Valid_7_delay_20_42 <= io_A_Valid_7_delay_19_43;
    io_A_Valid_7_delay_21_41 <= io_A_Valid_7_delay_20_42;
    io_A_Valid_7_delay_22_40 <= io_A_Valid_7_delay_21_41;
    io_A_Valid_7_delay_23_39 <= io_A_Valid_7_delay_22_40;
    io_A_Valid_7_delay_24_38 <= io_A_Valid_7_delay_23_39;
    io_A_Valid_7_delay_25_37 <= io_A_Valid_7_delay_24_38;
    io_A_Valid_7_delay_26_36 <= io_A_Valid_7_delay_25_37;
    io_A_Valid_7_delay_27_35 <= io_A_Valid_7_delay_26_36;
    io_A_Valid_7_delay_28_34 <= io_A_Valid_7_delay_27_35;
    io_A_Valid_7_delay_29_33 <= io_A_Valid_7_delay_28_34;
    io_A_Valid_7_delay_30_32 <= io_A_Valid_7_delay_29_33;
    io_A_Valid_7_delay_31_31 <= io_A_Valid_7_delay_30_32;
    io_A_Valid_7_delay_32_30 <= io_A_Valid_7_delay_31_31;
    io_A_Valid_7_delay_33_29 <= io_A_Valid_7_delay_32_30;
    io_A_Valid_7_delay_34_28 <= io_A_Valid_7_delay_33_29;
    io_A_Valid_7_delay_35_27 <= io_A_Valid_7_delay_34_28;
    io_A_Valid_7_delay_36_26 <= io_A_Valid_7_delay_35_27;
    io_A_Valid_7_delay_37_25 <= io_A_Valid_7_delay_36_26;
    io_A_Valid_7_delay_38_24 <= io_A_Valid_7_delay_37_25;
    io_A_Valid_7_delay_39_23 <= io_A_Valid_7_delay_38_24;
    io_A_Valid_7_delay_40_22 <= io_A_Valid_7_delay_39_23;
    io_A_Valid_7_delay_41_21 <= io_A_Valid_7_delay_40_22;
    io_A_Valid_7_delay_42_20 <= io_A_Valid_7_delay_41_21;
    io_A_Valid_7_delay_43_19 <= io_A_Valid_7_delay_42_20;
    io_A_Valid_7_delay_44_18 <= io_A_Valid_7_delay_43_19;
    io_A_Valid_7_delay_45_17 <= io_A_Valid_7_delay_44_18;
    io_A_Valid_7_delay_46_16 <= io_A_Valid_7_delay_45_17;
    io_A_Valid_7_delay_47_15 <= io_A_Valid_7_delay_46_16;
    io_A_Valid_7_delay_48_14 <= io_A_Valid_7_delay_47_15;
    io_A_Valid_7_delay_49_13 <= io_A_Valid_7_delay_48_14;
    io_A_Valid_7_delay_50_12 <= io_A_Valid_7_delay_49_13;
    io_A_Valid_7_delay_51_11 <= io_A_Valid_7_delay_50_12;
    io_A_Valid_7_delay_52_10 <= io_A_Valid_7_delay_51_11;
    io_A_Valid_7_delay_53_9 <= io_A_Valid_7_delay_52_10;
    io_A_Valid_7_delay_54_8 <= io_A_Valid_7_delay_53_9;
    io_A_Valid_7_delay_55_7 <= io_A_Valid_7_delay_54_8;
    io_A_Valid_7_delay_56_6 <= io_A_Valid_7_delay_55_7;
    io_A_Valid_7_delay_57_5 <= io_A_Valid_7_delay_56_6;
    io_A_Valid_7_delay_58_4 <= io_A_Valid_7_delay_57_5;
    io_A_Valid_7_delay_59_3 <= io_A_Valid_7_delay_58_4;
    io_A_Valid_7_delay_60_2 <= io_A_Valid_7_delay_59_3;
    io_A_Valid_7_delay_61_1 <= io_A_Valid_7_delay_60_2;
    io_A_Valid_7_delay_62 <= io_A_Valid_7_delay_61_1;
    io_B_Valid_62_delay_1_6 <= io_B_Valid_62;
    io_B_Valid_62_delay_2_5 <= io_B_Valid_62_delay_1_6;
    io_B_Valid_62_delay_3_4 <= io_B_Valid_62_delay_2_5;
    io_B_Valid_62_delay_4_3 <= io_B_Valid_62_delay_3_4;
    io_B_Valid_62_delay_5_2 <= io_B_Valid_62_delay_4_3;
    io_B_Valid_62_delay_6_1 <= io_B_Valid_62_delay_5_2;
    io_B_Valid_62_delay_7 <= io_B_Valid_62_delay_6_1;
    io_A_Valid_7_delay_1_62 <= io_A_Valid_7;
    io_A_Valid_7_delay_2_61 <= io_A_Valid_7_delay_1_62;
    io_A_Valid_7_delay_3_60 <= io_A_Valid_7_delay_2_61;
    io_A_Valid_7_delay_4_59 <= io_A_Valid_7_delay_3_60;
    io_A_Valid_7_delay_5_58 <= io_A_Valid_7_delay_4_59;
    io_A_Valid_7_delay_6_57 <= io_A_Valid_7_delay_5_58;
    io_A_Valid_7_delay_7_56 <= io_A_Valid_7_delay_6_57;
    io_A_Valid_7_delay_8_55 <= io_A_Valid_7_delay_7_56;
    io_A_Valid_7_delay_9_54 <= io_A_Valid_7_delay_8_55;
    io_A_Valid_7_delay_10_53 <= io_A_Valid_7_delay_9_54;
    io_A_Valid_7_delay_11_52 <= io_A_Valid_7_delay_10_53;
    io_A_Valid_7_delay_12_51 <= io_A_Valid_7_delay_11_52;
    io_A_Valid_7_delay_13_50 <= io_A_Valid_7_delay_12_51;
    io_A_Valid_7_delay_14_49 <= io_A_Valid_7_delay_13_50;
    io_A_Valid_7_delay_15_48 <= io_A_Valid_7_delay_14_49;
    io_A_Valid_7_delay_16_47 <= io_A_Valid_7_delay_15_48;
    io_A_Valid_7_delay_17_46 <= io_A_Valid_7_delay_16_47;
    io_A_Valid_7_delay_18_45 <= io_A_Valid_7_delay_17_46;
    io_A_Valid_7_delay_19_44 <= io_A_Valid_7_delay_18_45;
    io_A_Valid_7_delay_20_43 <= io_A_Valid_7_delay_19_44;
    io_A_Valid_7_delay_21_42 <= io_A_Valid_7_delay_20_43;
    io_A_Valid_7_delay_22_41 <= io_A_Valid_7_delay_21_42;
    io_A_Valid_7_delay_23_40 <= io_A_Valid_7_delay_22_41;
    io_A_Valid_7_delay_24_39 <= io_A_Valid_7_delay_23_40;
    io_A_Valid_7_delay_25_38 <= io_A_Valid_7_delay_24_39;
    io_A_Valid_7_delay_26_37 <= io_A_Valid_7_delay_25_38;
    io_A_Valid_7_delay_27_36 <= io_A_Valid_7_delay_26_37;
    io_A_Valid_7_delay_28_35 <= io_A_Valid_7_delay_27_36;
    io_A_Valid_7_delay_29_34 <= io_A_Valid_7_delay_28_35;
    io_A_Valid_7_delay_30_33 <= io_A_Valid_7_delay_29_34;
    io_A_Valid_7_delay_31_32 <= io_A_Valid_7_delay_30_33;
    io_A_Valid_7_delay_32_31 <= io_A_Valid_7_delay_31_32;
    io_A_Valid_7_delay_33_30 <= io_A_Valid_7_delay_32_31;
    io_A_Valid_7_delay_34_29 <= io_A_Valid_7_delay_33_30;
    io_A_Valid_7_delay_35_28 <= io_A_Valid_7_delay_34_29;
    io_A_Valid_7_delay_36_27 <= io_A_Valid_7_delay_35_28;
    io_A_Valid_7_delay_37_26 <= io_A_Valid_7_delay_36_27;
    io_A_Valid_7_delay_38_25 <= io_A_Valid_7_delay_37_26;
    io_A_Valid_7_delay_39_24 <= io_A_Valid_7_delay_38_25;
    io_A_Valid_7_delay_40_23 <= io_A_Valid_7_delay_39_24;
    io_A_Valid_7_delay_41_22 <= io_A_Valid_7_delay_40_23;
    io_A_Valid_7_delay_42_21 <= io_A_Valid_7_delay_41_22;
    io_A_Valid_7_delay_43_20 <= io_A_Valid_7_delay_42_21;
    io_A_Valid_7_delay_44_19 <= io_A_Valid_7_delay_43_20;
    io_A_Valid_7_delay_45_18 <= io_A_Valid_7_delay_44_19;
    io_A_Valid_7_delay_46_17 <= io_A_Valid_7_delay_45_18;
    io_A_Valid_7_delay_47_16 <= io_A_Valid_7_delay_46_17;
    io_A_Valid_7_delay_48_15 <= io_A_Valid_7_delay_47_16;
    io_A_Valid_7_delay_49_14 <= io_A_Valid_7_delay_48_15;
    io_A_Valid_7_delay_50_13 <= io_A_Valid_7_delay_49_14;
    io_A_Valid_7_delay_51_12 <= io_A_Valid_7_delay_50_13;
    io_A_Valid_7_delay_52_11 <= io_A_Valid_7_delay_51_12;
    io_A_Valid_7_delay_53_10 <= io_A_Valid_7_delay_52_11;
    io_A_Valid_7_delay_54_9 <= io_A_Valid_7_delay_53_10;
    io_A_Valid_7_delay_55_8 <= io_A_Valid_7_delay_54_9;
    io_A_Valid_7_delay_56_7 <= io_A_Valid_7_delay_55_8;
    io_A_Valid_7_delay_57_6 <= io_A_Valid_7_delay_56_7;
    io_A_Valid_7_delay_58_5 <= io_A_Valid_7_delay_57_6;
    io_A_Valid_7_delay_59_4 <= io_A_Valid_7_delay_58_5;
    io_A_Valid_7_delay_60_3 <= io_A_Valid_7_delay_59_4;
    io_A_Valid_7_delay_61_2 <= io_A_Valid_7_delay_60_3;
    io_A_Valid_7_delay_62_1 <= io_A_Valid_7_delay_61_2;
    io_A_Valid_7_delay_63 <= io_A_Valid_7_delay_62_1;
    io_B_Valid_63_delay_1_6 <= io_B_Valid_63;
    io_B_Valid_63_delay_2_5 <= io_B_Valid_63_delay_1_6;
    io_B_Valid_63_delay_3_4 <= io_B_Valid_63_delay_2_5;
    io_B_Valid_63_delay_4_3 <= io_B_Valid_63_delay_3_4;
    io_B_Valid_63_delay_5_2 <= io_B_Valid_63_delay_4_3;
    io_B_Valid_63_delay_6_1 <= io_B_Valid_63_delay_5_2;
    io_B_Valid_63_delay_7 <= io_B_Valid_63_delay_6_1;
  end


endmodule

//AxisDataConverter_7 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

//AxisDataConverter_6 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

//AxisDataConverter_5 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

//AxisDataConverter_4 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

//AxisDataConverter_3 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

//AxisDataConverter_2 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

//AxisDataConverter_1 replaced by AxisDataConverter

//Img2Col_WidthConverter_Fifo replaced by Img2Col_WidthConverter_Fifo

module AxisDataConverter (
  input               inStream_valid,
  output              inStream_ready,
  input      [63:0]   inStream_payload,
  output              outStream_valid,
  input               outStream_ready,
  output     [7:0]    outStream_payload,
  input               clk,
  input               reset
);

  wire       [2:0]    _zz__zz_outStream_payload_1;
  wire       [0:0]    _zz__zz_outStream_payload_1_1;
  wire       [63:0]   _zz__zz_outStream_payload_3;
  reg        [7:0]    _zz_outStream_payload_4;
  wire                outStream_fire;
  reg                 _zz_outStream_payload;
  reg        [2:0]    _zz_outStream_payload_1;
  reg        [2:0]    _zz_outStream_payload_2;
  wire                _zz_inStream_ready;
  wire       [63:0]   _zz_outStream_payload_3;

  assign _zz__zz_outStream_payload_1_1 = _zz_outStream_payload;
  assign _zz__zz_outStream_payload_1 = {2'd0, _zz__zz_outStream_payload_1_1};
  assign _zz__zz_outStream_payload_3 = inStream_payload;
  always @(*) begin
    case(_zz_outStream_payload_2)
      3'b000 : _zz_outStream_payload_4 = _zz_outStream_payload_3[7 : 0];
      3'b001 : _zz_outStream_payload_4 = _zz_outStream_payload_3[15 : 8];
      3'b010 : _zz_outStream_payload_4 = _zz_outStream_payload_3[23 : 16];
      3'b011 : _zz_outStream_payload_4 = _zz_outStream_payload_3[31 : 24];
      3'b100 : _zz_outStream_payload_4 = _zz_outStream_payload_3[39 : 32];
      3'b101 : _zz_outStream_payload_4 = _zz_outStream_payload_3[47 : 40];
      3'b110 : _zz_outStream_payload_4 = _zz_outStream_payload_3[55 : 48];
      default : _zz_outStream_payload_4 = _zz_outStream_payload_3[63 : 56];
    endcase
  end

  assign outStream_fire = (outStream_valid && outStream_ready);
  always @(*) begin
    _zz_outStream_payload = 1'b0;
    if(outStream_fire) begin
      _zz_outStream_payload = 1'b1;
    end
  end

  assign _zz_inStream_ready = (_zz_outStream_payload_2 == 3'b111);
  always @(*) begin
    _zz_outStream_payload_1 = (_zz_outStream_payload_2 + _zz__zz_outStream_payload_1);
    if(1'b0) begin
      _zz_outStream_payload_1 = 3'b000;
    end
  end

  assign outStream_valid = inStream_valid;
  assign _zz_outStream_payload_3 = _zz__zz_outStream_payload_3;
  assign outStream_payload = _zz_outStream_payload_4;
  assign inStream_ready = (outStream_ready && _zz_inStream_ready);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _zz_outStream_payload_2 <= 3'b000;
    end else begin
      _zz_outStream_payload_2 <= _zz_outStream_payload_1;
    end
  end


endmodule

module Img2Col_WidthConverter_Fifo (
  input               io_push_valid,
  output              io_push_ready,
  input      [63:0]   io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [63:0]   io_pop_payload,
  input               io_flush,
  output     [4:0]    io_occupancy,
  output     [4:0]    io_availability,
  input               clk,
  input               reset
);

  reg        [63:0]   _zz_logic_ram_port0;
  wire       [3:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [3:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [63:0]   _zz_logic_ram_port_1;
  wire       [3:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [3:0]    logic_pushPtr_valueNext;
  reg        [3:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [3:0]    logic_popPtr_valueNext;
  reg        [3:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1122;
  wire       [3:0]    logic_ptrDif;
  reg [63:0] logic_ram [0:15];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {3'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {3'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  assign _zz_logic_ram_port_1 = io_push_payload;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 4'b1111);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 4'b0000;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 4'b1111);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 4'b0000;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1122 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_pushPtr_value <= 4'b0000;
      logic_popPtr_value <= 4'b0000;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1122) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module Img2Col_Top (
  input               start,
  input               sData_valid,
  output              sData_ready,
  input      [63:0]   sData_payload,
  output     [63:0]   mData,
  input               mReady,
  output              mValid,
  input               Fifo_Clear,
  output              mLast,
  input      [4:0]    Stride,
  input      [4:0]    Kernel_Size,
  input      [15:0]   Window_Size,
  input      [15:0]   InFeature_Size,
  input      [15:0]   InFeature_Channel,
  input      [15:0]   OutFeature_Channel,
  input      [15:0]   OutFeature_Size,
  input      [15:0]   OutCol_Count_Times,
  input      [15:0]   InCol_Count_Times,
  input      [15:0]   OutRow_Count_Times,
  input      [15:0]   OutFeature_Channel_Count_Times,
  input      [12:0]   Sliding_Size,
  output              Test_Signal,
  input      [15:0]   Test_Generate_Period,
  output              Test_End,
  output              Raddr_Valid,
  output              LayerEnd,
  output              SA_Row_Cnt_Valid,
  input               clk,
  input               reset
);
  localparam IMG2COL_ENUM_IDLE = 7'd1;
  localparam IMG2COL_ENUM_INIT = 7'd2;
  localparam IMG2COL_ENUM_INIT_ADDR = 7'd4;
  localparam IMG2COL_ENUM_DATA_CACHE = 7'd8;
  localparam IMG2COL_ENUM_WAIT_COMPUTE = 7'd16;
  localparam IMG2COL_ENUM_UPDATE_ADDR = 7'd32;
  localparam IMG2COL_ENUM_START_COMPUTE = 7'd64;

  reg                 AddrFifo_io_push_valid;
  reg                 AddrFifo_io_pop_ready;
  wire                AddrFifo_io_flush;
  reg                 RaddrFifo0_io_push_valid;
  reg        [15:0]   RaddrFifo0_io_push_payload;
  reg                 RaddrFifo0_io_pop_ready;
  wire                RaddrFifo0_io_flush;
  wire                Img2Col_SubModule_start;
  wire                Img2Col_SubModule_NewAddrIn_valid;
  wire       [13:0]   DGB_addra;
  wire       [13:0]   DGB_addrb;
  wire                AddrFifo_io_push_ready;
  wire                AddrFifo_io_pop_valid;
  wire       [15:0]   AddrFifo_io_pop_payload;
  wire       [5:0]    AddrFifo_io_occupancy;
  wire       [5:0]    AddrFifo_io_availability;
  wire                RaddrFifo0_io_push_ready;
  wire                RaddrFifo0_io_pop_valid;
  wire       [15:0]   RaddrFifo0_io_pop_payload;
  wire       [5:0]    RaddrFifo0_io_occupancy;
  wire       [5:0]    RaddrFifo0_io_availability;
  wire                Img2Col_SubModule_NewAddrIn_ready;
  wire                Img2Col_SubModule_SA_Idle;
  wire       [15:0]   Img2Col_SubModule_Raddr;
  wire                Img2Col_SubModule_Raddr_Valid;
  wire                Img2Col_SubModule_SA_End;
  wire                Img2Col_SubModule_AddrReceived;
  wire                Img2Col_SubModule_SA_Row_Cnt_Valid;
  wire       [63:0]   DGB_doutb;
  wire       [4:0]    _zz_Addr_Init_Cnt_valid;
  wire       [4:0]    _zz_Addr_Init_Cnt_valid_1;
  wire       [15:0]   _zz_In_Col_Cnt_valid;
  wire       [4:0]    _zz_Row_Cache_Cnt_valid;
  wire       [15:0]   _zz_In_Row_Cnt_valid;
  wire       [15:0]   _zz_when_Data_Generate_V2_l217;
  wire       [4:0]    _zz_when_Data_Generate_V2_l217_1;
  wire       [15:0]   _zz_Out_Row_Cnt_valid;
  wire       [15:0]   _zz_Test_Valid;
  reg                 start_regNext;
  wire                when_Data_Generate_V2_l59;
  reg        [6:0]    Fsm_currentState;
  reg        [6:0]    Fsm_nextState;
  wire                Fsm_Init_End;
  wire                Fsm_Addr_Inited;
  wire                Fsm_Data_Cached;
  wire                Fsm_Addr_Updated;
  wire                Fsm_SA_Ready;
  wire                Fsm_Cache_End;
  wire                Fsm_Layer_End;
  wire                when_WaCounter_l19;
  reg        [2:0]    Init_Count_count;
  reg                 Init_Count_valid;
  wire                when_WaCounter_l14;
  wire                when_WaCounter_l40;
  reg        [4:0]    Addr_Init_Cnt_count;
  wire                Addr_Init_Cnt_valid;
  reg        [15:0]   WaddrOffset;
  wire                when_Data_Generate_V2_l170;
  wire                when_Data_Generate_V2_l175;
  wire                SubModule_AddrFifo_io_pop_fire;
  wire                when_Data_Generate_V2_l179;
  wire                when_Data_Generate_V2_l183;
  reg        [15:0]   Raddr_Initialization;
  wire                when_Data_Generate_V2_l193;
  wire                when_Data_Generate_V2_l197;
  reg        [4:0]    Cache_Row_Num;
  reg        [4:0]    Raddr_Updata_Cnt_Num;
  wire                sData_fire;
  reg        [15:0]   In_Col_Cnt_count;
  wire                In_Col_Cnt_valid;
  reg        [4:0]    Row_Cache_Cnt_count;
  wire                Row_Cache_Cnt_valid;
  reg        [15:0]   In_Row_Cnt_count;
  wire                In_Row_Cnt_valid;
  wire                when_Data_Generate_V2_l217;
  reg                 CacheEnd_Flag;
  wire                when_Data_Generate_V2_l228;
  wire                Img2ColOutput_Module_Ready_Receive_Addr;
  wire                when_Data_Generate_V2_l245;
  wire                SubModule_RaddrFifo0_io_pop_fire;
  reg        [15:0]   Out_Row_Cnt_count;
  wire                Out_Row_Cnt_valid;
  wire       [15:0]   Waddr;
  wire                sData_fire_1;
  reg                 SubModule_Img2Col_SubModule_Raddr_Valid_regNext;
  reg                 Out_Row_Cnt_valid_regNext;
  reg        [15:0]   Out_Row_Cnt_count_regNext;
  wire                Test_Valid;
  reg                 Test_Valid_regNext;
  `ifndef SYNTHESIS
  reg [103:0] Fsm_currentState_string;
  reg [103:0] Fsm_nextState_string;
  `endif


  assign _zz_Addr_Init_Cnt_valid = (_zz_Addr_Init_Cnt_valid_1 - 5'h01);
  assign _zz_Addr_Init_Cnt_valid_1 = (Kernel_Size + Stride);
  assign _zz_In_Col_Cnt_valid = (InCol_Count_Times - 16'h0001);
  assign _zz_Row_Cache_Cnt_valid = (Cache_Row_Num - 5'h01);
  assign _zz_In_Row_Cnt_valid = (InFeature_Size - 16'h0001);
  assign _zz_when_Data_Generate_V2_l217_1 = (Kernel_Size - 5'h01);
  assign _zz_when_Data_Generate_V2_l217 = {11'd0, _zz_when_Data_Generate_V2_l217_1};
  assign _zz_Out_Row_Cnt_valid = (OutRow_Count_Times - 16'h0001);
  assign _zz_Test_Valid = (Test_Generate_Period - 16'h0001);
  WaddrOffset_Fifo_2 AddrFifo (
    .io_push_valid   (AddrFifo_io_push_valid       ), //i
    .io_push_ready   (AddrFifo_io_push_ready       ), //o
    .io_push_payload (WaddrOffset[15:0]            ), //i
    .io_pop_valid    (AddrFifo_io_pop_valid        ), //o
    .io_pop_ready    (AddrFifo_io_pop_ready        ), //i
    .io_pop_payload  (AddrFifo_io_pop_payload[15:0]), //o
    .io_flush        (AddrFifo_io_flush            ), //i
    .io_occupancy    (AddrFifo_io_occupancy[5:0]   ), //o
    .io_availability (AddrFifo_io_availability[5:0]), //o
    .clk             (clk                          ), //i
    .reset           (reset                        )  //i
  );
  WaddrOffset_Fifo_2 RaddrFifo0 (
    .io_push_valid   (RaddrFifo0_io_push_valid        ), //i
    .io_push_ready   (RaddrFifo0_io_push_ready        ), //o
    .io_push_payload (RaddrFifo0_io_push_payload[15:0]), //i
    .io_pop_valid    (RaddrFifo0_io_pop_valid         ), //o
    .io_pop_ready    (RaddrFifo0_io_pop_ready         ), //i
    .io_pop_payload  (RaddrFifo0_io_pop_payload[15:0] ), //o
    .io_flush        (RaddrFifo0_io_flush             ), //i
    .io_occupancy    (RaddrFifo0_io_occupancy[5:0]    ), //o
    .io_availability (RaddrFifo0_io_availability[5:0] ), //o
    .clk             (clk                             ), //i
    .reset           (reset                           )  //i
  );
  Img2Col_OutPut Img2Col_SubModule (
    .start                          (Img2Col_SubModule_start             ), //i
    .NewAddrIn_valid                (Img2Col_SubModule_NewAddrIn_valid   ), //i
    .NewAddrIn_ready                (Img2Col_SubModule_NewAddrIn_ready   ), //o
    .NewAddrIn_payload              (RaddrFifo0_io_pop_payload[15:0]     ), //i
    .SA_Idle                        (Img2Col_SubModule_SA_Idle           ), //o
    .Raddr                          (Img2Col_SubModule_Raddr[15:0]       ), //o
    .Raddr_Valid                    (Img2Col_SubModule_Raddr_Valid       ), //o
    .SA_End                         (Img2Col_SubModule_SA_End            ), //o
    .Stride                         (Stride[4:0]                         ), //i
    .Kernel_Size                    (Kernel_Size[4:0]                    ), //i
    .Window_Size                    (Window_Size[15:0]                   ), //i
    .InFeature_Size                 (InFeature_Size[15:0]                ), //i
    .InFeature_Channel              (InFeature_Channel[15:0]             ), //i
    .OutFeature_Channel             (OutFeature_Channel[15:0]            ), //i
    .OutFeature_Size                (OutFeature_Size[15:0]               ), //i
    .OutCol_Count_Times             (OutCol_Count_Times[15:0]            ), //i
    .InCol_Count_Times              (InCol_Count_Times[15:0]             ), //i
    .OutFeature_Channel_Count_Times (OutFeature_Channel_Count_Times[15:0]), //i
    .Sliding_Size                   (Sliding_Size[12:0]                  ), //i
    .mReady                         (mReady                              ), //i
    .Fifo_Clear                     (Fifo_Clear                          ), //i
    .AddrReceived                   (Img2Col_SubModule_AddrReceived      ), //o
    .LayerEnd                       (Fsm_Layer_End                       ), //i
    .SA_Row_Cnt_Valid               (Img2Col_SubModule_SA_Row_Cnt_Valid  ), //o
    .clk                            (clk                                 ), //i
    .reset                          (reset                               )  //i
  );
  DataGen_Bram DGB (
    .clka  (clk                ), //i
    .addra (DGB_addra[13:0]    ), //i
    .dina  (sData_payload[63:0]), //i
    .ena   (sData_fire_1       ), //i
    .wea   (1'b1               ), //i
    .addrb (DGB_addrb[13:0]    ), //i
    .doutb (DGB_doutb[63:0]    ), //o
    .clkb  (clk                )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      IMG2COL_ENUM_IDLE : Fsm_currentState_string = "IDLE         ";
      IMG2COL_ENUM_INIT : Fsm_currentState_string = "INIT         ";
      IMG2COL_ENUM_INIT_ADDR : Fsm_currentState_string = "INIT_ADDR    ";
      IMG2COL_ENUM_DATA_CACHE : Fsm_currentState_string = "DATA_CACHE   ";
      IMG2COL_ENUM_WAIT_COMPUTE : Fsm_currentState_string = "WAIT_COMPUTE ";
      IMG2COL_ENUM_UPDATE_ADDR : Fsm_currentState_string = "UPDATE_ADDR  ";
      IMG2COL_ENUM_START_COMPUTE : Fsm_currentState_string = "START_COMPUTE";
      default : Fsm_currentState_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      IMG2COL_ENUM_IDLE : Fsm_nextState_string = "IDLE         ";
      IMG2COL_ENUM_INIT : Fsm_nextState_string = "INIT         ";
      IMG2COL_ENUM_INIT_ADDR : Fsm_nextState_string = "INIT_ADDR    ";
      IMG2COL_ENUM_DATA_CACHE : Fsm_nextState_string = "DATA_CACHE   ";
      IMG2COL_ENUM_WAIT_COMPUTE : Fsm_nextState_string = "WAIT_COMPUTE ";
      IMG2COL_ENUM_UPDATE_ADDR : Fsm_nextState_string = "UPDATE_ADDR  ";
      IMG2COL_ENUM_START_COMPUTE : Fsm_nextState_string = "START_COMPUTE";
      default : Fsm_nextState_string = "?????????????";
    endcase
  end
  `endif

  assign when_Data_Generate_V2_l59 = (start && (! start_regNext));
  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & IMG2COL_ENUM_IDLE) == IMG2COL_ENUM_IDLE) : begin
        if(when_Data_Generate_V2_l59) begin
          Fsm_nextState = IMG2COL_ENUM_INIT;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_IDLE;
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_INIT) == IMG2COL_ENUM_INIT) : begin
        if(Fsm_Init_End) begin
          Fsm_nextState = IMG2COL_ENUM_INIT_ADDR;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_INIT;
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_INIT_ADDR) == IMG2COL_ENUM_INIT_ADDR) : begin
        if(Fsm_Addr_Inited) begin
          Fsm_nextState = IMG2COL_ENUM_DATA_CACHE;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_INIT_ADDR;
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_DATA_CACHE) == IMG2COL_ENUM_DATA_CACHE) : begin
        if(Fsm_Data_Cached) begin
          Fsm_nextState = IMG2COL_ENUM_WAIT_COMPUTE;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_DATA_CACHE;
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_WAIT_COMPUTE) == IMG2COL_ENUM_WAIT_COMPUTE) : begin
        if(Fsm_Layer_End) begin
          Fsm_nextState = IMG2COL_ENUM_IDLE;
        end else begin
          if(Fsm_SA_Ready) begin
            Fsm_nextState = IMG2COL_ENUM_UPDATE_ADDR;
          end else begin
            Fsm_nextState = IMG2COL_ENUM_WAIT_COMPUTE;
          end
        end
      end
      (((Fsm_currentState) & IMG2COL_ENUM_UPDATE_ADDR) == IMG2COL_ENUM_UPDATE_ADDR) : begin
        if(Fsm_Addr_Updated) begin
          Fsm_nextState = IMG2COL_ENUM_START_COMPUTE;
        end else begin
          Fsm_nextState = IMG2COL_ENUM_UPDATE_ADDR;
        end
      end
      default : begin
        if(Fsm_Layer_End) begin
          Fsm_nextState = IMG2COL_ENUM_IDLE;
        end else begin
          if(Fsm_Cache_End) begin
            Fsm_nextState = IMG2COL_ENUM_WAIT_COMPUTE;
          end else begin
            Fsm_nextState = IMG2COL_ENUM_DATA_CACHE;
          end
        end
      end
    endcase
  end

  assign when_WaCounter_l19 = ((Fsm_currentState & IMG2COL_ENUM_INIT) != 7'b0000000);
  assign when_WaCounter_l14 = (Init_Count_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l14) begin
      Init_Count_valid = 1'b1;
    end else begin
      Init_Count_valid = 1'b0;
    end
  end

  assign Fsm_Init_End = Init_Count_valid;
  assign when_WaCounter_l40 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign Addr_Init_Cnt_valid = ((Addr_Init_Cnt_count == _zz_Addr_Init_Cnt_valid) && when_WaCounter_l40);
  assign Fsm_Addr_Inited = Addr_Init_Cnt_valid;
  always @(*) begin
    AddrFifo_io_push_valid = 1'b0;
    if(when_Data_Generate_V2_l170) begin
      AddrFifo_io_push_valid = 1'b1;
    end
    if(In_Col_Cnt_valid) begin
      AddrFifo_io_push_valid = 1'b1;
    end
  end

  always @(*) begin
    AddrFifo_io_pop_ready = 1'b0;
    if(when_Data_Generate_V2_l183) begin
      AddrFifo_io_pop_ready = 1'b1;
    end
    if(In_Col_Cnt_valid) begin
      AddrFifo_io_pop_ready = 1'b1;
    end
  end

  assign when_Data_Generate_V2_l170 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign when_Data_Generate_V2_l175 = ((Fsm_currentState & IMG2COL_ENUM_INIT) != 7'b0000000);
  assign SubModule_AddrFifo_io_pop_fire = (AddrFifo_io_pop_valid && AddrFifo_io_pop_ready);
  assign when_Data_Generate_V2_l179 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign when_Data_Generate_V2_l183 = (((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000) && ((Fsm_nextState & IMG2COL_ENUM_DATA_CACHE) != 7'b0000000));
  always @(*) begin
    RaddrFifo0_io_push_valid = 1'b0;
    if(when_Data_Generate_V2_l193) begin
      RaddrFifo0_io_push_valid = 1'b1;
    end
    if(when_Data_Generate_V2_l245) begin
      RaddrFifo0_io_push_valid = SubModule_RaddrFifo0_io_pop_fire;
    end
  end

  always @(*) begin
    RaddrFifo0_io_pop_ready = 1'b0;
    if(when_Data_Generate_V2_l245) begin
      RaddrFifo0_io_pop_ready = Img2ColOutput_Module_Ready_Receive_Addr;
    end
  end

  always @(*) begin
    RaddrFifo0_io_push_payload = RaddrFifo0_io_pop_payload;
    if(when_Data_Generate_V2_l193) begin
      RaddrFifo0_io_push_payload = Raddr_Initialization;
    end
    if(when_Data_Generate_V2_l245) begin
      RaddrFifo0_io_push_payload = RaddrFifo0_io_pop_payload;
    end
  end

  assign when_Data_Generate_V2_l193 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign when_Data_Generate_V2_l197 = ((Fsm_currentState & IMG2COL_ENUM_INIT_ADDR) != 7'b0000000);
  assign sData_fire = (sData_valid && sData_ready);
  assign In_Col_Cnt_valid = ((In_Col_Cnt_count == _zz_In_Col_Cnt_valid) && sData_fire);
  assign Row_Cache_Cnt_valid = ((Row_Cache_Cnt_count == _zz_Row_Cache_Cnt_valid) && In_Col_Cnt_valid);
  assign In_Row_Cnt_valid = ((In_Row_Cnt_count == _zz_In_Row_Cnt_valid) && In_Col_Cnt_valid);
  assign when_Data_Generate_V2_l217 = (_zz_when_Data_Generate_V2_l217 < In_Row_Cnt_count);
  always @(*) begin
    if(when_Data_Generate_V2_l217) begin
      Cache_Row_Num = Stride;
    end else begin
      Cache_Row_Num = Kernel_Size;
    end
  end

  always @(*) begin
    if(when_Data_Generate_V2_l217) begin
      Raddr_Updata_Cnt_Num = Stride;
    end else begin
      Raddr_Updata_Cnt_Num = Kernel_Size;
    end
  end

  assign Fsm_Data_Cached = Row_Cache_Cnt_valid;
  assign when_Data_Generate_V2_l228 = ((Fsm_currentState & IMG2COL_ENUM_IDLE) != 7'b0000000);
  assign Fsm_Cache_End = CacheEnd_Flag;
  assign sData_ready = ((Fsm_currentState & IMG2COL_ENUM_DATA_CACHE) != 7'b0000000);
  assign when_Data_Generate_V2_l245 = ((Fsm_currentState & IMG2COL_ENUM_UPDATE_ADDR) != 7'b0000000);
  assign SubModule_RaddrFifo0_io_pop_fire = (RaddrFifo0_io_pop_valid && RaddrFifo0_io_pop_ready);
  assign Img2Col_SubModule_start = ((Fsm_currentState & IMG2COL_ENUM_UPDATE_ADDR) != 7'b0000000);
  assign Fsm_SA_Ready = Img2Col_SubModule_SA_Idle;
  assign Img2ColOutput_Module_Ready_Receive_Addr = Img2Col_SubModule_NewAddrIn_ready;
  assign Img2Col_SubModule_NewAddrIn_valid = ((Fsm_currentState & IMG2COL_ENUM_UPDATE_ADDR) != 7'b0000000);
  assign SA_Row_Cnt_Valid = Img2Col_SubModule_SA_Row_Cnt_Valid;
  assign LayerEnd = Fsm_Layer_End;
  assign Fsm_Addr_Updated = Img2Col_SubModule_AddrReceived;
  assign Out_Row_Cnt_valid = ((Out_Row_Cnt_count == _zz_Out_Row_Cnt_valid) && Img2Col_SubModule_SA_End);
  assign Fsm_Layer_End = Out_Row_Cnt_valid;
  assign Waddr = (WaddrOffset + In_Col_Cnt_count);
  assign DGB_addra = Waddr[13:0];
  assign sData_fire_1 = (sData_valid && sData_ready);
  assign DGB_addrb = Img2Col_SubModule_Raddr[13:0];
  assign mData = DGB_doutb;
  assign mValid = SubModule_Img2Col_SubModule_Raddr_Valid_regNext;
  assign mLast = Out_Row_Cnt_valid_regNext;
  assign Test_Valid = (_zz_Test_Valid == Out_Row_Cnt_count_regNext);
  assign Test_Signal = Test_Valid;
  assign Test_End = ((! Test_Valid) && Test_Valid_regNext);
  assign AddrFifo_io_flush = ((Fsm_nextState & IMG2COL_ENUM_IDLE) != 7'b0000000);
  assign RaddrFifo0_io_flush = ((Fsm_nextState & IMG2COL_ENUM_IDLE) != 7'b0000000);
  assign Raddr_Valid = Img2Col_SubModule_Raddr_Valid;
  always @(posedge clk) begin
    start_regNext <= start;
    SubModule_Img2Col_SubModule_Raddr_Valid_regNext <= Img2Col_SubModule_Raddr_Valid;
    Out_Row_Cnt_valid_regNext <= Out_Row_Cnt_valid;
    Out_Row_Cnt_count_regNext <= Out_Row_Cnt_count;
    Test_Valid_regNext <= Test_Valid;
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= IMG2COL_ENUM_IDLE;
      Init_Count_count <= 3'b000;
      Addr_Init_Cnt_count <= 5'h0;
      WaddrOffset <= 16'h0;
      Raddr_Initialization <= 16'h0;
      In_Col_Cnt_count <= 16'h0;
      Row_Cache_Cnt_count <= 5'h0;
      In_Row_Cnt_count <= 16'h0;
      CacheEnd_Flag <= 1'b0;
      Out_Row_Cnt_count <= 16'h0;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l19) begin
        Init_Count_count <= (Init_Count_count + 3'b001);
        if(Init_Count_valid) begin
          Init_Count_count <= 3'b000;
        end
      end
      if(when_WaCounter_l40) begin
        if(Addr_Init_Cnt_valid) begin
          Addr_Init_Cnt_count <= 5'h0;
        end else begin
          Addr_Init_Cnt_count <= (Addr_Init_Cnt_count + 5'h01);
        end
      end
      if(when_Data_Generate_V2_l175) begin
        WaddrOffset <= 16'h0;
      end else begin
        if(SubModule_AddrFifo_io_pop_fire) begin
          WaddrOffset <= AddrFifo_io_pop_payload;
        end else begin
          if(when_Data_Generate_V2_l179) begin
            WaddrOffset <= (WaddrOffset + InCol_Count_Times);
          end
        end
      end
      if(when_Data_Generate_V2_l197) begin
        Raddr_Initialization <= (Raddr_Initialization + InCol_Count_Times);
      end else begin
        Raddr_Initialization <= 16'h0;
      end
      if(sData_fire) begin
        if(In_Col_Cnt_valid) begin
          In_Col_Cnt_count <= 16'h0;
        end else begin
          In_Col_Cnt_count <= (In_Col_Cnt_count + 16'h0001);
        end
      end
      if(In_Col_Cnt_valid) begin
        if(Row_Cache_Cnt_valid) begin
          Row_Cache_Cnt_count <= 5'h0;
        end else begin
          Row_Cache_Cnt_count <= (Row_Cache_Cnt_count + 5'h01);
        end
      end
      if(In_Col_Cnt_valid) begin
        if(In_Row_Cnt_valid) begin
          In_Row_Cnt_count <= 16'h0;
        end else begin
          In_Row_Cnt_count <= (In_Row_Cnt_count + 16'h0001);
        end
      end
      if(In_Row_Cnt_valid) begin
        CacheEnd_Flag <= 1'b1;
      end else begin
        if(when_Data_Generate_V2_l228) begin
          CacheEnd_Flag <= 1'b0;
        end
      end
      if(Img2Col_SubModule_SA_End) begin
        if(Out_Row_Cnt_valid) begin
          Out_Row_Cnt_count <= 16'h0;
        end else begin
          Out_Row_Cnt_count <= (Out_Row_Cnt_count + 16'h0001);
        end
      end
    end
  end


endmodule

//PE_511 replaced by PE

//PE_510 replaced by PE

//PE_509 replaced by PE

//PE_508 replaced by PE

//PE_507 replaced by PE

//PE_506 replaced by PE

//PE_505 replaced by PE

//PE_504 replaced by PE

//PE_503 replaced by PE

//PE_502 replaced by PE

//PE_501 replaced by PE

//PE_500 replaced by PE

//PE_499 replaced by PE

//PE_498 replaced by PE

//PE_497 replaced by PE

//PE_496 replaced by PE

//PE_495 replaced by PE

//PE_494 replaced by PE

//PE_493 replaced by PE

//PE_492 replaced by PE

//PE_491 replaced by PE

//PE_490 replaced by PE

//PE_489 replaced by PE

//PE_488 replaced by PE

//PE_487 replaced by PE

//PE_486 replaced by PE

//PE_485 replaced by PE

//PE_484 replaced by PE

//PE_483 replaced by PE

//PE_482 replaced by PE

//PE_481 replaced by PE

//PE_480 replaced by PE

//PE_479 replaced by PE

//PE_478 replaced by PE

//PE_477 replaced by PE

//PE_476 replaced by PE

//PE_475 replaced by PE

//PE_474 replaced by PE

//PE_473 replaced by PE

//PE_472 replaced by PE

//PE_471 replaced by PE

//PE_470 replaced by PE

//PE_469 replaced by PE

//PE_468 replaced by PE

//PE_467 replaced by PE

//PE_466 replaced by PE

//PE_465 replaced by PE

//PE_464 replaced by PE

//PE_463 replaced by PE

//PE_462 replaced by PE

//PE_461 replaced by PE

//PE_460 replaced by PE

//PE_459 replaced by PE

//PE_458 replaced by PE

//PE_457 replaced by PE

//PE_456 replaced by PE

//PE_455 replaced by PE

//PE_454 replaced by PE

//PE_453 replaced by PE

//PE_452 replaced by PE

//PE_451 replaced by PE

//PE_450 replaced by PE

//PE_449 replaced by PE

//PE_448 replaced by PE

//PE_447 replaced by PE

//PE_446 replaced by PE

//PE_445 replaced by PE

//PE_444 replaced by PE

//PE_443 replaced by PE

//PE_442 replaced by PE

//PE_441 replaced by PE

//PE_440 replaced by PE

//PE_439 replaced by PE

//PE_438 replaced by PE

//PE_437 replaced by PE

//PE_436 replaced by PE

//PE_435 replaced by PE

//PE_434 replaced by PE

//PE_433 replaced by PE

//PE_432 replaced by PE

//PE_431 replaced by PE

//PE_430 replaced by PE

//PE_429 replaced by PE

//PE_428 replaced by PE

//PE_427 replaced by PE

//PE_426 replaced by PE

//PE_425 replaced by PE

//PE_424 replaced by PE

//PE_423 replaced by PE

//PE_422 replaced by PE

//PE_421 replaced by PE

//PE_420 replaced by PE

//PE_419 replaced by PE

//PE_418 replaced by PE

//PE_417 replaced by PE

//PE_416 replaced by PE

//PE_415 replaced by PE

//PE_414 replaced by PE

//PE_413 replaced by PE

//PE_412 replaced by PE

//PE_411 replaced by PE

//PE_410 replaced by PE

//PE_409 replaced by PE

//PE_408 replaced by PE

//PE_407 replaced by PE

//PE_406 replaced by PE

//PE_405 replaced by PE

//PE_404 replaced by PE

//PE_403 replaced by PE

//PE_402 replaced by PE

//PE_401 replaced by PE

//PE_400 replaced by PE

//PE_399 replaced by PE

//PE_398 replaced by PE

//PE_397 replaced by PE

//PE_396 replaced by PE

//PE_395 replaced by PE

//PE_394 replaced by PE

//PE_393 replaced by PE

//PE_392 replaced by PE

//PE_391 replaced by PE

//PE_390 replaced by PE

//PE_389 replaced by PE

//PE_388 replaced by PE

//PE_387 replaced by PE

//PE_386 replaced by PE

//PE_385 replaced by PE

//PE_384 replaced by PE

//PE_383 replaced by PE

//PE_382 replaced by PE

//PE_381 replaced by PE

//PE_380 replaced by PE

//PE_379 replaced by PE

//PE_378 replaced by PE

//PE_377 replaced by PE

//PE_376 replaced by PE

//PE_375 replaced by PE

//PE_374 replaced by PE

//PE_373 replaced by PE

//PE_372 replaced by PE

//PE_371 replaced by PE

//PE_370 replaced by PE

//PE_369 replaced by PE

//PE_368 replaced by PE

//PE_367 replaced by PE

//PE_366 replaced by PE

//PE_365 replaced by PE

//PE_364 replaced by PE

//PE_363 replaced by PE

//PE_362 replaced by PE

//PE_361 replaced by PE

//PE_360 replaced by PE

//PE_359 replaced by PE

//PE_358 replaced by PE

//PE_357 replaced by PE

//PE_356 replaced by PE

//PE_355 replaced by PE

//PE_354 replaced by PE

//PE_353 replaced by PE

//PE_352 replaced by PE

//PE_351 replaced by PE

//PE_350 replaced by PE

//PE_349 replaced by PE

//PE_348 replaced by PE

//PE_347 replaced by PE

//PE_346 replaced by PE

//PE_345 replaced by PE

//PE_344 replaced by PE

//PE_343 replaced by PE

//PE_342 replaced by PE

//PE_341 replaced by PE

//PE_340 replaced by PE

//PE_339 replaced by PE

//PE_338 replaced by PE

//PE_337 replaced by PE

//PE_336 replaced by PE

//PE_335 replaced by PE

//PE_334 replaced by PE

//PE_333 replaced by PE

//PE_332 replaced by PE

//PE_331 replaced by PE

//PE_330 replaced by PE

//PE_329 replaced by PE

//PE_328 replaced by PE

//PE_327 replaced by PE

//PE_326 replaced by PE

//PE_325 replaced by PE

//PE_324 replaced by PE

//PE_323 replaced by PE

//PE_322 replaced by PE

//PE_321 replaced by PE

//PE_320 replaced by PE

//PE_319 replaced by PE

//PE_318 replaced by PE

//PE_317 replaced by PE

//PE_316 replaced by PE

//PE_315 replaced by PE

//PE_314 replaced by PE

//PE_313 replaced by PE

//PE_312 replaced by PE

//PE_311 replaced by PE

//PE_310 replaced by PE

//PE_309 replaced by PE

//PE_308 replaced by PE

//PE_307 replaced by PE

//PE_306 replaced by PE

//PE_305 replaced by PE

//PE_304 replaced by PE

//PE_303 replaced by PE

//PE_302 replaced by PE

//PE_301 replaced by PE

//PE_300 replaced by PE

//PE_299 replaced by PE

//PE_298 replaced by PE

//PE_297 replaced by PE

//PE_296 replaced by PE

//PE_295 replaced by PE

//PE_294 replaced by PE

//PE_293 replaced by PE

//PE_292 replaced by PE

//PE_291 replaced by PE

//PE_290 replaced by PE

//PE_289 replaced by PE

//PE_288 replaced by PE

//PE_287 replaced by PE

//PE_286 replaced by PE

//PE_285 replaced by PE

//PE_284 replaced by PE

//PE_283 replaced by PE

//PE_282 replaced by PE

//PE_281 replaced by PE

//PE_280 replaced by PE

//PE_279 replaced by PE

//PE_278 replaced by PE

//PE_277 replaced by PE

//PE_276 replaced by PE

//PE_275 replaced by PE

//PE_274 replaced by PE

//PE_273 replaced by PE

//PE_272 replaced by PE

//PE_271 replaced by PE

//PE_270 replaced by PE

//PE_269 replaced by PE

//PE_268 replaced by PE

//PE_267 replaced by PE

//PE_266 replaced by PE

//PE_265 replaced by PE

//PE_264 replaced by PE

//PE_263 replaced by PE

//PE_262 replaced by PE

//PE_261 replaced by PE

//PE_260 replaced by PE

//PE_259 replaced by PE

//PE_258 replaced by PE

//PE_257 replaced by PE

//PE_256 replaced by PE

//PE_255 replaced by PE

//PE_254 replaced by PE

//PE_253 replaced by PE

//PE_252 replaced by PE

//PE_251 replaced by PE

//PE_250 replaced by PE

//PE_249 replaced by PE

//PE_248 replaced by PE

//PE_247 replaced by PE

//PE_246 replaced by PE

//PE_245 replaced by PE

//PE_244 replaced by PE

//PE_243 replaced by PE

//PE_242 replaced by PE

//PE_241 replaced by PE

//PE_240 replaced by PE

//PE_239 replaced by PE

//PE_238 replaced by PE

//PE_237 replaced by PE

//PE_236 replaced by PE

//PE_235 replaced by PE

//PE_234 replaced by PE

//PE_233 replaced by PE

//PE_232 replaced by PE

//PE_231 replaced by PE

//PE_230 replaced by PE

//PE_229 replaced by PE

//PE_228 replaced by PE

//PE_227 replaced by PE

//PE_226 replaced by PE

//PE_225 replaced by PE

//PE_224 replaced by PE

//PE_223 replaced by PE

//PE_222 replaced by PE

//PE_221 replaced by PE

//PE_220 replaced by PE

//PE_219 replaced by PE

//PE_218 replaced by PE

//PE_217 replaced by PE

//PE_216 replaced by PE

//PE_215 replaced by PE

//PE_214 replaced by PE

//PE_213 replaced by PE

//PE_212 replaced by PE

//PE_211 replaced by PE

//PE_210 replaced by PE

//PE_209 replaced by PE

//PE_208 replaced by PE

//PE_207 replaced by PE

//PE_206 replaced by PE

//PE_205 replaced by PE

//PE_204 replaced by PE

//PE_203 replaced by PE

//PE_202 replaced by PE

//PE_201 replaced by PE

//PE_200 replaced by PE

//PE_199 replaced by PE

//PE_198 replaced by PE

//PE_197 replaced by PE

//PE_196 replaced by PE

//PE_195 replaced by PE

//PE_194 replaced by PE

//PE_193 replaced by PE

//PE_192 replaced by PE

//PE_191 replaced by PE

//PE_190 replaced by PE

//PE_189 replaced by PE

//PE_188 replaced by PE

//PE_187 replaced by PE

//PE_186 replaced by PE

//PE_185 replaced by PE

//PE_184 replaced by PE

//PE_183 replaced by PE

//PE_182 replaced by PE

//PE_181 replaced by PE

//PE_180 replaced by PE

//PE_179 replaced by PE

//PE_178 replaced by PE

//PE_177 replaced by PE

//PE_176 replaced by PE

//PE_175 replaced by PE

//PE_174 replaced by PE

//PE_173 replaced by PE

//PE_172 replaced by PE

//PE_171 replaced by PE

//PE_170 replaced by PE

//PE_169 replaced by PE

//PE_168 replaced by PE

//PE_167 replaced by PE

//PE_166 replaced by PE

//PE_165 replaced by PE

//PE_164 replaced by PE

//PE_163 replaced by PE

//PE_162 replaced by PE

//PE_161 replaced by PE

//PE_160 replaced by PE

//PE_159 replaced by PE

//PE_158 replaced by PE

//PE_157 replaced by PE

//PE_156 replaced by PE

//PE_155 replaced by PE

//PE_154 replaced by PE

//PE_153 replaced by PE

//PE_152 replaced by PE

//PE_151 replaced by PE

//PE_150 replaced by PE

//PE_149 replaced by PE

//PE_148 replaced by PE

//PE_147 replaced by PE

//PE_146 replaced by PE

//PE_145 replaced by PE

//PE_144 replaced by PE

//PE_143 replaced by PE

//PE_142 replaced by PE

//PE_141 replaced by PE

//PE_140 replaced by PE

//PE_139 replaced by PE

//PE_138 replaced by PE

//PE_137 replaced by PE

//PE_136 replaced by PE

//PE_135 replaced by PE

//PE_134 replaced by PE

//PE_133 replaced by PE

//PE_132 replaced by PE

//PE_131 replaced by PE

//PE_130 replaced by PE

//PE_129 replaced by PE

//PE_128 replaced by PE

//PE_127 replaced by PE

//PE_126 replaced by PE

//PE_125 replaced by PE

//PE_124 replaced by PE

//PE_123 replaced by PE

//PE_122 replaced by PE

//PE_121 replaced by PE

//PE_120 replaced by PE

//PE_119 replaced by PE

//PE_118 replaced by PE

//PE_117 replaced by PE

//PE_116 replaced by PE

//PE_115 replaced by PE

//PE_114 replaced by PE

//PE_113 replaced by PE

//PE_112 replaced by PE

//PE_111 replaced by PE

//PE_110 replaced by PE

//PE_109 replaced by PE

//PE_108 replaced by PE

//PE_107 replaced by PE

//PE_106 replaced by PE

//PE_105 replaced by PE

//PE_104 replaced by PE

//PE_103 replaced by PE

//PE_102 replaced by PE

//PE_101 replaced by PE

//PE_100 replaced by PE

//PE_99 replaced by PE

//PE_98 replaced by PE

//PE_97 replaced by PE

//PE_96 replaced by PE

//PE_95 replaced by PE

//PE_94 replaced by PE

//PE_93 replaced by PE

//PE_92 replaced by PE

//PE_91 replaced by PE

//PE_90 replaced by PE

//PE_89 replaced by PE

//PE_88 replaced by PE

//PE_87 replaced by PE

//PE_86 replaced by PE

//PE_85 replaced by PE

//PE_84 replaced by PE

//PE_83 replaced by PE

//PE_82 replaced by PE

//PE_81 replaced by PE

//PE_80 replaced by PE

//PE_79 replaced by PE

//PE_78 replaced by PE

//PE_77 replaced by PE

//PE_76 replaced by PE

//PE_75 replaced by PE

//PE_74 replaced by PE

//PE_73 replaced by PE

//PE_72 replaced by PE

//PE_71 replaced by PE

//PE_70 replaced by PE

//PE_69 replaced by PE

//PE_68 replaced by PE

//PE_67 replaced by PE

//PE_66 replaced by PE

//PE_65 replaced by PE

//PE_64 replaced by PE

//PE_63 replaced by PE

//PE_62 replaced by PE

//PE_61 replaced by PE

//PE_60 replaced by PE

//PE_59 replaced by PE

//PE_58 replaced by PE

//PE_57 replaced by PE

//PE_56 replaced by PE

//PE_55 replaced by PE

//PE_54 replaced by PE

//PE_53 replaced by PE

//PE_52 replaced by PE

//PE_51 replaced by PE

//PE_50 replaced by PE

//PE_49 replaced by PE

//PE_48 replaced by PE

//PE_47 replaced by PE

//PE_46 replaced by PE

//PE_45 replaced by PE

//PE_44 replaced by PE

//PE_43 replaced by PE

//PE_42 replaced by PE

//PE_41 replaced by PE

//PE_40 replaced by PE

//PE_39 replaced by PE

//PE_38 replaced by PE

//PE_37 replaced by PE

//PE_36 replaced by PE

//PE_35 replaced by PE

//PE_34 replaced by PE

//PE_33 replaced by PE

//PE_32 replaced by PE

//PE_31 replaced by PE

//PE_30 replaced by PE

//PE_29 replaced by PE

//PE_28 replaced by PE

//PE_27 replaced by PE

//PE_26 replaced by PE

//PE_25 replaced by PE

//PE_24 replaced by PE

//PE_23 replaced by PE

//PE_22 replaced by PE

//PE_21 replaced by PE

//PE_20 replaced by PE

//PE_19 replaced by PE

//PE_18 replaced by PE

//PE_17 replaced by PE

//PE_16 replaced by PE

//PE_15 replaced by PE

//PE_14 replaced by PE

//PE_13 replaced by PE

//PE_12 replaced by PE

//PE_11 replaced by PE

//PE_10 replaced by PE

//PE_9 replaced by PE

//PE_8 replaced by PE

//PE_7 replaced by PE

//PE_6 replaced by PE

//PE_5 replaced by PE

//PE_4 replaced by PE

//PE_3 replaced by PE

//PE_2 replaced by PE

//PE_1 replaced by PE

module PE (
  input      [7:0]    activate,
  input      [7:0]    weight,
  input               valid,
  input      [15:0]   signCount,
  output     [7:0]    acount,
  output     [7:0]    bcount,
  output reg [31:0]   PE_OUT,
  output              finish,
  input               clk,
  input               reset
);

  wire       [15:0]   dsp_P;
  wire       [31:0]   _zz_reg1;
  wire       [31:0]   _zz_reg1_1;
  wire       [31:0]   _zz_reg1_2;
  reg        [31:0]   reg1;
  reg                 valid_regNext;
  reg                 valid_regNext_regNext;
  reg        [15:0]   finishCnt_count;
  wire                finishCnt_valid;
  reg                 valid_regNext_1;
  reg        [7:0]    activate_regNext;
  reg        [7:0]    weight_regNext;

  assign _zz_reg1 = {{16{dsp_P[15]}}, dsp_P};
  assign _zz_reg1_1 = 32'h0;
  assign _zz_reg1_2 = {{16{dsp_P[15]}}, dsp_P};
  dsp_marco dsp (
    .CLK (clk          ), //i
    .A   (activate[7:0]), //i
    .B   (weight[7:0]  ), //i
    .P   (dsp_P[15:0]  )  //o
  );
  assign finishCnt_valid = ((finishCnt_count == signCount) && valid_regNext_regNext);
  assign finish = finishCnt_valid;
  always @(*) begin
    PE_OUT = 32'h0;
    if(finishCnt_valid) begin
      PE_OUT = reg1;
    end
  end

  assign acount = activate_regNext;
  assign bcount = weight_regNext;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      reg1 <= 32'h0;
      finishCnt_count <= 16'h0;
    end else begin
      if(valid_regNext_regNext) begin
        if(finishCnt_valid) begin
          finishCnt_count <= 16'h0;
        end else begin
          finishCnt_count <= (finishCnt_count + 16'h0001);
        end
      end
      if(finishCnt_valid) begin
        reg1 <= (valid ? _zz_reg1 : _zz_reg1_1);
      end else begin
        if(valid_regNext_1) begin
          reg1 <= ($signed(_zz_reg1_2) + $signed(reg1));
        end
      end
    end
  end

  always @(posedge clk) begin
    valid_regNext <= valid;
    valid_regNext_regNext <= valid_regNext;
    valid_regNext_1 <= valid;
    activate_regNext <= activate;
    weight_regNext <= weight;
  end


endmodule

module Img2Col_OutPut (
  input               start,
  input               NewAddrIn_valid,
  output              NewAddrIn_ready,
  input      [15:0]   NewAddrIn_payload,
  output              SA_Idle,
  output     [15:0]   Raddr,
  output              Raddr_Valid,
  output              SA_End,
  input      [4:0]    Stride,
  input      [4:0]    Kernel_Size,
  input      [15:0]   Window_Size,
  input      [15:0]   InFeature_Size,
  input      [15:0]   InFeature_Channel,
  input      [15:0]   OutFeature_Channel,
  input      [15:0]   OutFeature_Size,
  input      [15:0]   OutCol_Count_Times,
  input      [15:0]   InCol_Count_Times,
  input      [15:0]   OutFeature_Channel_Count_Times,
  input      [12:0]   Sliding_Size,
  input               mReady,
  input               Fifo_Clear,
  output reg          AddrReceived,
  input               LayerEnd,
  output              SA_Row_Cnt_Valid,
  input               clk,
  input               reset
);
  localparam IMG2COL_OUTPUT_ENUM_IDLE = 7'd1;
  localparam IMG2COL_OUTPUT_ENUM_INIT = 7'd2;
  localparam IMG2COL_OUTPUT_ENUM_INIT_ADDR = 7'd4;
  localparam IMG2COL_OUTPUT_ENUM_SA_COMPUTE = 7'd8;
  localparam IMG2COL_OUTPUT_ENUM_UPDATE_ADDR = 7'd16;
  localparam IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY = 7'd32;
  localparam IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR = 7'd64;

  reg                 RaddrFifo1_io_push_valid;
  reg        [15:0]   RaddrFifo1_io_push_payload;
  reg                 RaddrFifo1_io_pop_ready;
  wire                RaddrFifo1_io_flush;
  wire                RaddrFifo1_io_push_ready;
  wire                RaddrFifo1_io_pop_valid;
  wire       [15:0]   RaddrFifo1_io_pop_payload;
  wire       [5:0]    RaddrFifo1_io_occupancy;
  wire       [5:0]    RaddrFifo1_io_availability;
  wire       [4:0]    _zz_Raddr_Init_Cnt_valid;
  wire       [4:0]    _zz_Raddr_Update_Cnt_valid;
  wire       [12:0]   _zz_In_Channel_Process_Cnt_valid;
  wire       [12:0]   _zz_In_Channel_Process_Cnt_valid_1;
  wire       [15:0]   _zz_Window_Col_Cnt_valid;
  wire       [4:0]    _zz_Window_Col_Cnt_valid_1;
  wire       [15:0]   _zz_Window_Row_Cnt_valid;
  wire       [4:0]    _zz_Window_Row_Cnt_valid_1;
  wire       [15:0]   _zz_Out_Channel_Cnt_valid;
  wire       [15:0]   _zz_Out_Col_Cnt_valid;
  wire       [15:0]   _zz_when_Data_Generate_V2_l498;
  wire       [15:0]   _zz_when_Data_Generate_V2_l498_1;
  wire       [15:0]   _zz_WindowSize_Cnt_valid;
  wire       [15:0]   _zz_WindowSize_Cnt_valid_1;
  wire       [31:0]   _zz_Kernel_Base_Addr;
  wire       [15:0]   _zz_Kernel_Base_Addr_1;
  wire       [31:0]   _zz_Kernel_Addr;
  wire       [15:0]   _zz_Kernel_Addr_1;
  wire       [31:0]   _zz_Kernel_Addr_2;
  wire       [31:0]   _zz_Kernel_Addr_3;
  wire       [31:0]   _zz_Kernel_Addr_4;
  wire       [31:0]   _zz_Raddr;
  wire       [31:0]   _zz_Raddr_1;
  reg                 start_regNext;
  wire                when_Data_Generate_V2_l344;
  reg        [6:0]    Fsm_currentState;
  reg        [6:0]    Fsm_nextState;
  wire                Fsm_Init_End;
  wire                Fsm_Addr_Inited;
  wire                Fsm_SA_Computed;
  wire                Fsm_Addr_Updated;
  wire                Fsm_LayerEnd;
  wire                Fsm_NextReady;
  wire                Fsm_Fifo_Clear;
  wire                when_Data_Generate_V2_l376;
  wire                when_WaCounter_l19;
  reg        [2:0]    Init_Count_count;
  reg                 Init_Count_valid;
  wire                when_WaCounter_l14;
  reg        [15:0]   Row_Base_Addr;
  wire                Img2Col_SubModule_RaddrFifo1_io_pop_fire;
  wire                Img2Col_SubModule_RaddrFifo1_io_push_fire;
  wire                when_WaCounter_l40;
  reg        [4:0]    Raddr_Init_Cnt_count;
  wire                Raddr_Init_Cnt_valid;
  wire                Img2Col_SubModule_RaddrFifo1_io_push_fire_1;
  wire                when_WaCounter_l40_1;
  reg        [4:0]    Raddr_Update_Cnt_count;
  wire                Raddr_Update_Cnt_valid;
  wire                when_Data_Generate_V2_l463;
  wire                when_WaCounter_l40_2;
  reg        [2:0]    SA_Row_Cnt_count;
  reg                 SA_Row_Cnt_valid_1;
  reg        [12:0]   In_Channel_Process_Cnt_count;
  wire                In_Channel_Process_Cnt_valid;
  reg        [15:0]   Window_Col_Cnt_count;
  wire                Window_Col_Cnt_valid;
  reg        [15:0]   Window_Row_Cnt_count;
  wire                Window_Row_Cnt_valid;
  reg        [15:0]   Out_Channel_Cnt_count;
  wire                Out_Channel_Cnt_valid;
  reg        [15:0]   Out_Col_Cnt_count;
  wire                Out_Col_Cnt_valid;
  reg        [15:0]   OutFeature_Col_Lefted;
  wire                when_Data_Generate_V2_l495;
  wire                when_Data_Generate_V2_l498;
  reg        [12:0]   WindowSize_Cnt_count;
  wire                WindowSize_Cnt_valid;
  reg        [31:0]   Kernel_Addr;
  reg        [31:0]   Kernel_Base_Addr;
  wire                when_Data_Generate_V2_l523;
  wire                when_Data_Generate_V2_l533;
  wire                Img2Col_SubModule_RaddrFifo1_io_push_fire_2;
  wire                when_Data_Generate_V2_l537;
  `ifndef SYNTHESIS
  reg [119:0] Fsm_currentState_string;
  reg [119:0] Fsm_nextState_string;
  `endif


  assign _zz_Raddr_Init_Cnt_valid = (Kernel_Size - 5'h01);
  assign _zz_Raddr_Update_Cnt_valid = (Stride - 5'h01);
  assign _zz_In_Channel_Process_Cnt_valid = (_zz_In_Channel_Process_Cnt_valid_1 - 13'h0001);
  assign _zz_In_Channel_Process_Cnt_valid_1 = (InFeature_Channel >>> 3);
  assign _zz_Window_Col_Cnt_valid_1 = (Kernel_Size - 5'h01);
  assign _zz_Window_Col_Cnt_valid = {11'd0, _zz_Window_Col_Cnt_valid_1};
  assign _zz_Window_Row_Cnt_valid_1 = (Kernel_Size - 5'h01);
  assign _zz_Window_Row_Cnt_valid = {11'd0, _zz_Window_Row_Cnt_valid_1};
  assign _zz_Out_Channel_Cnt_valid = (OutFeature_Channel_Count_Times - 16'h0001);
  assign _zz_Out_Col_Cnt_valid = (OutCol_Count_Times - 16'h0001);
  assign _zz_when_Data_Generate_V2_l498 = {13'd0, SA_Row_Cnt_count};
  assign _zz_when_Data_Generate_V2_l498_1 = (OutFeature_Col_Lefted - 16'h0001);
  assign _zz_WindowSize_Cnt_valid = {3'd0, WindowSize_Cnt_count};
  assign _zz_WindowSize_Cnt_valid_1 = (Window_Size - 16'h0001);
  assign _zz_Kernel_Base_Addr_1 = ({3'd0,Sliding_Size} <<< 3);
  assign _zz_Kernel_Base_Addr = {16'd0, _zz_Kernel_Base_Addr_1};
  assign _zz_Kernel_Addr_1 = ({3'd0,Sliding_Size} <<< 3);
  assign _zz_Kernel_Addr = {16'd0, _zz_Kernel_Addr_1};
  assign _zz_Kernel_Addr_2 = (Kernel_Base_Addr + _zz_Kernel_Addr_3);
  assign _zz_Kernel_Addr_3 = {19'd0, WindowSize_Cnt_count};
  assign _zz_Kernel_Addr_4 = {19'd0, Sliding_Size};
  assign _zz_Raddr = (Kernel_Addr + _zz_Raddr_1);
  assign _zz_Raddr_1 = {16'd0, Row_Base_Addr};
  WaddrOffset_Fifo_2 RaddrFifo1 (
    .io_push_valid   (RaddrFifo1_io_push_valid        ), //i
    .io_push_ready   (RaddrFifo1_io_push_ready        ), //o
    .io_push_payload (RaddrFifo1_io_push_payload[15:0]), //i
    .io_pop_valid    (RaddrFifo1_io_pop_valid         ), //o
    .io_pop_ready    (RaddrFifo1_io_pop_ready         ), //i
    .io_pop_payload  (RaddrFifo1_io_pop_payload[15:0] ), //o
    .io_flush        (RaddrFifo1_io_flush             ), //i
    .io_occupancy    (RaddrFifo1_io_occupancy[5:0]    ), //o
    .io_availability (RaddrFifo1_io_availability[5:0] ), //o
    .clk             (clk                             ), //i
    .reset           (reset                           )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(Fsm_currentState)
      IMG2COL_OUTPUT_ENUM_IDLE : Fsm_currentState_string = "IDLE           ";
      IMG2COL_OUTPUT_ENUM_INIT : Fsm_currentState_string = "INIT           ";
      IMG2COL_OUTPUT_ENUM_INIT_ADDR : Fsm_currentState_string = "INIT_ADDR      ";
      IMG2COL_OUTPUT_ENUM_SA_COMPUTE : Fsm_currentState_string = "SA_COMPUTE     ";
      IMG2COL_OUTPUT_ENUM_UPDATE_ADDR : Fsm_currentState_string = "UPDATE_ADDR    ";
      IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY : Fsm_currentState_string = "WAIT_NEXT_READY";
      IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR : Fsm_currentState_string = "WAIT_FIFO_CLEAR";
      default : Fsm_currentState_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(Fsm_nextState)
      IMG2COL_OUTPUT_ENUM_IDLE : Fsm_nextState_string = "IDLE           ";
      IMG2COL_OUTPUT_ENUM_INIT : Fsm_nextState_string = "INIT           ";
      IMG2COL_OUTPUT_ENUM_INIT_ADDR : Fsm_nextState_string = "INIT_ADDR      ";
      IMG2COL_OUTPUT_ENUM_SA_COMPUTE : Fsm_nextState_string = "SA_COMPUTE     ";
      IMG2COL_OUTPUT_ENUM_UPDATE_ADDR : Fsm_nextState_string = "UPDATE_ADDR    ";
      IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY : Fsm_nextState_string = "WAIT_NEXT_READY";
      IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR : Fsm_nextState_string = "WAIT_FIFO_CLEAR";
      default : Fsm_nextState_string = "???????????????";
    endcase
  end
  `endif

  assign when_Data_Generate_V2_l344 = (start && (! start_regNext));
  always @(*) begin
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_IDLE) == IMG2COL_OUTPUT_ENUM_IDLE) : begin
        if(when_Data_Generate_V2_l344) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_INIT;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_IDLE;
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_INIT) == IMG2COL_OUTPUT_ENUM_INIT) : begin
        if(Fsm_Init_End) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_INIT_ADDR;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_INIT;
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_INIT_ADDR) == IMG2COL_OUTPUT_ENUM_INIT_ADDR) : begin
        if(Fsm_Addr_Inited) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_INIT_ADDR;
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY) == IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY) : begin
        if(Fsm_NextReady) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_SA_COMPUTE;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY;
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) == IMG2COL_OUTPUT_ENUM_SA_COMPUTE) : begin
        if(Fsm_LayerEnd) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_IDLE;
        end else begin
          if(Fsm_SA_Computed) begin
            Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR;
          end else begin
            if(when_Data_Generate_V2_l376) begin
              Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY;
            end else begin
              Fsm_nextState = IMG2COL_OUTPUT_ENUM_SA_COMPUTE;
            end
          end
        end
      end
      (((Fsm_currentState) & IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR) == IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR) : begin
        if(Fsm_Fifo_Clear) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_UPDATE_ADDR;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_FIFO_CLEAR;
        end
      end
      default : begin
        if(Fsm_Addr_Updated) begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY;
        end else begin
          Fsm_nextState = IMG2COL_OUTPUT_ENUM_UPDATE_ADDR;
        end
      end
    endcase
  end

  assign when_Data_Generate_V2_l376 = (! Fsm_NextReady);
  assign when_WaCounter_l19 = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT) != 7'b0000000);
  assign when_WaCounter_l14 = (Init_Count_count == 3'b101);
  always @(*) begin
    if(when_WaCounter_l14) begin
      Init_Count_valid = 1'b1;
    end else begin
      Init_Count_valid = 1'b0;
    end
  end

  assign Fsm_Init_End = Init_Count_valid;
  assign Fsm_Fifo_Clear = Fifo_Clear;
  assign NewAddrIn_ready = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT_ADDR) != 7'b0000000) || ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 7'b0000000));
  always @(*) begin
    RaddrFifo1_io_push_valid = 1'b0;
    if(when_Data_Generate_V2_l533) begin
      RaddrFifo1_io_push_valid = NewAddrIn_valid;
    end else begin
      if(when_Data_Generate_V2_l537) begin
        RaddrFifo1_io_push_valid = NewAddrIn_valid;
      end else begin
        RaddrFifo1_io_push_valid = Window_Col_Cnt_valid;
      end
    end
  end

  always @(*) begin
    RaddrFifo1_io_pop_ready = 1'b0;
    if(when_Data_Generate_V2_l463) begin
      RaddrFifo1_io_pop_ready = 1'b1;
    end
    if(!when_Data_Generate_V2_l533) begin
      if(when_Data_Generate_V2_l537) begin
        RaddrFifo1_io_pop_ready = Img2Col_SubModule_RaddrFifo1_io_push_fire_2;
      end
    end
    if(Window_Col_Cnt_valid) begin
      RaddrFifo1_io_pop_ready = 1'b1;
    end
  end

  assign Img2Col_SubModule_RaddrFifo1_io_pop_fire = (RaddrFifo1_io_pop_valid && RaddrFifo1_io_pop_ready);
  assign Img2Col_SubModule_RaddrFifo1_io_push_fire = (RaddrFifo1_io_push_valid && RaddrFifo1_io_push_ready);
  assign when_WaCounter_l40 = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT_ADDR) != 7'b0000000) && Img2Col_SubModule_RaddrFifo1_io_push_fire);
  assign Raddr_Init_Cnt_valid = ((Raddr_Init_Cnt_count == _zz_Raddr_Init_Cnt_valid) && when_WaCounter_l40);
  assign Fsm_Addr_Inited = Raddr_Init_Cnt_valid;
  assign Img2Col_SubModule_RaddrFifo1_io_push_fire_1 = (RaddrFifo1_io_push_valid && RaddrFifo1_io_push_ready);
  assign when_WaCounter_l40_1 = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 7'b0000000) && Img2Col_SubModule_RaddrFifo1_io_push_fire_1);
  assign Raddr_Update_Cnt_valid = ((Raddr_Update_Cnt_count == _zz_Raddr_Update_Cnt_valid) && when_WaCounter_l40_1);
  assign Fsm_Addr_Updated = Raddr_Update_Cnt_valid;
  assign Fsm_NextReady = mReady;
  always @(*) begin
    AddrReceived = 1'b0;
    if(when_Data_Generate_V2_l463) begin
      AddrReceived = 1'b1;
    end
  end

  assign when_Data_Generate_V2_l463 = ((((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT_ADDR) != 7'b0000000) && ((Fsm_nextState & IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY) != 7'b0000000)) || (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 7'b0000000) && ((Fsm_nextState & IMG2COL_OUTPUT_ENUM_WAIT_NEXT_READY) != 7'b0000000)));
  assign when_WaCounter_l40_2 = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) != 7'b0000000) && mReady);
  always @(*) begin
    SA_Row_Cnt_valid_1 = ((SA_Row_Cnt_count == 3'b111) && when_WaCounter_l40_2);
    if(when_Data_Generate_V2_l498) begin
      SA_Row_Cnt_valid_1 = 1'b1;
    end
  end

  assign SA_Row_Cnt_Valid = SA_Row_Cnt_valid_1;
  assign In_Channel_Process_Cnt_valid = ((In_Channel_Process_Cnt_count == _zz_In_Channel_Process_Cnt_valid) && SA_Row_Cnt_valid_1);
  assign Window_Col_Cnt_valid = ((Window_Col_Cnt_count == _zz_Window_Col_Cnt_valid) && In_Channel_Process_Cnt_valid);
  assign Window_Row_Cnt_valid = ((Window_Row_Cnt_count == _zz_Window_Row_Cnt_valid) && Window_Col_Cnt_valid);
  assign Out_Channel_Cnt_valid = ((Out_Channel_Cnt_count == _zz_Out_Channel_Cnt_valid) && Window_Row_Cnt_valid);
  assign Out_Col_Cnt_valid = ((Out_Col_Cnt_count == _zz_Out_Col_Cnt_valid) && Out_Channel_Cnt_valid);
  assign SA_End = Out_Col_Cnt_valid;
  assign when_Data_Generate_V2_l495 = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT) != 7'b0000000);
  assign when_Data_Generate_V2_l498 = (((_zz_when_Data_Generate_V2_l498 == _zz_when_Data_Generate_V2_l498_1) && mReady) && ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) != 7'b0000000));
  assign WindowSize_Cnt_valid = ((_zz_WindowSize_Cnt_valid == _zz_WindowSize_Cnt_valid_1) && SA_Row_Cnt_valid_1);
  assign when_Data_Generate_V2_l523 = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) != 7'b0000000) && mReady);
  assign Raddr = _zz_Raddr[15:0];
  assign Fsm_SA_Computed = Out_Col_Cnt_valid;
  assign SA_Idle = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_IDLE) != 7'b0000000) || ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 7'b0000000));
  assign when_Data_Generate_V2_l533 = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_INIT_ADDR) != 7'b0000000);
  always @(*) begin
    if(when_Data_Generate_V2_l533) begin
      RaddrFifo1_io_push_payload = NewAddrIn_payload;
    end else begin
      if(when_Data_Generate_V2_l537) begin
        RaddrFifo1_io_push_payload = NewAddrIn_payload;
      end else begin
        RaddrFifo1_io_push_payload = Row_Base_Addr;
      end
    end
  end

  assign Img2Col_SubModule_RaddrFifo1_io_push_fire_2 = (RaddrFifo1_io_push_valid && RaddrFifo1_io_push_ready);
  assign when_Data_Generate_V2_l537 = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_UPDATE_ADDR) != 7'b0000000);
  assign Raddr_Valid = (((Fsm_currentState & IMG2COL_OUTPUT_ENUM_SA_COMPUTE) != 7'b0000000) && mReady);
  assign Fsm_LayerEnd = LayerEnd;
  assign RaddrFifo1_io_flush = ((Fsm_currentState & IMG2COL_OUTPUT_ENUM_IDLE) != 7'b0000000);
  always @(posedge clk) begin
    start_regNext <= start;
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      Fsm_currentState <= IMG2COL_OUTPUT_ENUM_IDLE;
      Init_Count_count <= 3'b000;
      Row_Base_Addr <= 16'h0;
      Raddr_Init_Cnt_count <= 5'h0;
      Raddr_Update_Cnt_count <= 5'h0;
      SA_Row_Cnt_count <= 3'b000;
      In_Channel_Process_Cnt_count <= 13'h0;
      Window_Col_Cnt_count <= 16'h0;
      Window_Row_Cnt_count <= 16'h0;
      Out_Channel_Cnt_count <= 16'h0;
      Out_Col_Cnt_count <= 16'h0;
      OutFeature_Col_Lefted <= 16'h0;
      WindowSize_Cnt_count <= 13'h0;
      Kernel_Addr <= 32'h0;
      Kernel_Base_Addr <= 32'h0;
    end else begin
      Fsm_currentState <= Fsm_nextState;
      if(when_WaCounter_l19) begin
        Init_Count_count <= (Init_Count_count + 3'b001);
        if(Init_Count_valid) begin
          Init_Count_count <= 3'b000;
        end
      end
      if(Img2Col_SubModule_RaddrFifo1_io_pop_fire) begin
        Row_Base_Addr <= RaddrFifo1_io_pop_payload;
      end
      if(when_WaCounter_l40) begin
        if(Raddr_Init_Cnt_valid) begin
          Raddr_Init_Cnt_count <= 5'h0;
        end else begin
          Raddr_Init_Cnt_count <= (Raddr_Init_Cnt_count + 5'h01);
        end
      end
      if(when_WaCounter_l40_1) begin
        if(Raddr_Update_Cnt_valid) begin
          Raddr_Update_Cnt_count <= 5'h0;
        end else begin
          Raddr_Update_Cnt_count <= (Raddr_Update_Cnt_count + 5'h01);
        end
      end
      if(when_WaCounter_l40_2) begin
        if(SA_Row_Cnt_valid_1) begin
          SA_Row_Cnt_count <= 3'b000;
        end else begin
          SA_Row_Cnt_count <= (SA_Row_Cnt_count + 3'b001);
        end
      end
      if(SA_Row_Cnt_valid_1) begin
        if(In_Channel_Process_Cnt_valid) begin
          In_Channel_Process_Cnt_count <= 13'h0;
        end else begin
          In_Channel_Process_Cnt_count <= (In_Channel_Process_Cnt_count + 13'h0001);
        end
      end
      if(In_Channel_Process_Cnt_valid) begin
        if(Window_Col_Cnt_valid) begin
          Window_Col_Cnt_count <= 16'h0;
        end else begin
          Window_Col_Cnt_count <= (Window_Col_Cnt_count + 16'h0001);
        end
      end
      if(Window_Col_Cnt_valid) begin
        if(Window_Row_Cnt_valid) begin
          Window_Row_Cnt_count <= 16'h0;
        end else begin
          Window_Row_Cnt_count <= (Window_Row_Cnt_count + 16'h0001);
        end
      end
      if(Window_Row_Cnt_valid) begin
        if(Out_Channel_Cnt_valid) begin
          Out_Channel_Cnt_count <= 16'h0;
        end else begin
          Out_Channel_Cnt_count <= (Out_Channel_Cnt_count + 16'h0001);
        end
      end
      if(Out_Channel_Cnt_valid) begin
        if(Out_Col_Cnt_valid) begin
          Out_Col_Cnt_count <= 16'h0;
        end else begin
          Out_Col_Cnt_count <= (Out_Col_Cnt_count + 16'h0001);
        end
      end
      if(Out_Col_Cnt_valid) begin
        OutFeature_Col_Lefted <= OutFeature_Size;
      end else begin
        if(Out_Channel_Cnt_valid) begin
          OutFeature_Col_Lefted <= (OutFeature_Col_Lefted - 16'h0008);
        end else begin
          if(when_Data_Generate_V2_l495) begin
            OutFeature_Col_Lefted <= OutFeature_Size;
          end
        end
      end
      if(when_Data_Generate_V2_l498) begin
        SA_Row_Cnt_count <= 3'b000;
      end
      if(SA_Row_Cnt_valid_1) begin
        if(WindowSize_Cnt_valid) begin
          WindowSize_Cnt_count <= 13'h0;
        end else begin
          WindowSize_Cnt_count <= (WindowSize_Cnt_count + 13'h0001);
        end
      end
      if(Out_Col_Cnt_valid) begin
        Kernel_Base_Addr <= 32'h0;
      end else begin
        if(Out_Channel_Cnt_valid) begin
          Kernel_Base_Addr <= (Kernel_Base_Addr + _zz_Kernel_Base_Addr);
        end
      end
      if(Out_Col_Cnt_valid) begin
        Kernel_Addr <= 32'h0;
      end else begin
        if(Out_Channel_Cnt_valid) begin
          Kernel_Addr <= (Kernel_Base_Addr + _zz_Kernel_Addr);
        end else begin
          if(Window_Row_Cnt_valid) begin
            Kernel_Addr <= Kernel_Base_Addr;
          end else begin
            if(WindowSize_Cnt_valid) begin
              Kernel_Addr <= Kernel_Base_Addr;
            end else begin
              if(SA_Row_Cnt_valid_1) begin
                Kernel_Addr <= (_zz_Kernel_Addr_2 + 32'h00000001);
              end else begin
                if(when_Data_Generate_V2_l523) begin
                  Kernel_Addr <= (Kernel_Addr + _zz_Kernel_Addr_4);
                end
              end
            end
          end
        end
      end
    end
  end


endmodule

//WaddrOffset_Fifo_1 replaced by WaddrOffset_Fifo_2

//WaddrOffset_Fifo replaced by WaddrOffset_Fifo_2

module WaddrOffset_Fifo_2 (
  input               io_push_valid,
  output              io_push_ready,
  input      [15:0]   io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [15:0]   io_pop_payload,
  input               io_flush,
  output reg [5:0]    io_occupancy,
  output reg [5:0]    io_availability,
  input               clk,
  input               reset
);

  reg        [15:0]   _zz_logic_ram_port0;
  wire       [5:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [5:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [15:0]   _zz_logic_ram_port_1;
  wire       [5:0]    _zz_io_occupancy;
  wire       [5:0]    _zz_io_availability;
  wire       [5:0]    _zz_io_availability_1;
  wire       [5:0]    _zz_io_availability_2;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [5:0]    logic_pushPtr_valueNext;
  reg        [5:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [5:0]    logic_popPtr_valueNext;
  reg        [5:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1122;
  wire       [5:0]    logic_ptrDif;
  reg [15:0] logic_ram [0:32];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {5'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {5'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_occupancy = (6'h21 + logic_ptrDif);
  assign _zz_io_availability = (6'h21 + _zz_io_availability_1);
  assign _zz_io_availability_1 = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_availability_2 = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  assign _zz_logic_ram_port_1 = io_push_payload;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 6'h20);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    if(logic_pushPtr_willOverflow) begin
      logic_pushPtr_valueNext = 6'h0;
    end else begin
      logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    end
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 6'h0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 6'h20);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    if(logic_popPtr_willOverflow) begin
      logic_popPtr_valueNext = 6'h0;
    end else begin
      logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    end
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 6'h0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1122 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  always @(*) begin
    if(logic_ptrMatch) begin
      io_occupancy = (logic_risingOccupancy ? 6'h21 : 6'h0);
    end else begin
      io_occupancy = ((logic_popPtr_value < logic_pushPtr_value) ? logic_ptrDif : _zz_io_occupancy);
    end
  end

  always @(*) begin
    if(logic_ptrMatch) begin
      io_availability = (logic_risingOccupancy ? 6'h0 : 6'h21);
    end else begin
      io_availability = ((logic_popPtr_value < logic_pushPtr_value) ? _zz_io_availability : _zz_io_availability_2);
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_pushPtr_value <= 6'h0;
      logic_popPtr_value <= 6'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1122) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule
